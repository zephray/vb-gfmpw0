magic
tech gf180mcuC
magscale 1 5
timestamp 1670290360
<< obsm1 >>
rect 672 855 149296 148329
<< metal2 >>
rect 2184 149600 2240 150000
rect 3472 149600 3528 150000
rect 4760 149600 4816 150000
rect 6048 149600 6104 150000
rect 7336 149600 7392 150000
rect 8624 149600 8680 150000
rect 9912 149600 9968 150000
rect 11200 149600 11256 150000
rect 12488 149600 12544 150000
rect 13776 149600 13832 150000
rect 15064 149600 15120 150000
rect 16352 149600 16408 150000
rect 17640 149600 17696 150000
rect 18928 149600 18984 150000
rect 20216 149600 20272 150000
rect 21504 149600 21560 150000
rect 22792 149600 22848 150000
rect 24080 149600 24136 150000
rect 25368 149600 25424 150000
rect 26656 149600 26712 150000
rect 27944 149600 28000 150000
rect 29232 149600 29288 150000
rect 30520 149600 30576 150000
rect 31808 149600 31864 150000
rect 33096 149600 33152 150000
rect 34384 149600 34440 150000
rect 35672 149600 35728 150000
rect 36960 149600 37016 150000
rect 38248 149600 38304 150000
rect 39536 149600 39592 150000
rect 40824 149600 40880 150000
rect 42112 149600 42168 150000
rect 43400 149600 43456 150000
rect 44688 149600 44744 150000
rect 45976 149600 46032 150000
rect 47264 149600 47320 150000
rect 48552 149600 48608 150000
rect 49840 149600 49896 150000
rect 51128 149600 51184 150000
rect 52416 149600 52472 150000
rect 53704 149600 53760 150000
rect 54992 149600 55048 150000
rect 56280 149600 56336 150000
rect 57568 149600 57624 150000
rect 58856 149600 58912 150000
rect 60144 149600 60200 150000
rect 61432 149600 61488 150000
rect 62720 149600 62776 150000
rect 64008 149600 64064 150000
rect 65296 149600 65352 150000
rect 66584 149600 66640 150000
rect 67872 149600 67928 150000
rect 69160 149600 69216 150000
rect 70448 149600 70504 150000
rect 71736 149600 71792 150000
rect 73024 149600 73080 150000
rect 74312 149600 74368 150000
rect 75600 149600 75656 150000
rect 76888 149600 76944 150000
rect 78176 149600 78232 150000
rect 79464 149600 79520 150000
rect 80752 149600 80808 150000
rect 82040 149600 82096 150000
rect 83328 149600 83384 150000
rect 84616 149600 84672 150000
rect 85904 149600 85960 150000
rect 87192 149600 87248 150000
rect 88480 149600 88536 150000
rect 89768 149600 89824 150000
rect 91056 149600 91112 150000
rect 92344 149600 92400 150000
rect 93632 149600 93688 150000
rect 94920 149600 94976 150000
rect 96208 149600 96264 150000
rect 97496 149600 97552 150000
rect 98784 149600 98840 150000
rect 100072 149600 100128 150000
rect 101360 149600 101416 150000
rect 102648 149600 102704 150000
rect 103936 149600 103992 150000
rect 105224 149600 105280 150000
rect 106512 149600 106568 150000
rect 107800 149600 107856 150000
rect 109088 149600 109144 150000
rect 110376 149600 110432 150000
rect 111664 149600 111720 150000
rect 112952 149600 113008 150000
rect 114240 149600 114296 150000
rect 115528 149600 115584 150000
rect 116816 149600 116872 150000
rect 118104 149600 118160 150000
rect 119392 149600 119448 150000
rect 120680 149600 120736 150000
rect 121968 149600 122024 150000
rect 123256 149600 123312 150000
rect 124544 149600 124600 150000
rect 125832 149600 125888 150000
rect 127120 149600 127176 150000
rect 128408 149600 128464 150000
rect 129696 149600 129752 150000
rect 130984 149600 131040 150000
rect 132272 149600 132328 150000
rect 133560 149600 133616 150000
rect 134848 149600 134904 150000
rect 136136 149600 136192 150000
rect 137424 149600 137480 150000
rect 138712 149600 138768 150000
rect 140000 149600 140056 150000
rect 141288 149600 141344 150000
rect 142576 149600 142632 150000
rect 143864 149600 143920 150000
rect 145152 149600 145208 150000
rect 146440 149600 146496 150000
rect 147728 149600 147784 150000
rect 7728 0 7784 400
rect 8176 0 8232 400
rect 8624 0 8680 400
rect 9072 0 9128 400
rect 9520 0 9576 400
rect 9968 0 10024 400
rect 10416 0 10472 400
rect 10864 0 10920 400
rect 11312 0 11368 400
rect 11760 0 11816 400
rect 12208 0 12264 400
rect 12656 0 12712 400
rect 13104 0 13160 400
rect 13552 0 13608 400
rect 14000 0 14056 400
rect 14448 0 14504 400
rect 14896 0 14952 400
rect 15344 0 15400 400
rect 15792 0 15848 400
rect 16240 0 16296 400
rect 16688 0 16744 400
rect 17136 0 17192 400
rect 17584 0 17640 400
rect 18032 0 18088 400
rect 18480 0 18536 400
rect 18928 0 18984 400
rect 19376 0 19432 400
rect 19824 0 19880 400
rect 20272 0 20328 400
rect 20720 0 20776 400
rect 21168 0 21224 400
rect 21616 0 21672 400
rect 22064 0 22120 400
rect 22512 0 22568 400
rect 22960 0 23016 400
rect 23408 0 23464 400
rect 23856 0 23912 400
rect 24304 0 24360 400
rect 24752 0 24808 400
rect 25200 0 25256 400
rect 25648 0 25704 400
rect 26096 0 26152 400
rect 26544 0 26600 400
rect 26992 0 27048 400
rect 27440 0 27496 400
rect 27888 0 27944 400
rect 28336 0 28392 400
rect 28784 0 28840 400
rect 29232 0 29288 400
rect 29680 0 29736 400
rect 30128 0 30184 400
rect 30576 0 30632 400
rect 31024 0 31080 400
rect 31472 0 31528 400
rect 31920 0 31976 400
rect 32368 0 32424 400
rect 32816 0 32872 400
rect 33264 0 33320 400
rect 33712 0 33768 400
rect 34160 0 34216 400
rect 34608 0 34664 400
rect 35056 0 35112 400
rect 35504 0 35560 400
rect 35952 0 36008 400
rect 36400 0 36456 400
rect 36848 0 36904 400
rect 37296 0 37352 400
rect 37744 0 37800 400
rect 38192 0 38248 400
rect 38640 0 38696 400
rect 39088 0 39144 400
rect 39536 0 39592 400
rect 39984 0 40040 400
rect 40432 0 40488 400
rect 40880 0 40936 400
rect 41328 0 41384 400
rect 41776 0 41832 400
rect 42224 0 42280 400
rect 42672 0 42728 400
rect 43120 0 43176 400
rect 43568 0 43624 400
rect 44016 0 44072 400
rect 44464 0 44520 400
rect 44912 0 44968 400
rect 45360 0 45416 400
rect 45808 0 45864 400
rect 46256 0 46312 400
rect 46704 0 46760 400
rect 47152 0 47208 400
rect 47600 0 47656 400
rect 48048 0 48104 400
rect 48496 0 48552 400
rect 48944 0 49000 400
rect 49392 0 49448 400
rect 49840 0 49896 400
rect 50288 0 50344 400
rect 50736 0 50792 400
rect 51184 0 51240 400
rect 51632 0 51688 400
rect 52080 0 52136 400
rect 52528 0 52584 400
rect 52976 0 53032 400
rect 53424 0 53480 400
rect 53872 0 53928 400
rect 54320 0 54376 400
rect 54768 0 54824 400
rect 55216 0 55272 400
rect 55664 0 55720 400
rect 56112 0 56168 400
rect 56560 0 56616 400
rect 57008 0 57064 400
rect 57456 0 57512 400
rect 57904 0 57960 400
rect 58352 0 58408 400
rect 58800 0 58856 400
rect 59248 0 59304 400
rect 59696 0 59752 400
rect 60144 0 60200 400
rect 60592 0 60648 400
rect 61040 0 61096 400
rect 61488 0 61544 400
rect 61936 0 61992 400
rect 62384 0 62440 400
rect 62832 0 62888 400
rect 63280 0 63336 400
rect 63728 0 63784 400
rect 64176 0 64232 400
rect 64624 0 64680 400
rect 65072 0 65128 400
rect 65520 0 65576 400
rect 65968 0 66024 400
rect 66416 0 66472 400
rect 66864 0 66920 400
rect 67312 0 67368 400
rect 67760 0 67816 400
rect 68208 0 68264 400
rect 68656 0 68712 400
rect 69104 0 69160 400
rect 69552 0 69608 400
rect 70000 0 70056 400
rect 70448 0 70504 400
rect 70896 0 70952 400
rect 71344 0 71400 400
rect 71792 0 71848 400
rect 72240 0 72296 400
rect 72688 0 72744 400
rect 73136 0 73192 400
rect 73584 0 73640 400
rect 74032 0 74088 400
rect 74480 0 74536 400
rect 74928 0 74984 400
rect 75376 0 75432 400
rect 75824 0 75880 400
rect 76272 0 76328 400
rect 76720 0 76776 400
rect 77168 0 77224 400
rect 77616 0 77672 400
rect 78064 0 78120 400
rect 78512 0 78568 400
rect 78960 0 79016 400
rect 79408 0 79464 400
rect 79856 0 79912 400
rect 80304 0 80360 400
rect 80752 0 80808 400
rect 81200 0 81256 400
rect 81648 0 81704 400
rect 82096 0 82152 400
rect 82544 0 82600 400
rect 82992 0 83048 400
rect 83440 0 83496 400
rect 83888 0 83944 400
rect 84336 0 84392 400
rect 84784 0 84840 400
rect 85232 0 85288 400
rect 85680 0 85736 400
rect 86128 0 86184 400
rect 86576 0 86632 400
rect 87024 0 87080 400
rect 87472 0 87528 400
rect 87920 0 87976 400
rect 88368 0 88424 400
rect 88816 0 88872 400
rect 89264 0 89320 400
rect 89712 0 89768 400
rect 90160 0 90216 400
rect 90608 0 90664 400
rect 91056 0 91112 400
rect 91504 0 91560 400
rect 91952 0 92008 400
rect 92400 0 92456 400
rect 92848 0 92904 400
rect 93296 0 93352 400
rect 93744 0 93800 400
rect 94192 0 94248 400
rect 94640 0 94696 400
rect 95088 0 95144 400
rect 95536 0 95592 400
rect 95984 0 96040 400
rect 96432 0 96488 400
rect 96880 0 96936 400
rect 97328 0 97384 400
rect 97776 0 97832 400
rect 98224 0 98280 400
rect 98672 0 98728 400
rect 99120 0 99176 400
rect 99568 0 99624 400
rect 100016 0 100072 400
rect 100464 0 100520 400
rect 100912 0 100968 400
rect 101360 0 101416 400
rect 101808 0 101864 400
rect 102256 0 102312 400
rect 102704 0 102760 400
rect 103152 0 103208 400
rect 103600 0 103656 400
rect 104048 0 104104 400
rect 104496 0 104552 400
rect 104944 0 105000 400
rect 105392 0 105448 400
rect 105840 0 105896 400
rect 106288 0 106344 400
rect 106736 0 106792 400
rect 107184 0 107240 400
rect 107632 0 107688 400
rect 108080 0 108136 400
rect 108528 0 108584 400
rect 108976 0 109032 400
rect 109424 0 109480 400
rect 109872 0 109928 400
rect 110320 0 110376 400
rect 110768 0 110824 400
rect 111216 0 111272 400
rect 111664 0 111720 400
rect 112112 0 112168 400
rect 112560 0 112616 400
rect 113008 0 113064 400
rect 113456 0 113512 400
rect 113904 0 113960 400
rect 114352 0 114408 400
rect 114800 0 114856 400
rect 115248 0 115304 400
rect 115696 0 115752 400
rect 116144 0 116200 400
rect 116592 0 116648 400
rect 117040 0 117096 400
rect 117488 0 117544 400
rect 117936 0 117992 400
rect 118384 0 118440 400
rect 118832 0 118888 400
rect 119280 0 119336 400
rect 119728 0 119784 400
rect 120176 0 120232 400
rect 120624 0 120680 400
rect 121072 0 121128 400
rect 121520 0 121576 400
rect 121968 0 122024 400
rect 122416 0 122472 400
rect 122864 0 122920 400
rect 123312 0 123368 400
rect 123760 0 123816 400
rect 124208 0 124264 400
rect 124656 0 124712 400
rect 125104 0 125160 400
rect 125552 0 125608 400
rect 126000 0 126056 400
rect 126448 0 126504 400
rect 126896 0 126952 400
rect 127344 0 127400 400
rect 127792 0 127848 400
rect 128240 0 128296 400
rect 128688 0 128744 400
rect 129136 0 129192 400
rect 129584 0 129640 400
rect 130032 0 130088 400
rect 130480 0 130536 400
rect 130928 0 130984 400
rect 131376 0 131432 400
rect 131824 0 131880 400
rect 132272 0 132328 400
rect 132720 0 132776 400
rect 133168 0 133224 400
rect 133616 0 133672 400
rect 134064 0 134120 400
rect 134512 0 134568 400
rect 134960 0 135016 400
rect 135408 0 135464 400
rect 135856 0 135912 400
rect 136304 0 136360 400
rect 136752 0 136808 400
rect 137200 0 137256 400
rect 137648 0 137704 400
rect 138096 0 138152 400
rect 138544 0 138600 400
rect 138992 0 139048 400
rect 139440 0 139496 400
rect 139888 0 139944 400
rect 140336 0 140392 400
rect 140784 0 140840 400
rect 141232 0 141288 400
rect 141680 0 141736 400
rect 142128 0 142184 400
<< obsm2 >>
rect 686 149570 2154 149674
rect 2270 149570 3442 149674
rect 3558 149570 4730 149674
rect 4846 149570 6018 149674
rect 6134 149570 7306 149674
rect 7422 149570 8594 149674
rect 8710 149570 9882 149674
rect 9998 149570 11170 149674
rect 11286 149570 12458 149674
rect 12574 149570 13746 149674
rect 13862 149570 15034 149674
rect 15150 149570 16322 149674
rect 16438 149570 17610 149674
rect 17726 149570 18898 149674
rect 19014 149570 20186 149674
rect 20302 149570 21474 149674
rect 21590 149570 22762 149674
rect 22878 149570 24050 149674
rect 24166 149570 25338 149674
rect 25454 149570 26626 149674
rect 26742 149570 27914 149674
rect 28030 149570 29202 149674
rect 29318 149570 30490 149674
rect 30606 149570 31778 149674
rect 31894 149570 33066 149674
rect 33182 149570 34354 149674
rect 34470 149570 35642 149674
rect 35758 149570 36930 149674
rect 37046 149570 38218 149674
rect 38334 149570 39506 149674
rect 39622 149570 40794 149674
rect 40910 149570 42082 149674
rect 42198 149570 43370 149674
rect 43486 149570 44658 149674
rect 44774 149570 45946 149674
rect 46062 149570 47234 149674
rect 47350 149570 48522 149674
rect 48638 149570 49810 149674
rect 49926 149570 51098 149674
rect 51214 149570 52386 149674
rect 52502 149570 53674 149674
rect 53790 149570 54962 149674
rect 55078 149570 56250 149674
rect 56366 149570 57538 149674
rect 57654 149570 58826 149674
rect 58942 149570 60114 149674
rect 60230 149570 61402 149674
rect 61518 149570 62690 149674
rect 62806 149570 63978 149674
rect 64094 149570 65266 149674
rect 65382 149570 66554 149674
rect 66670 149570 67842 149674
rect 67958 149570 69130 149674
rect 69246 149570 70418 149674
rect 70534 149570 71706 149674
rect 71822 149570 72994 149674
rect 73110 149570 74282 149674
rect 74398 149570 75570 149674
rect 75686 149570 76858 149674
rect 76974 149570 78146 149674
rect 78262 149570 79434 149674
rect 79550 149570 80722 149674
rect 80838 149570 82010 149674
rect 82126 149570 83298 149674
rect 83414 149570 84586 149674
rect 84702 149570 85874 149674
rect 85990 149570 87162 149674
rect 87278 149570 88450 149674
rect 88566 149570 89738 149674
rect 89854 149570 91026 149674
rect 91142 149570 92314 149674
rect 92430 149570 93602 149674
rect 93718 149570 94890 149674
rect 95006 149570 96178 149674
rect 96294 149570 97466 149674
rect 97582 149570 98754 149674
rect 98870 149570 100042 149674
rect 100158 149570 101330 149674
rect 101446 149570 102618 149674
rect 102734 149570 103906 149674
rect 104022 149570 105194 149674
rect 105310 149570 106482 149674
rect 106598 149570 107770 149674
rect 107886 149570 109058 149674
rect 109174 149570 110346 149674
rect 110462 149570 111634 149674
rect 111750 149570 112922 149674
rect 113038 149570 114210 149674
rect 114326 149570 115498 149674
rect 115614 149570 116786 149674
rect 116902 149570 118074 149674
rect 118190 149570 119362 149674
rect 119478 149570 120650 149674
rect 120766 149570 121938 149674
rect 122054 149570 123226 149674
rect 123342 149570 124514 149674
rect 124630 149570 125802 149674
rect 125918 149570 127090 149674
rect 127206 149570 128378 149674
rect 128494 149570 129666 149674
rect 129782 149570 130954 149674
rect 131070 149570 132242 149674
rect 132358 149570 133530 149674
rect 133646 149570 134818 149674
rect 134934 149570 136106 149674
rect 136222 149570 137394 149674
rect 137510 149570 138682 149674
rect 138798 149570 139970 149674
rect 140086 149570 141258 149674
rect 141374 149570 142546 149674
rect 142662 149570 143834 149674
rect 143950 149570 145122 149674
rect 145238 149570 146410 149674
rect 146526 149570 147698 149674
rect 147814 149570 149338 149674
rect 686 430 149338 149570
rect 686 400 7698 430
rect 7814 400 8146 430
rect 8262 400 8594 430
rect 8710 400 9042 430
rect 9158 400 9490 430
rect 9606 400 9938 430
rect 10054 400 10386 430
rect 10502 400 10834 430
rect 10950 400 11282 430
rect 11398 400 11730 430
rect 11846 400 12178 430
rect 12294 400 12626 430
rect 12742 400 13074 430
rect 13190 400 13522 430
rect 13638 400 13970 430
rect 14086 400 14418 430
rect 14534 400 14866 430
rect 14982 400 15314 430
rect 15430 400 15762 430
rect 15878 400 16210 430
rect 16326 400 16658 430
rect 16774 400 17106 430
rect 17222 400 17554 430
rect 17670 400 18002 430
rect 18118 400 18450 430
rect 18566 400 18898 430
rect 19014 400 19346 430
rect 19462 400 19794 430
rect 19910 400 20242 430
rect 20358 400 20690 430
rect 20806 400 21138 430
rect 21254 400 21586 430
rect 21702 400 22034 430
rect 22150 400 22482 430
rect 22598 400 22930 430
rect 23046 400 23378 430
rect 23494 400 23826 430
rect 23942 400 24274 430
rect 24390 400 24722 430
rect 24838 400 25170 430
rect 25286 400 25618 430
rect 25734 400 26066 430
rect 26182 400 26514 430
rect 26630 400 26962 430
rect 27078 400 27410 430
rect 27526 400 27858 430
rect 27974 400 28306 430
rect 28422 400 28754 430
rect 28870 400 29202 430
rect 29318 400 29650 430
rect 29766 400 30098 430
rect 30214 400 30546 430
rect 30662 400 30994 430
rect 31110 400 31442 430
rect 31558 400 31890 430
rect 32006 400 32338 430
rect 32454 400 32786 430
rect 32902 400 33234 430
rect 33350 400 33682 430
rect 33798 400 34130 430
rect 34246 400 34578 430
rect 34694 400 35026 430
rect 35142 400 35474 430
rect 35590 400 35922 430
rect 36038 400 36370 430
rect 36486 400 36818 430
rect 36934 400 37266 430
rect 37382 400 37714 430
rect 37830 400 38162 430
rect 38278 400 38610 430
rect 38726 400 39058 430
rect 39174 400 39506 430
rect 39622 400 39954 430
rect 40070 400 40402 430
rect 40518 400 40850 430
rect 40966 400 41298 430
rect 41414 400 41746 430
rect 41862 400 42194 430
rect 42310 400 42642 430
rect 42758 400 43090 430
rect 43206 400 43538 430
rect 43654 400 43986 430
rect 44102 400 44434 430
rect 44550 400 44882 430
rect 44998 400 45330 430
rect 45446 400 45778 430
rect 45894 400 46226 430
rect 46342 400 46674 430
rect 46790 400 47122 430
rect 47238 400 47570 430
rect 47686 400 48018 430
rect 48134 400 48466 430
rect 48582 400 48914 430
rect 49030 400 49362 430
rect 49478 400 49810 430
rect 49926 400 50258 430
rect 50374 400 50706 430
rect 50822 400 51154 430
rect 51270 400 51602 430
rect 51718 400 52050 430
rect 52166 400 52498 430
rect 52614 400 52946 430
rect 53062 400 53394 430
rect 53510 400 53842 430
rect 53958 400 54290 430
rect 54406 400 54738 430
rect 54854 400 55186 430
rect 55302 400 55634 430
rect 55750 400 56082 430
rect 56198 400 56530 430
rect 56646 400 56978 430
rect 57094 400 57426 430
rect 57542 400 57874 430
rect 57990 400 58322 430
rect 58438 400 58770 430
rect 58886 400 59218 430
rect 59334 400 59666 430
rect 59782 400 60114 430
rect 60230 400 60562 430
rect 60678 400 61010 430
rect 61126 400 61458 430
rect 61574 400 61906 430
rect 62022 400 62354 430
rect 62470 400 62802 430
rect 62918 400 63250 430
rect 63366 400 63698 430
rect 63814 400 64146 430
rect 64262 400 64594 430
rect 64710 400 65042 430
rect 65158 400 65490 430
rect 65606 400 65938 430
rect 66054 400 66386 430
rect 66502 400 66834 430
rect 66950 400 67282 430
rect 67398 400 67730 430
rect 67846 400 68178 430
rect 68294 400 68626 430
rect 68742 400 69074 430
rect 69190 400 69522 430
rect 69638 400 69970 430
rect 70086 400 70418 430
rect 70534 400 70866 430
rect 70982 400 71314 430
rect 71430 400 71762 430
rect 71878 400 72210 430
rect 72326 400 72658 430
rect 72774 400 73106 430
rect 73222 400 73554 430
rect 73670 400 74002 430
rect 74118 400 74450 430
rect 74566 400 74898 430
rect 75014 400 75346 430
rect 75462 400 75794 430
rect 75910 400 76242 430
rect 76358 400 76690 430
rect 76806 400 77138 430
rect 77254 400 77586 430
rect 77702 400 78034 430
rect 78150 400 78482 430
rect 78598 400 78930 430
rect 79046 400 79378 430
rect 79494 400 79826 430
rect 79942 400 80274 430
rect 80390 400 80722 430
rect 80838 400 81170 430
rect 81286 400 81618 430
rect 81734 400 82066 430
rect 82182 400 82514 430
rect 82630 400 82962 430
rect 83078 400 83410 430
rect 83526 400 83858 430
rect 83974 400 84306 430
rect 84422 400 84754 430
rect 84870 400 85202 430
rect 85318 400 85650 430
rect 85766 400 86098 430
rect 86214 400 86546 430
rect 86662 400 86994 430
rect 87110 400 87442 430
rect 87558 400 87890 430
rect 88006 400 88338 430
rect 88454 400 88786 430
rect 88902 400 89234 430
rect 89350 400 89682 430
rect 89798 400 90130 430
rect 90246 400 90578 430
rect 90694 400 91026 430
rect 91142 400 91474 430
rect 91590 400 91922 430
rect 92038 400 92370 430
rect 92486 400 92818 430
rect 92934 400 93266 430
rect 93382 400 93714 430
rect 93830 400 94162 430
rect 94278 400 94610 430
rect 94726 400 95058 430
rect 95174 400 95506 430
rect 95622 400 95954 430
rect 96070 400 96402 430
rect 96518 400 96850 430
rect 96966 400 97298 430
rect 97414 400 97746 430
rect 97862 400 98194 430
rect 98310 400 98642 430
rect 98758 400 99090 430
rect 99206 400 99538 430
rect 99654 400 99986 430
rect 100102 400 100434 430
rect 100550 400 100882 430
rect 100998 400 101330 430
rect 101446 400 101778 430
rect 101894 400 102226 430
rect 102342 400 102674 430
rect 102790 400 103122 430
rect 103238 400 103570 430
rect 103686 400 104018 430
rect 104134 400 104466 430
rect 104582 400 104914 430
rect 105030 400 105362 430
rect 105478 400 105810 430
rect 105926 400 106258 430
rect 106374 400 106706 430
rect 106822 400 107154 430
rect 107270 400 107602 430
rect 107718 400 108050 430
rect 108166 400 108498 430
rect 108614 400 108946 430
rect 109062 400 109394 430
rect 109510 400 109842 430
rect 109958 400 110290 430
rect 110406 400 110738 430
rect 110854 400 111186 430
rect 111302 400 111634 430
rect 111750 400 112082 430
rect 112198 400 112530 430
rect 112646 400 112978 430
rect 113094 400 113426 430
rect 113542 400 113874 430
rect 113990 400 114322 430
rect 114438 400 114770 430
rect 114886 400 115218 430
rect 115334 400 115666 430
rect 115782 400 116114 430
rect 116230 400 116562 430
rect 116678 400 117010 430
rect 117126 400 117458 430
rect 117574 400 117906 430
rect 118022 400 118354 430
rect 118470 400 118802 430
rect 118918 400 119250 430
rect 119366 400 119698 430
rect 119814 400 120146 430
rect 120262 400 120594 430
rect 120710 400 121042 430
rect 121158 400 121490 430
rect 121606 400 121938 430
rect 122054 400 122386 430
rect 122502 400 122834 430
rect 122950 400 123282 430
rect 123398 400 123730 430
rect 123846 400 124178 430
rect 124294 400 124626 430
rect 124742 400 125074 430
rect 125190 400 125522 430
rect 125638 400 125970 430
rect 126086 400 126418 430
rect 126534 400 126866 430
rect 126982 400 127314 430
rect 127430 400 127762 430
rect 127878 400 128210 430
rect 128326 400 128658 430
rect 128774 400 129106 430
rect 129222 400 129554 430
rect 129670 400 130002 430
rect 130118 400 130450 430
rect 130566 400 130898 430
rect 131014 400 131346 430
rect 131462 400 131794 430
rect 131910 400 132242 430
rect 132358 400 132690 430
rect 132806 400 133138 430
rect 133254 400 133586 430
rect 133702 400 134034 430
rect 134150 400 134482 430
rect 134598 400 134930 430
rect 135046 400 135378 430
rect 135494 400 135826 430
rect 135942 400 136274 430
rect 136390 400 136722 430
rect 136838 400 137170 430
rect 137286 400 137618 430
rect 137734 400 138066 430
rect 138182 400 138514 430
rect 138630 400 138962 430
rect 139078 400 139410 430
rect 139526 400 139858 430
rect 139974 400 140306 430
rect 140422 400 140754 430
rect 140870 400 141202 430
rect 141318 400 141650 430
rect 141766 400 142098 430
rect 142214 400 149338 430
<< obsm3 >>
rect 681 1554 149343 148890
<< metal4 >>
rect 2224 1538 2384 148206
rect 9904 1538 10064 148206
rect 17584 1538 17744 148206
rect 25264 1538 25424 148206
rect 32944 1538 33104 148206
rect 40624 1538 40784 148206
rect 48304 1538 48464 148206
rect 55984 1538 56144 148206
rect 63664 1538 63824 148206
rect 71344 1538 71504 148206
rect 79024 1538 79184 148206
rect 86704 1538 86864 148206
rect 94384 1538 94544 148206
rect 102064 1538 102224 148206
rect 109744 1538 109904 148206
rect 117424 1538 117584 148206
rect 125104 1538 125264 148206
rect 132784 1538 132944 148206
rect 140464 1538 140624 148206
rect 148144 1538 148304 148206
<< obsm4 >>
rect 1974 148236 146986 148895
rect 1974 6449 2194 148236
rect 2414 6449 9874 148236
rect 10094 6449 17554 148236
rect 17774 6449 25234 148236
rect 25454 6449 32914 148236
rect 33134 6449 40594 148236
rect 40814 6449 48274 148236
rect 48494 6449 55954 148236
rect 56174 6449 63634 148236
rect 63854 6449 71314 148236
rect 71534 6449 78994 148236
rect 79214 6449 86674 148236
rect 86894 6449 94354 148236
rect 94574 6449 102034 148236
rect 102254 6449 109714 148236
rect 109934 6449 117394 148236
rect 117614 6449 125074 148236
rect 125294 6449 132754 148236
rect 132974 6449 140434 148236
rect 140654 6449 146986 148236
<< labels >>
rlabel metal2 s 2184 149600 2240 150000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 40824 149600 40880 150000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 44688 149600 44744 150000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 48552 149600 48608 150000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 52416 149600 52472 150000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 56280 149600 56336 150000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 60144 149600 60200 150000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 64008 149600 64064 150000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 67872 149600 67928 150000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 71736 149600 71792 150000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 75600 149600 75656 150000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 6048 149600 6104 150000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 79464 149600 79520 150000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 83328 149600 83384 150000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 87192 149600 87248 150000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 91056 149600 91112 150000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 94920 149600 94976 150000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 98784 149600 98840 150000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 102648 149600 102704 150000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 106512 149600 106568 150000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 110376 149600 110432 150000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 114240 149600 114296 150000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9912 149600 9968 150000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 118104 149600 118160 150000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 121968 149600 122024 150000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 125832 149600 125888 150000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 129696 149600 129752 150000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 133560 149600 133616 150000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 137424 149600 137480 150000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 141288 149600 141344 150000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 145152 149600 145208 150000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13776 149600 13832 150000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17640 149600 17696 150000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21504 149600 21560 150000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 25368 149600 25424 150000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 29232 149600 29288 150000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 33096 149600 33152 150000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 36960 149600 37016 150000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3472 149600 3528 150000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 42112 149600 42168 150000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 45976 149600 46032 150000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 49840 149600 49896 150000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 53704 149600 53760 150000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 57568 149600 57624 150000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 61432 149600 61488 150000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 65296 149600 65352 150000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 69160 149600 69216 150000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 73024 149600 73080 150000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 76888 149600 76944 150000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7336 149600 7392 150000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 80752 149600 80808 150000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 84616 149600 84672 150000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 88480 149600 88536 150000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 92344 149600 92400 150000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 96208 149600 96264 150000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 100072 149600 100128 150000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 103936 149600 103992 150000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 107800 149600 107856 150000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 111664 149600 111720 150000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 115528 149600 115584 150000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 11200 149600 11256 150000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 119392 149600 119448 150000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 123256 149600 123312 150000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 127120 149600 127176 150000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 130984 149600 131040 150000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 134848 149600 134904 150000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 138712 149600 138768 150000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 142576 149600 142632 150000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 146440 149600 146496 150000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 15064 149600 15120 150000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 18928 149600 18984 150000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 22792 149600 22848 150000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 26656 149600 26712 150000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 30520 149600 30576 150000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 34384 149600 34440 150000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 38248 149600 38304 150000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4760 149600 4816 150000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 43400 149600 43456 150000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 47264 149600 47320 150000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 51128 149600 51184 150000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 54992 149600 55048 150000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 58856 149600 58912 150000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 62720 149600 62776 150000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 66584 149600 66640 150000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 70448 149600 70504 150000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 74312 149600 74368 150000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 78176 149600 78232 150000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 8624 149600 8680 150000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 82040 149600 82096 150000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 85904 149600 85960 150000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 89768 149600 89824 150000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 93632 149600 93688 150000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 97496 149600 97552 150000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 101360 149600 101416 150000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 105224 149600 105280 150000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 109088 149600 109144 150000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 112952 149600 113008 150000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 116816 149600 116872 150000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 12488 149600 12544 150000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 120680 149600 120736 150000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 124544 149600 124600 150000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 128408 149600 128464 150000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 132272 149600 132328 150000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 136136 149600 136192 150000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 140000 149600 140056 150000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 143864 149600 143920 150000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 147728 149600 147784 150000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16352 149600 16408 150000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20216 149600 20272 150000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24080 149600 24136 150000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 27944 149600 28000 150000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 31808 149600 31864 150000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 35672 149600 35728 150000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 39536 149600 39592 150000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 141232 0 141288 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 141680 0 141736 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 142128 0 142184 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 55216 0 55272 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 68656 0 68712 400 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 70000 0 70056 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 71344 0 71400 400 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 72688 0 72744 400 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 75376 0 75432 400 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 76720 0 76776 400 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 78064 0 78120 400 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 80752 0 80808 400 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 56560 0 56616 400 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 84784 0 84840 400 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 86128 0 86184 400 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 87472 0 87528 400 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 88816 0 88872 400 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 90160 0 90216 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 91504 0 91560 400 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 92848 0 92904 400 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 94192 0 94248 400 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 95536 0 95592 400 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 96880 0 96936 400 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 98224 0 98280 400 6 la_data_in[32]
port 143 nsew signal input
rlabel metal2 s 99568 0 99624 400 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 100912 0 100968 400 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 102256 0 102312 400 6 la_data_in[35]
port 146 nsew signal input
rlabel metal2 s 103600 0 103656 400 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 104944 0 105000 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 106288 0 106344 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal2 s 107632 0 107688 400 6 la_data_in[39]
port 150 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 la_data_in[3]
port 151 nsew signal input
rlabel metal2 s 108976 0 109032 400 6 la_data_in[40]
port 152 nsew signal input
rlabel metal2 s 110320 0 110376 400 6 la_data_in[41]
port 153 nsew signal input
rlabel metal2 s 111664 0 111720 400 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 113008 0 113064 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 114352 0 114408 400 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 115696 0 115752 400 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 117040 0 117096 400 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 118384 0 118440 400 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 119728 0 119784 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal2 s 121072 0 121128 400 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 60592 0 60648 400 6 la_data_in[4]
port 162 nsew signal input
rlabel metal2 s 122416 0 122472 400 6 la_data_in[50]
port 163 nsew signal input
rlabel metal2 s 123760 0 123816 400 6 la_data_in[51]
port 164 nsew signal input
rlabel metal2 s 125104 0 125160 400 6 la_data_in[52]
port 165 nsew signal input
rlabel metal2 s 126448 0 126504 400 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 127792 0 127848 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal2 s 129136 0 129192 400 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 130480 0 130536 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 131824 0 131880 400 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 133168 0 133224 400 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 134512 0 134568 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal2 s 61936 0 61992 400 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 135856 0 135912 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal2 s 137200 0 137256 400 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 138544 0 138600 400 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 la_data_in[6]
port 178 nsew signal input
rlabel metal2 s 64624 0 64680 400 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal2 s 67312 0 67368 400 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 la_data_out[0]
port 182 nsew signal output
rlabel metal2 s 69104 0 69160 400 6 la_data_out[10]
port 183 nsew signal output
rlabel metal2 s 70448 0 70504 400 6 la_data_out[11]
port 184 nsew signal output
rlabel metal2 s 71792 0 71848 400 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 73136 0 73192 400 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 74480 0 74536 400 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 75824 0 75880 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 78512 0 78568 400 6 la_data_out[17]
port 190 nsew signal output
rlabel metal2 s 79856 0 79912 400 6 la_data_out[18]
port 191 nsew signal output
rlabel metal2 s 81200 0 81256 400 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 57008 0 57064 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal2 s 82544 0 82600 400 6 la_data_out[20]
port 194 nsew signal output
rlabel metal2 s 83888 0 83944 400 6 la_data_out[21]
port 195 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 86576 0 86632 400 6 la_data_out[23]
port 197 nsew signal output
rlabel metal2 s 87920 0 87976 400 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 89264 0 89320 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal2 s 90608 0 90664 400 6 la_data_out[26]
port 200 nsew signal output
rlabel metal2 s 91952 0 92008 400 6 la_data_out[27]
port 201 nsew signal output
rlabel metal2 s 93296 0 93352 400 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 94640 0 94696 400 6 la_data_out[29]
port 203 nsew signal output
rlabel metal2 s 58352 0 58408 400 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 95984 0 96040 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 97328 0 97384 400 6 la_data_out[31]
port 206 nsew signal output
rlabel metal2 s 98672 0 98728 400 6 la_data_out[32]
port 207 nsew signal output
rlabel metal2 s 100016 0 100072 400 6 la_data_out[33]
port 208 nsew signal output
rlabel metal2 s 101360 0 101416 400 6 la_data_out[34]
port 209 nsew signal output
rlabel metal2 s 102704 0 102760 400 6 la_data_out[35]
port 210 nsew signal output
rlabel metal2 s 104048 0 104104 400 6 la_data_out[36]
port 211 nsew signal output
rlabel metal2 s 105392 0 105448 400 6 la_data_out[37]
port 212 nsew signal output
rlabel metal2 s 106736 0 106792 400 6 la_data_out[38]
port 213 nsew signal output
rlabel metal2 s 108080 0 108136 400 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 59696 0 59752 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 109424 0 109480 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 110768 0 110824 400 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 112112 0 112168 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal2 s 113456 0 113512 400 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 114800 0 114856 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 116144 0 116200 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 117488 0 117544 400 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 118832 0 118888 400 6 la_data_out[47]
port 223 nsew signal output
rlabel metal2 s 120176 0 120232 400 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 121520 0 121576 400 6 la_data_out[49]
port 225 nsew signal output
rlabel metal2 s 61040 0 61096 400 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 122864 0 122920 400 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 124208 0 124264 400 6 la_data_out[51]
port 228 nsew signal output
rlabel metal2 s 125552 0 125608 400 6 la_data_out[52]
port 229 nsew signal output
rlabel metal2 s 126896 0 126952 400 6 la_data_out[53]
port 230 nsew signal output
rlabel metal2 s 128240 0 128296 400 6 la_data_out[54]
port 231 nsew signal output
rlabel metal2 s 129584 0 129640 400 6 la_data_out[55]
port 232 nsew signal output
rlabel metal2 s 130928 0 130984 400 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 132272 0 132328 400 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 133616 0 133672 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 134960 0 135016 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal2 s 62384 0 62440 400 6 la_data_out[5]
port 237 nsew signal output
rlabel metal2 s 136304 0 136360 400 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 137648 0 137704 400 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 138992 0 139048 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal2 s 140336 0 140392 400 6 la_data_out[63]
port 241 nsew signal output
rlabel metal2 s 63728 0 63784 400 6 la_data_out[6]
port 242 nsew signal output
rlabel metal2 s 65072 0 65128 400 6 la_data_out[7]
port 243 nsew signal output
rlabel metal2 s 66416 0 66472 400 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 67760 0 67816 400 6 la_data_out[9]
port 245 nsew signal output
rlabel metal2 s 56112 0 56168 400 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 70896 0 70952 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 72240 0 72296 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 la_oenb[14]
port 251 nsew signal input
rlabel metal2 s 76272 0 76328 400 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 77616 0 77672 400 6 la_oenb[16]
port 253 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 80304 0 80360 400 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal2 s 82992 0 83048 400 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 84336 0 84392 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal2 s 85680 0 85736 400 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 87024 0 87080 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal2 s 88368 0 88424 400 6 la_oenb[24]
port 262 nsew signal input
rlabel metal2 s 89712 0 89768 400 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 91056 0 91112 400 6 la_oenb[26]
port 264 nsew signal input
rlabel metal2 s 92400 0 92456 400 6 la_oenb[27]
port 265 nsew signal input
rlabel metal2 s 93744 0 93800 400 6 la_oenb[28]
port 266 nsew signal input
rlabel metal2 s 95088 0 95144 400 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 96432 0 96488 400 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 97776 0 97832 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 99120 0 99176 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 100464 0 100520 400 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 101808 0 101864 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal2 s 103152 0 103208 400 6 la_oenb[35]
port 274 nsew signal input
rlabel metal2 s 104496 0 104552 400 6 la_oenb[36]
port 275 nsew signal input
rlabel metal2 s 105840 0 105896 400 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 107184 0 107240 400 6 la_oenb[38]
port 277 nsew signal input
rlabel metal2 s 108528 0 108584 400 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 60144 0 60200 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 109872 0 109928 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal2 s 111216 0 111272 400 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 112560 0 112616 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 113904 0 113960 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal2 s 115248 0 115304 400 6 la_oenb[44]
port 284 nsew signal input
rlabel metal2 s 116592 0 116648 400 6 la_oenb[45]
port 285 nsew signal input
rlabel metal2 s 117936 0 117992 400 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 119280 0 119336 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 120624 0 120680 400 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 121968 0 122024 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal2 s 61488 0 61544 400 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 123312 0 123368 400 6 la_oenb[50]
port 291 nsew signal input
rlabel metal2 s 124656 0 124712 400 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 126000 0 126056 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 127344 0 127400 400 6 la_oenb[53]
port 294 nsew signal input
rlabel metal2 s 128688 0 128744 400 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 130032 0 130088 400 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 131376 0 131432 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal2 s 132720 0 132776 400 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 134064 0 134120 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_oenb[59]
port 300 nsew signal input
rlabel metal2 s 62832 0 62888 400 6 la_oenb[5]
port 301 nsew signal input
rlabel metal2 s 136752 0 136808 400 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 138096 0 138152 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 139440 0 139496 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal2 s 140784 0 140840 400 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 64176 0 64232 400 6 la_oenb[6]
port 306 nsew signal input
rlabel metal2 s 65520 0 65576 400 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 66864 0 66920 400 6 la_oenb[8]
port 308 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 2224 1538 2384 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 148206 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 148206 6 vss
port 311 nsew ground bidirectional
rlabel metal2 s 7728 0 7784 400 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wb_rst_i
port 313 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 37744 0 37800 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 40432 0 40488 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal2 s 51184 0 51240 400 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal2 s 53872 0 53928 400 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 38192 0 38248 400 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 27888 0 27944 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal2 s 29232 0 29288 400 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 30576 0 30632 400 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal2 s 31920 0 31976 400 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 33264 0 33320 400 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal2 s 35952 0 36008 400 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 37296 0 37352 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal2 s 44016 0 44072 400 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 46704 0 46760 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 49392 0 49448 400 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 50736 0 50792 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal2 s 53424 0 53480 400 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 22512 0 22568 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 23856 0 23912 400 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 25200 0 25256 400 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wbs_stb_i
port 416 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 150000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 62449974
string GDS_FILE /home/wenting/caravel_user_project/openlane/vb_wrapper/runs/22_12_05_20_12/results/signoff/vb_wrapper.magic.gds
string GDS_START 404270
<< end >>

