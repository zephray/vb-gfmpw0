magic
tech gf180mcuC
magscale 1 10
timestamp 1670290910
<< metal1 >>
rect 324258 198270 324270 198322
rect 324322 198319 324334 198322
rect 325042 198319 325054 198322
rect 324322 198273 325054 198319
rect 324322 198270 324334 198273
rect 325042 198270 325054 198273
rect 325106 198270 325118 198322
<< via1 >>
rect 324270 198270 324322 198322
rect 325054 198270 325106 198322
<< metal2 >>
rect 10108 595644 10948 595700
rect 11032 595672 11256 597000
rect 9212 520884 9268 520894
rect 4172 516628 4228 516638
rect 4172 503188 4228 516572
rect 4172 503122 4228 503132
rect 5852 502516 5908 502526
rect 5852 501508 5908 502460
rect 5852 501442 5908 501452
rect 9212 206388 9268 520828
rect 10108 503300 10164 595644
rect 10892 595476 10948 595644
rect 11004 595560 11256 595672
rect 31948 595644 33012 595700
rect 33096 595672 33320 597000
rect 11004 595476 11060 595560
rect 10892 595420 11060 595476
rect 14252 586404 14308 586414
rect 14252 565348 14308 586348
rect 31948 583828 32004 595644
rect 32956 595476 33012 595644
rect 33068 595560 33320 595672
rect 55160 595672 55384 597000
rect 55160 595560 55412 595672
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 99260 595560 99512 595672
rect 121324 595560 121576 595672
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 143416 595560 143668 595672
rect 165480 595560 165732 595672
rect 187544 595560 187796 595672
rect 33068 595476 33124 595560
rect 32956 595420 33124 595476
rect 55356 593124 55412 595560
rect 55356 593058 55412 593068
rect 31948 583762 32004 583772
rect 14252 565282 14308 565292
rect 27692 530964 27748 530974
rect 10108 503234 10164 503244
rect 12572 527604 12628 527614
rect 12572 275604 12628 527548
rect 22652 519204 22708 519214
rect 19292 514164 19348 514174
rect 12572 275538 12628 275548
rect 14252 510804 14308 510814
rect 14252 262164 14308 510748
rect 17612 504084 17668 504094
rect 15932 499044 15988 499054
rect 15932 458724 15988 498988
rect 17612 473844 17668 504028
rect 17612 473778 17668 473788
rect 15932 458658 15988 458668
rect 19292 317604 19348 514108
rect 22652 361284 22708 519148
rect 22652 361218 22708 361228
rect 19292 317538 19348 317548
rect 14252 262098 14308 262108
rect 9212 206322 9268 206332
rect 10108 195748 10164 195758
rect 4172 94948 4228 94958
rect 4172 93492 4228 94892
rect 4172 93426 4228 93436
rect 4172 41188 4228 41198
rect 4172 36932 4228 41132
rect 4172 36866 4228 36876
rect 4284 27748 4340 27758
rect 4172 26068 4228 26078
rect 4172 8820 4228 26012
rect 4284 22932 4340 27692
rect 4284 22866 4340 22876
rect 4172 8754 4228 8764
rect 10108 420 10164 195692
rect 22652 192388 22708 192398
rect 11788 31108 11844 31118
rect 11228 480 11396 532
rect 11228 476 11592 480
rect 11228 420 11284 476
rect 10108 364 11284 420
rect 11340 392 11592 476
rect 11368 -960 11592 392
rect 11788 420 11844 31052
rect 18508 12628 18564 12638
rect 17276 6244 17332 6254
rect 15372 5012 15428 5022
rect 13132 480 13300 532
rect 15372 480 15428 4956
rect 17276 480 17332 6188
rect 13132 476 13496 480
rect 13132 420 13188 476
rect 11788 364 13188 420
rect 13244 392 13496 476
rect 13272 -960 13496 392
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18508 420 18564 12572
rect 22652 5012 22708 192332
rect 27692 191604 27748 530908
rect 77308 526708 77364 595560
rect 99260 572908 99316 595560
rect 121324 572908 121380 595560
rect 143612 585508 143668 595560
rect 165676 590212 165732 595560
rect 187740 593236 187796 595560
rect 187740 593170 187796 593180
rect 208348 595644 209524 595700
rect 209608 595672 209832 597000
rect 165676 590146 165732 590156
rect 167132 590212 167188 590222
rect 143612 585442 143668 585452
rect 99148 572852 99316 572908
rect 120988 572852 121380 572908
rect 99148 550228 99204 572852
rect 99148 550162 99204 550172
rect 77308 526642 77364 526652
rect 120988 525140 121044 572852
rect 167132 551908 167188 590156
rect 167132 551842 167188 551852
rect 120988 525074 121044 525084
rect 206668 529396 206724 529406
rect 44492 522564 44548 522574
rect 44492 233604 44548 522508
rect 203308 520996 203364 521006
rect 158732 517748 158788 517758
rect 155372 517636 155428 517646
rect 98252 507556 98308 507566
rect 98252 487284 98308 507500
rect 98252 487218 98308 487228
rect 44492 233538 44548 233548
rect 144508 199220 144564 199230
rect 65548 199108 65604 199118
rect 57036 195860 57092 195870
rect 27692 191538 27748 191548
rect 29372 194068 29428 194078
rect 27692 190708 27748 190718
rect 22652 4946 22708 4956
rect 24892 9268 24948 9278
rect 22988 4340 23044 4350
rect 21084 4116 21140 4126
rect 18844 480 19012 532
rect 21084 480 21140 4060
rect 22988 480 23044 4284
rect 24892 480 24948 9212
rect 27692 4340 27748 190652
rect 27692 4274 27748 4284
rect 28700 4340 28756 4350
rect 26796 4228 26852 4238
rect 26796 480 26852 4172
rect 28700 480 28756 4284
rect 29372 4228 29428 194012
rect 36988 189140 37044 189150
rect 31948 189028 32004 189038
rect 30268 44548 30324 44558
rect 30268 20188 30324 44492
rect 30268 20132 30436 20188
rect 29372 4162 29428 4172
rect 18844 476 19208 480
rect 18844 420 18900 476
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18508 364 18900 420
rect 18956 392 19208 476
rect 18984 -960 19208 392
rect 20888 392 21140 480
rect 22792 392 23044 480
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30380 480 30436 20132
rect 30380 392 30632 480
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 31948 420 32004 188972
rect 33628 14308 33684 14318
rect 32172 480 32340 532
rect 32172 476 32536 480
rect 32172 420 32228 476
rect 31948 364 32228 420
rect 32284 392 32536 476
rect 32312 -960 32536 392
rect 33628 420 33684 14252
rect 36316 4452 36372 4462
rect 34076 480 34244 532
rect 36316 480 36372 4396
rect 34076 476 34440 480
rect 34076 420 34132 476
rect 33628 364 34132 420
rect 34188 392 34440 476
rect 34216 -960 34440 392
rect 36120 392 36372 480
rect 36988 420 37044 189084
rect 45388 187348 45444 187358
rect 41132 178948 41188 178958
rect 40124 4116 40180 4126
rect 37884 480 38052 532
rect 40124 480 40180 4060
rect 41132 4116 41188 178892
rect 44492 56308 44548 56318
rect 41132 4050 41188 4060
rect 41916 5012 41972 5022
rect 41916 480 41972 4956
rect 44492 5012 44548 56252
rect 45388 20188 45444 187292
rect 47068 180628 47124 180638
rect 45388 20132 45668 20188
rect 44492 4946 44548 4956
rect 43932 4564 43988 4574
rect 43932 480 43988 4508
rect 37884 476 38248 480
rect 37884 420 37940 476
rect 36120 -960 36344 392
rect 36988 364 37940 420
rect 37996 392 38248 476
rect 38024 -960 38248 392
rect 39928 392 40180 480
rect 39928 -960 40152 392
rect 41832 -960 42056 480
rect 43736 392 43988 480
rect 45612 480 45668 20132
rect 45612 392 45864 480
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47068 420 47124 180572
rect 52108 160468 52164 160478
rect 48748 52948 48804 52958
rect 47404 480 47572 532
rect 47404 476 47768 480
rect 47404 420 47460 476
rect 47068 364 47460 420
rect 47516 392 47768 476
rect 47544 -960 47768 392
rect 48748 420 48804 52892
rect 51548 4676 51604 4686
rect 49308 480 49476 532
rect 51548 480 51604 4620
rect 49308 476 49672 480
rect 49308 420 49364 476
rect 48748 364 49364 420
rect 49420 392 49672 476
rect 49448 -960 49672 392
rect 51352 392 51604 480
rect 52108 420 52164 160412
rect 53788 54628 53844 54638
rect 53116 480 53284 532
rect 53116 476 53480 480
rect 53116 420 53172 476
rect 51352 -960 51576 392
rect 52108 364 53172 420
rect 53228 392 53480 476
rect 53256 -960 53480 392
rect 53788 420 53844 54572
rect 57036 4788 57092 195804
rect 62972 165508 63028 165518
rect 58828 158788 58884 158798
rect 58828 20188 58884 158732
rect 58828 20132 58996 20188
rect 57036 4732 57204 4788
rect 55020 480 55188 532
rect 57148 480 57204 4732
rect 58940 480 58996 20132
rect 62860 4788 62916 4798
rect 61068 4116 61124 4126
rect 61068 480 61124 4060
rect 62860 480 62916 4732
rect 62972 4116 63028 165452
rect 62972 4050 63028 4060
rect 63868 157108 63924 157118
rect 55020 476 55384 480
rect 55020 420 55076 476
rect 53788 364 55076 420
rect 55132 392 55384 476
rect 55160 -960 55384 392
rect 57064 -960 57288 480
rect 58940 392 59192 480
rect 58968 -960 59192 392
rect 60872 392 61124 480
rect 60872 -960 61096 392
rect 62776 -960 63000 480
rect 63868 420 63924 157052
rect 64540 480 64708 532
rect 64540 476 64904 480
rect 64540 420 64596 476
rect 63868 364 64596 420
rect 64652 392 64904 476
rect 64680 -960 64904 392
rect 65548 420 65604 199052
rect 113372 197540 113428 197550
rect 94892 197428 94948 197438
rect 80668 185668 80724 185678
rect 72268 182308 72324 182318
rect 71372 167188 71428 167198
rect 68012 61348 68068 61358
rect 68012 4788 68068 61292
rect 68012 4722 68068 4732
rect 68908 37828 68964 37838
rect 68684 4116 68740 4126
rect 66444 480 66612 532
rect 68684 480 68740 4060
rect 66444 476 66808 480
rect 66444 420 66500 476
rect 65548 364 66500 420
rect 66556 392 66808 476
rect 66584 -960 66808 392
rect 68488 392 68740 480
rect 68908 420 68964 37772
rect 71372 4116 71428 167132
rect 71372 4050 71428 4060
rect 70252 480 70420 532
rect 72268 480 72324 182252
rect 75628 155428 75684 155438
rect 74396 4116 74452 4126
rect 74396 480 74452 4060
rect 70252 476 70616 480
rect 70252 420 70308 476
rect 68488 -960 68712 392
rect 68908 364 70308 420
rect 70364 392 70616 476
rect 72268 392 72520 480
rect 70392 -960 70616 392
rect 72296 -960 72520 392
rect 74200 392 74452 480
rect 75628 420 75684 155372
rect 78092 66388 78148 66398
rect 78092 4116 78148 66332
rect 78092 4050 78148 4060
rect 78204 7588 78260 7598
rect 75964 480 76132 532
rect 78204 480 78260 7532
rect 80108 4116 80164 4126
rect 80108 480 80164 4060
rect 75964 476 76328 480
rect 75964 420 76020 476
rect 74200 -960 74424 392
rect 75628 364 76020 420
rect 76076 392 76328 476
rect 76104 -960 76328 392
rect 78008 392 78260 480
rect 79912 392 80164 480
rect 80668 420 80724 185612
rect 89068 183988 89124 183998
rect 87388 175588 87444 175598
rect 84812 147028 84868 147038
rect 82348 17668 82404 17678
rect 81676 480 81844 532
rect 81676 476 82040 480
rect 81676 420 81732 476
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 80668 364 81732 420
rect 81788 392 82040 476
rect 81816 -960 82040 392
rect 82348 420 82404 17612
rect 84812 4116 84868 146972
rect 87388 20188 87444 175532
rect 87388 20132 87556 20188
rect 84812 4050 84868 4060
rect 85820 4788 85876 4798
rect 83580 480 83748 532
rect 85820 480 85876 4732
rect 83580 476 83944 480
rect 83580 420 83636 476
rect 82348 364 83636 420
rect 83692 392 83944 476
rect 83720 -960 83944 392
rect 85624 392 85876 480
rect 87500 480 87556 20132
rect 87500 392 87752 480
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89068 420 89124 183932
rect 90748 32900 90804 32910
rect 89292 480 89460 532
rect 89292 476 89656 480
rect 89292 420 89348 476
rect 89068 364 89348 420
rect 89404 392 89656 476
rect 89432 -960 89656 392
rect 90748 420 90804 32844
rect 93436 5124 93492 5134
rect 91196 480 91364 532
rect 93436 480 93492 5068
rect 94892 5124 94948 197372
rect 104188 194180 104244 194190
rect 97468 192500 97524 192510
rect 94892 5058 94948 5068
rect 95340 6020 95396 6030
rect 95340 480 95396 5964
rect 97244 4116 97300 4126
rect 97244 480 97300 4060
rect 91196 476 91560 480
rect 91196 420 91252 476
rect 90748 364 91252 420
rect 91308 392 91560 476
rect 91336 -960 91560 392
rect 93240 392 93492 480
rect 95144 392 95396 480
rect 97048 392 97300 480
rect 97468 420 97524 192444
rect 99932 185780 99988 185790
rect 99932 4116 99988 185724
rect 99932 4050 99988 4060
rect 100828 153748 100884 153758
rect 98812 480 98980 532
rect 100828 480 100884 153692
rect 102956 10948 103012 10958
rect 102956 480 103012 10892
rect 98812 476 99176 480
rect 98812 420 98868 476
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 97468 364 98868 420
rect 98924 392 99176 476
rect 100828 392 101080 480
rect 98952 -960 99176 392
rect 100856 -960 101080 392
rect 102760 392 103012 480
rect 104188 420 104244 194124
rect 105868 184100 105924 184110
rect 104524 480 104692 532
rect 104524 476 104888 480
rect 104524 420 104580 476
rect 102760 -960 102984 392
rect 104188 364 104580 420
rect 104636 392 104888 476
rect 104664 -960 104888 392
rect 105868 420 105924 184044
rect 109228 173908 109284 173918
rect 107548 148708 107604 148718
rect 106428 480 106596 532
rect 106428 476 106792 480
rect 106428 420 106484 476
rect 105868 364 106484 420
rect 106540 392 106792 476
rect 106568 -960 106792 392
rect 107548 420 107604 148652
rect 108332 480 108500 532
rect 108332 476 108696 480
rect 108332 420 108388 476
rect 107548 364 108388 420
rect 108444 392 108696 476
rect 108472 -960 108696 392
rect 109228 420 109284 173852
rect 113372 12628 113428 197484
rect 132636 195972 132692 195982
rect 117628 182420 117684 182430
rect 115948 172228 116004 172238
rect 113372 12562 113428 12572
rect 113484 24388 113540 24398
rect 112476 4116 112532 4126
rect 110236 480 110404 532
rect 112476 480 112532 4060
rect 113484 4116 113540 24332
rect 115948 20188 116004 172172
rect 115948 20132 116116 20188
rect 113484 4050 113540 4060
rect 114380 2548 114436 2558
rect 114380 480 114436 2492
rect 110236 476 110600 480
rect 110236 420 110292 476
rect 109228 364 110292 420
rect 110348 392 110600 476
rect 110376 -960 110600 392
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116060 480 116116 20132
rect 116060 392 116312 480
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117628 420 117684 182364
rect 120988 170548 121044 170558
rect 119308 42980 119364 42990
rect 117852 480 118020 532
rect 117852 476 118216 480
rect 117852 420 117908 476
rect 117628 364 117908 420
rect 117964 392 118216 476
rect 117992 -960 118216 392
rect 119308 420 119364 42924
rect 119756 480 119924 532
rect 119756 476 120120 480
rect 119756 420 119812 476
rect 119308 364 119812 420
rect 119868 392 120120 476
rect 119896 -960 120120 392
rect 120988 420 121044 170492
rect 126028 168868 126084 168878
rect 124348 19348 124404 19358
rect 122668 15988 122724 15998
rect 121660 480 121828 532
rect 121660 476 122024 480
rect 121660 420 121716 476
rect 120988 364 121716 420
rect 121772 392 122024 476
rect 121800 -960 122024 392
rect 122668 420 122724 15932
rect 123564 480 123732 532
rect 123564 476 123928 480
rect 123564 420 123620 476
rect 122668 364 123620 420
rect 123676 392 123928 476
rect 123704 -960 123928 392
rect 124348 420 124404 19292
rect 125468 480 125636 532
rect 125468 476 125832 480
rect 125468 420 125524 476
rect 124348 364 125524 420
rect 125580 392 125832 476
rect 125608 -960 125832 392
rect 126028 420 126084 168812
rect 129276 152068 129332 152078
rect 129276 4228 129332 152012
rect 131068 21028 131124 21038
rect 131068 20188 131124 20972
rect 131068 20132 131348 20188
rect 129276 4172 129444 4228
rect 127372 480 127540 532
rect 129388 480 129444 4172
rect 131292 480 131348 20132
rect 132636 4228 132692 195916
rect 137788 194292 137844 194302
rect 134428 187460 134484 187470
rect 132636 4172 132804 4228
rect 127372 476 127736 480
rect 127372 420 127428 476
rect 126028 364 127428 420
rect 127484 392 127736 476
rect 129388 392 129640 480
rect 131292 392 131544 480
rect 127512 -960 127736 392
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 132748 420 132804 4172
rect 133084 480 133252 532
rect 133084 476 133448 480
rect 133084 420 133140 476
rect 132748 364 133140 420
rect 133196 392 133448 476
rect 133224 -960 133448 392
rect 134428 420 134484 187404
rect 136108 177268 136164 177278
rect 134988 480 135156 532
rect 134988 476 135352 480
rect 134988 420 135044 476
rect 134428 364 135044 420
rect 135100 392 135352 476
rect 135128 -960 135352 392
rect 136108 420 136164 177212
rect 136892 480 137060 532
rect 136892 476 137256 480
rect 136892 420 136948 476
rect 136108 364 136948 420
rect 137004 392 137256 476
rect 137032 -960 137256 392
rect 137788 420 137844 194236
rect 139468 182532 139524 182542
rect 138796 480 138964 532
rect 138796 476 139160 480
rect 138796 420 138852 476
rect 137788 364 138852 420
rect 138908 392 139160 476
rect 138936 -960 139160 392
rect 139468 420 139524 182476
rect 142828 179060 142884 179070
rect 142716 174020 142772 174030
rect 142716 4116 142772 173964
rect 142716 4050 142772 4060
rect 140700 480 140868 532
rect 142828 480 142884 179004
rect 144508 20188 144564 199164
rect 154476 190820 154532 190830
rect 149436 167300 149492 167310
rect 144508 20132 144676 20188
rect 144620 480 144676 20132
rect 147868 17780 147924 17790
rect 146524 4116 146580 4126
rect 146524 480 146580 4060
rect 140700 476 141064 480
rect 140700 420 140756 476
rect 139468 364 140756 420
rect 140812 392 141064 476
rect 140840 -960 141064 392
rect 142744 -960 142968 480
rect 144620 392 144872 480
rect 146524 392 146776 480
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 147868 420 147924 17724
rect 149436 5012 149492 167244
rect 151228 29428 151284 29438
rect 149436 4946 149492 4956
rect 150332 5012 150388 5022
rect 148316 480 148484 532
rect 150332 480 150388 4956
rect 148316 476 148680 480
rect 148316 420 148372 476
rect 147868 364 148372 420
rect 148428 392 148680 476
rect 150332 392 150584 480
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 151228 420 151284 29372
rect 154364 9380 154420 9390
rect 152124 480 152292 532
rect 154364 480 154420 9324
rect 154476 4116 154532 190764
rect 155372 63924 155428 517580
rect 157052 515956 157108 515966
rect 157052 105924 157108 515900
rect 157052 105858 157108 105868
rect 157948 150388 158004 150398
rect 155372 63858 155428 63868
rect 154476 4050 154532 4060
rect 156044 4116 156100 4126
rect 152124 476 152488 480
rect 152124 420 152180 476
rect 151228 364 152180 420
rect 152236 392 152488 476
rect 152264 -960 152488 392
rect 154168 392 154420 480
rect 156044 480 156100 4060
rect 157948 480 158004 150332
rect 158732 149604 158788 517692
rect 163772 516180 163828 516190
rect 163772 403284 163828 516124
rect 185612 514388 185668 514398
rect 173852 512484 173908 512494
rect 167132 509460 167188 509470
rect 167132 445284 167188 509404
rect 167132 445218 167188 445228
rect 170492 507444 170548 507454
rect 163772 403218 163828 403228
rect 162988 180740 163044 180750
rect 158732 149538 158788 149548
rect 161308 165620 161364 165630
rect 159852 12628 159908 12638
rect 159852 480 159908 12572
rect 156044 392 156296 480
rect 157948 392 158200 480
rect 159852 392 160104 480
rect 154168 -960 154392 392
rect 156072 -960 156296 392
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161308 420 161364 165564
rect 161644 480 161812 532
rect 161644 476 162008 480
rect 161644 420 161700 476
rect 161308 364 161700 420
rect 161756 392 162008 476
rect 161784 -960 162008 392
rect 162988 420 163044 180684
rect 166348 162148 166404 162158
rect 165788 7700 165844 7710
rect 163548 480 163716 532
rect 165788 480 165844 7644
rect 163548 476 163912 480
rect 163548 420 163604 476
rect 162988 364 163604 420
rect 163660 392 163912 476
rect 163688 -960 163912 392
rect 165592 392 165844 480
rect 166348 420 166404 162092
rect 170492 50484 170548 507388
rect 173068 135268 173124 135278
rect 170492 50418 170548 50428
rect 171388 93268 171444 93278
rect 170492 49588 170548 49598
rect 169596 4116 169652 4126
rect 167356 480 167524 532
rect 169596 480 169652 4060
rect 170492 4116 170548 49532
rect 170492 4050 170548 4060
rect 171388 480 171444 93212
rect 173068 20188 173124 135212
rect 173852 134484 173908 512428
rect 178892 507780 178948 507790
rect 178108 189252 178164 189262
rect 173852 134418 173908 134428
rect 174748 177380 174804 177390
rect 173068 20132 173236 20188
rect 173180 480 173236 20132
rect 167356 476 167720 480
rect 167356 420 167412 476
rect 165592 -960 165816 392
rect 166348 364 167412 420
rect 167468 392 167720 476
rect 167496 -960 167720 392
rect 169400 392 169652 480
rect 169400 -960 169624 392
rect 171304 -960 171528 480
rect 173180 392 173432 480
rect 173208 -960 173432 392
rect 174748 420 174804 177324
rect 176428 22708 176484 22718
rect 174972 480 175140 532
rect 174972 476 175336 480
rect 174972 420 175028 476
rect 174748 364 175028 420
rect 175084 392 175336 476
rect 175112 -960 175336 392
rect 176428 420 176484 22652
rect 176876 480 177044 532
rect 176876 476 177240 480
rect 176876 420 176932 476
rect 176428 364 176932 420
rect 176988 392 177240 476
rect 177016 -960 177240 392
rect 178108 420 178164 189196
rect 178892 176484 178948 507724
rect 182252 506100 182308 506110
rect 180572 505988 180628 505998
rect 180572 346164 180628 505932
rect 182252 388164 182308 506044
rect 182252 388098 182308 388108
rect 180572 346098 180628 346108
rect 185612 220164 185668 514332
rect 203308 514108 203364 520940
rect 203308 514052 203700 514108
rect 190652 512820 190708 512830
rect 188972 502516 189028 502526
rect 188972 304164 189028 502460
rect 190652 431844 190708 512764
rect 192332 511140 192388 511150
rect 190652 431778 190708 431788
rect 191436 500724 191492 500734
rect 188972 304098 189028 304108
rect 185612 220098 185668 220108
rect 178892 176418 178948 176428
rect 179788 198324 179844 198334
rect 178780 480 178948 532
rect 178780 476 179144 480
rect 178780 420 178836 476
rect 178108 364 178836 420
rect 178892 392 179144 476
rect 178920 -960 179144 392
rect 179788 420 179844 198268
rect 182252 197876 182308 197886
rect 181468 21140 181524 21150
rect 180684 480 180852 532
rect 180684 476 181048 480
rect 180684 420 180740 476
rect 179788 364 180740 420
rect 180796 392 181048 476
rect 180824 -960 181048 392
rect 181468 420 181524 21084
rect 182252 9268 182308 197820
rect 182252 9202 182308 9212
rect 185612 175700 185668 175710
rect 184716 5012 184772 5022
rect 182588 480 182756 532
rect 184716 480 184772 4956
rect 185612 5012 185668 175644
rect 188972 172340 189028 172350
rect 185612 4946 185668 4956
rect 188412 16100 188468 16110
rect 186732 4116 186788 4126
rect 186732 480 186788 4060
rect 182588 476 182952 480
rect 182588 420 182644 476
rect 181468 364 182644 420
rect 182700 392 182952 476
rect 182728 -960 182952 392
rect 184632 -960 184856 480
rect 186536 392 186788 480
rect 188412 480 188468 16044
rect 188972 4116 189028 172284
rect 191436 58884 191492 500668
rect 192332 247044 192388 511084
rect 197372 509572 197428 509582
rect 194012 507892 194068 507902
rect 194012 332724 194068 507836
rect 195692 504532 195748 504542
rect 195692 374724 195748 504476
rect 195692 374658 195748 374668
rect 194012 332658 194068 332668
rect 197372 290724 197428 509516
rect 199836 502404 199892 502414
rect 199052 501060 199108 501070
rect 199052 416724 199108 501004
rect 199052 416658 199108 416668
rect 197372 290658 197428 290668
rect 192332 246978 192388 246988
rect 197372 197988 197428 197998
rect 191436 58818 191492 58828
rect 194012 192612 194068 192622
rect 191548 47908 191604 47918
rect 188972 4050 189028 4060
rect 190540 4116 190596 4126
rect 190540 480 190596 4060
rect 188412 392 188664 480
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 392 190596 480
rect 191548 420 191604 47852
rect 193228 37940 193284 37950
rect 192108 480 192276 532
rect 192108 476 192472 480
rect 192108 420 192164 476
rect 190344 -960 190568 392
rect 191548 364 192164 420
rect 192220 392 192472 476
rect 192248 -960 192472 392
rect 193228 420 193284 37884
rect 194012 4116 194068 192556
rect 194012 4050 194068 4060
rect 194908 179172 194964 179182
rect 194012 480 194180 532
rect 194012 476 194376 480
rect 194012 420 194068 476
rect 193228 364 194068 420
rect 194124 392 194376 476
rect 194152 -960 194376 392
rect 194908 420 194964 179116
rect 197372 44548 197428 197932
rect 197372 44482 197428 44492
rect 196588 36148 196644 36158
rect 195916 480 196084 532
rect 195916 476 196280 480
rect 195916 420 195972 476
rect 194908 364 195972 420
rect 196028 392 196280 476
rect 196056 -960 196280 392
rect 196588 420 196644 36092
rect 199836 34468 199892 502348
rect 203644 499940 203700 514052
rect 206668 499940 206724 529340
rect 208348 523348 208404 595644
rect 209468 595476 209524 595644
rect 209580 595560 209832 595672
rect 230188 595644 231588 595700
rect 231672 595672 231896 597000
rect 209580 595476 209636 595560
rect 209468 595420 209636 595476
rect 208348 523282 208404 523292
rect 213388 524244 213444 524254
rect 213388 514108 213444 524188
rect 223468 516068 223524 516078
rect 218428 514276 218484 514286
rect 218428 514108 218484 514220
rect 223468 514108 223524 516012
rect 213388 514052 214004 514108
rect 218428 514052 219156 514108
rect 223468 514052 224308 514108
rect 212156 504196 212212 504206
rect 209580 502404 209636 502414
rect 203644 499884 204456 499940
rect 206668 499884 207032 499940
rect 209580 499912 209636 502348
rect 212156 499912 212212 504140
rect 213948 499940 214004 514052
rect 217308 500724 217364 500734
rect 213948 499884 214760 499940
rect 217308 499912 217364 500668
rect 219100 499940 219156 514052
rect 221788 509236 221844 509246
rect 221788 499940 221844 509180
rect 224252 499940 224308 514052
rect 230188 503524 230244 595644
rect 231532 595476 231588 595644
rect 231644 595560 231896 595672
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 253736 595560 253988 595672
rect 275800 595560 276052 595672
rect 231644 595476 231700 595560
rect 231532 595420 231700 595476
rect 253932 591332 253988 595560
rect 253932 591266 253988 591276
rect 257852 591332 257908 591342
rect 257852 535220 257908 591276
rect 275996 591332 276052 595560
rect 297388 595644 297780 595700
rect 297864 595672 298088 597000
rect 275996 591266 276052 591276
rect 279692 591332 279748 591342
rect 279692 536788 279748 591276
rect 297388 543508 297444 595644
rect 297724 595476 297780 595644
rect 297836 595560 298088 595672
rect 319228 595644 319844 595700
rect 319928 595672 320152 597000
rect 297836 595476 297892 595560
rect 297724 595420 297892 595476
rect 319228 578788 319284 595644
rect 319788 595476 319844 595644
rect 319900 595560 320152 595672
rect 341068 595644 341908 595700
rect 341992 595672 342216 597000
rect 319900 595476 319956 595560
rect 319788 595420 319956 595476
rect 319228 578722 319284 578732
rect 297388 543442 297444 543452
rect 314972 561204 315028 561214
rect 279692 536722 279748 536732
rect 257852 535154 257908 535164
rect 311612 536004 311668 536014
rect 307468 531860 307524 531870
rect 235228 527716 235284 527726
rect 231868 519316 231924 519326
rect 231868 514108 231924 519260
rect 231868 514052 232036 514108
rect 230188 503458 230244 503468
rect 230300 512596 230356 512606
rect 227612 500724 227668 500734
rect 219100 499884 219912 499940
rect 221788 499884 222488 499940
rect 224252 499884 225064 499940
rect 227612 499912 227668 500668
rect 230300 499940 230356 512540
rect 230216 499884 230356 499940
rect 231980 499940 232036 514052
rect 235228 499940 235284 527660
rect 260428 526036 260484 526046
rect 241948 525924 242004 525934
rect 239372 515844 239428 515854
rect 237916 503972 237972 503982
rect 231980 499884 232792 499940
rect 235228 499884 235368 499940
rect 237916 499912 237972 503916
rect 239372 503972 239428 515788
rect 241948 514108 242004 525868
rect 250348 522788 250404 522798
rect 245308 521108 245364 521118
rect 241948 514052 242340 514108
rect 239372 503906 239428 503916
rect 240268 510916 240324 510926
rect 240268 499940 240324 510860
rect 242284 499940 242340 514052
rect 245308 499940 245364 521052
rect 246988 519428 247044 519438
rect 246988 514108 247044 519372
rect 246988 514052 247492 514108
rect 247436 499940 247492 514052
rect 250348 499940 250404 522732
rect 255388 517524 255444 517534
rect 252588 509348 252644 509358
rect 252588 499940 252644 509292
rect 255388 499940 255444 517468
rect 258524 504308 258580 504318
rect 240268 499884 240520 499940
rect 242284 499884 243096 499940
rect 245308 499884 245672 499940
rect 247436 499884 248248 499940
rect 250348 499884 250824 499940
rect 252588 499884 253400 499940
rect 255388 499884 255976 499940
rect 258524 499912 258580 504252
rect 260428 499940 260484 525980
rect 304108 522676 304164 522686
rect 278908 517860 278964 517870
rect 268828 514500 268884 514510
rect 263676 500836 263732 500846
rect 260428 499884 261128 499940
rect 263676 499912 263732 500780
rect 268828 499912 268884 514444
rect 273868 506212 273924 506222
rect 271404 502852 271460 502862
rect 271404 499912 271460 502796
rect 273868 499940 273924 506156
rect 275772 505876 275828 505886
rect 275772 499940 275828 505820
rect 278908 499940 278964 517804
rect 286076 512708 286132 512718
rect 280924 505764 280980 505774
rect 280924 499940 280980 505708
rect 286076 499940 286132 512652
rect 296380 511028 296436 511038
rect 288988 507668 289044 507678
rect 288988 499940 289044 507612
rect 294588 504420 294644 504430
rect 292012 500948 292068 500958
rect 273868 499884 274008 499940
rect 275772 499884 276584 499940
rect 278908 499884 279160 499940
rect 280924 499884 281736 499940
rect 286076 499884 286888 499940
rect 288988 499884 289464 499940
rect 292012 499912 292068 500892
rect 294588 499912 294644 504364
rect 296380 499940 296436 510972
rect 299068 509124 299124 509134
rect 299068 499940 299124 509068
rect 302316 501172 302372 501182
rect 296380 499884 297192 499940
rect 299068 499884 299768 499940
rect 302316 499912 302372 501116
rect 304108 499940 304164 522620
rect 304108 499884 304920 499940
rect 307468 499912 307524 531804
rect 310044 503972 310100 503982
rect 310044 499912 310100 503916
rect 311612 503972 311668 535948
rect 314188 535108 314244 535118
rect 314188 514108 314244 535052
rect 314188 514052 314468 514108
rect 311612 503906 311668 503916
rect 312620 504644 312676 504654
rect 312620 499912 312676 504588
rect 314412 499940 314468 514052
rect 314972 504644 315028 561148
rect 333452 547764 333508 547774
rect 324268 538468 324324 538478
rect 314972 504578 315028 504588
rect 317548 528388 317604 528398
rect 317548 499940 317604 528332
rect 319228 525028 319284 525038
rect 319228 514108 319284 524972
rect 322588 519988 322644 519998
rect 319228 514052 319620 514108
rect 319564 499940 319620 514052
rect 322588 499940 322644 519932
rect 324268 514108 324324 538412
rect 327628 533428 327684 533438
rect 324268 514052 324772 514108
rect 324716 499940 324772 514052
rect 327628 499940 327684 533372
rect 333452 531860 333508 547708
rect 339388 541828 339444 541838
rect 333452 531794 333508 531804
rect 334348 540148 334404 540158
rect 332668 531748 332724 531758
rect 330652 503412 330708 503422
rect 314412 499884 315224 499940
rect 317548 499884 317800 499940
rect 319564 499884 320376 499940
rect 322588 499884 322952 499940
rect 324716 499884 325528 499940
rect 327628 499884 328104 499940
rect 330652 499912 330708 503356
rect 332668 499940 332724 531692
rect 334348 514108 334404 540092
rect 339388 514108 339444 541772
rect 341068 521332 341124 595644
rect 341852 595476 341908 595644
rect 341964 595560 342216 595672
rect 362908 595644 363972 595700
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 341964 595476 342020 595560
rect 341852 595420 342020 595476
rect 362012 590548 362068 590558
rect 351148 578788 351204 578798
rect 343532 574644 343588 574654
rect 341068 521266 341124 521276
rect 342748 528500 342804 528510
rect 334348 514052 335076 514108
rect 339388 514052 340228 514108
rect 335020 499940 335076 514052
rect 338380 503636 338436 503646
rect 332668 499884 333256 499940
rect 335020 499884 335832 499940
rect 338380 499912 338436 503580
rect 340172 499940 340228 514052
rect 342748 499940 342804 528444
rect 343532 528388 343588 574588
rect 343532 528322 343588 528332
rect 346108 521332 346164 521342
rect 340172 499884 340984 499940
rect 342748 499884 343560 499940
rect 346108 499912 346164 521276
rect 348684 503748 348740 503758
rect 348684 499912 348740 503692
rect 351148 499940 351204 578732
rect 356188 543508 356244 543518
rect 352828 536788 352884 536798
rect 352828 514108 352884 536732
rect 352828 514052 353108 514108
rect 353052 499940 353108 514052
rect 356188 499940 356244 543452
rect 357868 535220 357924 535230
rect 357868 514108 357924 535164
rect 362012 528500 362068 590492
rect 362012 528434 362068 528444
rect 361228 523348 361284 523358
rect 357868 514052 358260 514108
rect 358204 499940 358260 514052
rect 361228 499940 361284 523292
rect 362908 503748 362964 595644
rect 363916 595476 363972 595644
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 473788 595644 474292 595700
rect 474376 595672 474600 597000
rect 364028 595476 364084 595560
rect 363916 595420 364084 595476
rect 365372 593236 365428 593246
rect 365372 503972 365428 593180
rect 380492 593124 380548 593134
rect 367948 585508 368004 585518
rect 367948 514108 368004 585452
rect 371308 551908 371364 551918
rect 367948 514052 368564 514108
rect 365372 503906 365428 503916
rect 366716 503972 366772 503982
rect 362908 503682 362964 503692
rect 364140 503524 364196 503534
rect 351148 499884 351288 499940
rect 353052 499884 353864 499940
rect 356188 499884 356440 499940
rect 358204 499884 359016 499940
rect 361228 499884 361592 499940
rect 364140 499912 364196 503468
rect 366716 499912 366772 503916
rect 368508 499940 368564 514052
rect 371308 499940 371364 551852
rect 378028 550228 378084 550238
rect 376348 526708 376404 526718
rect 372988 525140 373044 525150
rect 372988 514108 373044 525084
rect 372988 514052 373716 514108
rect 373660 499940 373716 514052
rect 376348 499940 376404 526652
rect 378028 514108 378084 550172
rect 378028 514052 378868 514108
rect 378812 499940 378868 514052
rect 380492 503972 380548 593068
rect 386092 590548 386148 595560
rect 386092 590482 386148 590492
rect 386428 583828 386484 583838
rect 386428 514108 386484 583772
rect 394828 572964 394884 572974
rect 389788 565348 389844 565358
rect 386428 514052 386596 514108
rect 380492 503906 380548 503916
rect 382172 503972 382228 503982
rect 368508 499884 369320 499940
rect 371308 499884 371896 499940
rect 373660 499884 374472 499940
rect 376348 499884 377048 499940
rect 378812 499884 379624 499940
rect 382172 499912 382228 503916
rect 384748 503300 384804 503310
rect 384748 499912 384804 503244
rect 386540 499940 386596 514052
rect 389788 499940 389844 565292
rect 391468 557844 391524 557854
rect 391468 514108 391524 557788
rect 393932 529284 393988 529294
rect 393932 514948 393988 529228
rect 393932 514882 393988 514892
rect 391468 514052 391748 514108
rect 391692 499940 391748 514052
rect 394828 499940 394884 572908
rect 396508 544404 396564 544414
rect 396508 514108 396564 544348
rect 401548 514948 401604 514958
rect 401548 514108 401604 514892
rect 396508 514052 396900 514108
rect 401548 514052 402052 514108
rect 396844 499940 396900 514052
rect 400204 503188 400260 503198
rect 386540 499884 387352 499940
rect 389788 499884 389928 499940
rect 391692 499884 392504 499940
rect 394828 499884 395080 499940
rect 396844 499884 397656 499940
rect 400204 499912 400260 503132
rect 401996 499940 402052 514052
rect 407932 504084 407988 504094
rect 405356 501508 405412 501518
rect 401996 499884 402808 499940
rect 405356 499912 405412 501452
rect 407932 499912 407988 504028
rect 408268 503636 408324 595560
rect 430220 572908 430276 595560
rect 430108 572852 430276 572908
rect 451052 590212 451108 590222
rect 430108 541828 430164 572852
rect 430108 541762 430164 541772
rect 451052 540148 451108 590156
rect 452284 590212 452340 595560
rect 452284 590146 452340 590156
rect 451052 540082 451108 540092
rect 463708 530964 463764 530974
rect 448588 527604 448644 527614
rect 433468 519204 433524 519214
rect 425068 516180 425124 516190
rect 425068 514108 425124 516124
rect 425068 514052 425236 514108
rect 414988 512820 415044 512830
rect 408268 503570 408324 503580
rect 409948 507556 410004 507566
rect 409948 499940 410004 507500
rect 414988 499940 415044 512764
rect 417452 509460 417508 509470
rect 417452 499940 417508 509404
rect 423388 506100 423444 506110
rect 420812 501060 420868 501070
rect 409948 499884 410536 499940
rect 414988 499884 415688 499940
rect 417452 499884 418264 499940
rect 420812 499912 420868 501004
rect 423388 499912 423444 506044
rect 425180 499940 425236 514052
rect 430332 505988 430388 505998
rect 428540 504532 428596 504542
rect 425180 499884 425992 499940
rect 428540 499912 428596 504476
rect 430332 499940 430388 505932
rect 433468 499940 433524 519148
rect 440188 514164 440244 514174
rect 440188 514052 440692 514108
rect 435484 507892 435540 507902
rect 435484 499940 435540 507836
rect 438844 502516 438900 502526
rect 430332 499884 431144 499940
rect 433468 499884 433720 499940
rect 435484 499884 436296 499940
rect 438844 499912 438900 502460
rect 440636 499940 440692 514052
rect 445788 510804 445844 510814
rect 443548 509572 443604 509582
rect 443548 499940 443604 509516
rect 445788 499940 445844 510748
rect 448588 499940 448644 527548
rect 455308 522564 455364 522574
rect 453628 514388 453684 514398
rect 450940 511140 450996 511150
rect 450940 499940 450996 511084
rect 453628 499940 453684 514332
rect 455308 514108 455364 522508
rect 458668 520884 458724 520894
rect 455308 514052 456148 514108
rect 456092 499940 456148 514052
rect 458668 499940 458724 520828
rect 463708 514108 463764 530908
rect 472108 517748 472164 517758
rect 463708 514052 463876 514108
rect 462028 507780 462084 507790
rect 440636 499884 441448 499940
rect 443548 499884 444024 499940
rect 445788 499884 446600 499940
rect 448588 499884 449176 499940
rect 450940 499884 451752 499940
rect 453628 499884 454328 499940
rect 456092 499884 456904 499940
rect 458668 499884 459480 499940
rect 462028 499912 462084 507724
rect 463820 499940 463876 514052
rect 468972 512484 469028 512494
rect 468972 499940 469028 512428
rect 472108 499940 472164 517692
rect 473788 503412 473844 595644
rect 474236 595476 474292 595644
rect 474348 595560 474600 595672
rect 495628 595644 496356 595700
rect 496440 595672 496664 597000
rect 474348 595476 474404 595560
rect 474236 595420 474404 595476
rect 495628 531748 495684 595644
rect 496300 595476 496356 595644
rect 496412 595560 496664 595672
rect 517468 595644 518420 595700
rect 518504 595672 518728 597000
rect 496412 595476 496468 595560
rect 496300 595420 496468 595476
rect 517468 533428 517524 595644
rect 518364 595476 518420 595644
rect 518476 595560 518728 595672
rect 539308 595644 540484 595700
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 518476 595476 518532 595560
rect 518364 595420 518532 595476
rect 517468 533362 517524 533372
rect 495628 531682 495684 531692
rect 523292 526036 523348 526046
rect 519932 521108 519988 521118
rect 487228 517636 487284 517646
rect 478828 515956 478884 515966
rect 478828 514108 478884 515900
rect 478828 514052 479332 514108
rect 473788 503346 473844 503356
rect 474908 502628 474964 502638
rect 463820 499884 464632 499940
rect 468972 499884 469784 499940
rect 472108 499884 472360 499940
rect 474908 499912 474964 502572
rect 477484 502516 477540 502526
rect 477484 499912 477540 502460
rect 479276 499940 479332 514052
rect 484428 507444 484484 507454
rect 482636 501060 482692 501070
rect 479276 499884 480088 499940
rect 482636 499912 482692 501004
rect 484428 499940 484484 507388
rect 487228 499940 487284 517580
rect 518252 512596 518308 512606
rect 516572 509236 516628 509246
rect 506492 506212 506548 506222
rect 495516 502964 495572 502974
rect 492940 502740 492996 502750
rect 490364 502404 490420 502414
rect 484428 499884 485240 499940
rect 487228 499884 487816 499940
rect 490364 499912 490420 502348
rect 492940 499912 492996 502684
rect 495516 499912 495572 502908
rect 500668 502628 500724 502638
rect 499100 501172 499156 501182
rect 467180 499380 467236 499390
rect 467180 499314 467236 499324
rect 266252 499268 266308 499278
rect 266252 499202 266308 499212
rect 284284 499268 284340 499278
rect 284284 499202 284340 499212
rect 413084 499268 413140 499278
rect 413084 499202 413140 499212
rect 498988 499044 499044 499054
rect 212828 198212 212884 198222
rect 209916 197652 209972 197662
rect 206668 190932 206724 190942
rect 199836 34402 199892 34412
rect 201628 187572 201684 187582
rect 199836 31220 199892 31230
rect 199836 4788 199892 31164
rect 201628 20188 201684 187516
rect 203308 185892 203364 185902
rect 201628 20132 201796 20188
rect 199836 4732 200004 4788
rect 197820 480 197988 532
rect 199948 480 200004 4732
rect 201740 480 201796 20132
rect 197820 476 198184 480
rect 197820 420 197876 476
rect 196588 364 197876 420
rect 197932 392 198184 476
rect 197960 -960 198184 392
rect 199864 -960 200088 480
rect 201740 392 201992 480
rect 201768 -960 201992 392
rect 203308 420 203364 185836
rect 205772 4116 205828 4126
rect 203532 480 203700 532
rect 205772 480 205828 4060
rect 203532 476 203896 480
rect 203532 420 203588 476
rect 203308 364 203588 420
rect 203644 392 203896 476
rect 203672 -960 203896 392
rect 205576 392 205828 480
rect 206668 420 206724 190876
rect 207452 51268 207508 51278
rect 207452 4116 207508 51212
rect 207452 4050 207508 4060
rect 208348 39508 208404 39518
rect 207340 480 207508 532
rect 207340 476 207704 480
rect 207340 420 207396 476
rect 205576 -960 205800 392
rect 206668 364 207396 420
rect 207452 392 207704 476
rect 207480 -960 207704 392
rect 208348 420 208404 39452
rect 209916 25172 209972 197596
rect 211708 196084 211764 196094
rect 209916 25106 209972 25116
rect 210028 194404 210084 194414
rect 209244 480 209412 532
rect 209244 476 209608 480
rect 209244 420 209300 476
rect 208348 364 209300 420
rect 209356 392 209608 476
rect 209384 -960 209608 392
rect 210028 420 210084 194348
rect 211148 480 211316 532
rect 211148 476 211512 480
rect 211148 420 211204 476
rect 210028 364 211204 420
rect 211260 392 211512 476
rect 211288 -960 211512 392
rect 211708 420 211764 196028
rect 212828 195748 212884 198156
rect 215516 198212 215572 200088
rect 215516 198146 215572 198156
rect 212828 195682 212884 195692
rect 214956 197316 215012 197326
rect 214956 5124 215012 197260
rect 216412 31108 216468 200088
rect 217308 192388 217364 200088
rect 217308 192322 217364 192332
rect 216412 31042 216468 31052
rect 214956 5058 215012 5068
rect 215068 25172 215124 25182
rect 213052 480 213220 532
rect 215068 480 215124 25116
rect 218204 6244 218260 200088
rect 219100 197540 219156 200088
rect 219100 197474 219156 197484
rect 218204 6178 218260 6188
rect 217196 5796 217252 5806
rect 217196 480 217252 5740
rect 213052 476 213416 480
rect 213052 420 213108 476
rect 211708 364 213108 420
rect 213164 392 213416 476
rect 215068 392 215320 480
rect 213192 -960 213416 392
rect 215096 -960 215320 392
rect 217000 392 217252 480
rect 218876 5124 218932 5134
rect 218876 480 218932 5068
rect 219996 4228 220052 200088
rect 219996 4162 220052 4172
rect 220108 195748 220164 195758
rect 218876 392 219128 480
rect 217000 -960 217224 392
rect 218904 -960 219128 392
rect 220108 420 220164 195692
rect 220892 190708 220948 200088
rect 221788 197764 221844 200088
rect 221788 197698 221844 197708
rect 222684 194068 222740 200088
rect 222684 194002 222740 194012
rect 220892 190642 220948 190652
rect 223580 4340 223636 200088
rect 224476 197988 224532 200088
rect 224476 197922 224532 197932
rect 223692 197764 223748 197774
rect 223692 197316 223748 197708
rect 223692 197250 223748 197260
rect 224252 197540 224308 197550
rect 224252 157108 224308 197484
rect 225372 189028 225428 200088
rect 225372 188962 225428 188972
rect 224252 157042 224308 157052
rect 223580 4274 223636 4284
rect 225932 29540 225988 29550
rect 224812 4228 224868 4238
rect 222908 2660 222964 2670
rect 220668 480 220836 532
rect 222908 480 222964 2604
rect 224812 480 224868 4172
rect 225932 4228 225988 29484
rect 226268 14308 226324 200088
rect 226268 14242 226324 14252
rect 225932 4162 225988 4172
rect 226716 11060 226772 11070
rect 226716 480 226772 11004
rect 227164 4452 227220 200088
rect 228060 189140 228116 200088
rect 228060 189074 228116 189084
rect 228956 178948 229012 200088
rect 228956 178882 229012 178892
rect 229852 56308 229908 200088
rect 229852 56242 229908 56252
rect 230300 44548 230356 44558
rect 227164 4386 227220 4396
rect 228508 19460 228564 19470
rect 228508 480 228564 19404
rect 230300 480 230356 44492
rect 230748 4564 230804 200088
rect 231644 187348 231700 200088
rect 231644 187282 231700 187292
rect 232540 180628 232596 200088
rect 232540 180562 232596 180572
rect 233436 52948 233492 200088
rect 233436 52882 233492 52892
rect 233548 200060 234360 200116
rect 230748 4498 230804 4508
rect 231868 46228 231924 46238
rect 220668 476 221032 480
rect 220668 420 220724 476
rect 220108 364 220724 420
rect 220780 392 221032 476
rect 220808 -960 221032 392
rect 222712 392 222964 480
rect 224616 392 224868 480
rect 226520 392 226772 480
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 480
rect 230300 392 230552 480
rect 230328 -960 230552 392
rect 231868 420 231924 46172
rect 233548 4676 233604 200060
rect 234332 198212 234388 198222
rect 234332 158788 234388 198156
rect 235228 160468 235284 200088
rect 235228 160402 235284 160412
rect 234332 158722 234388 158732
rect 236124 54628 236180 200088
rect 237020 195860 237076 200088
rect 237916 198212 237972 200088
rect 237916 198146 237972 198156
rect 237020 195794 237076 195804
rect 238812 165508 238868 200088
rect 238812 165442 238868 165452
rect 239708 61348 239764 200088
rect 240604 197540 240660 200088
rect 241500 199108 241556 200088
rect 241500 199042 241556 199052
rect 240604 197474 240660 197484
rect 241948 197540 242004 197550
rect 241948 194404 242004 197484
rect 241948 194338 242004 194348
rect 242396 167188 242452 200088
rect 242396 167122 242452 167132
rect 239708 61282 239764 61292
rect 236124 54562 236180 54572
rect 243292 37828 243348 200088
rect 244188 182308 244244 200088
rect 244188 182242 244244 182252
rect 245084 66388 245140 200088
rect 245980 155428 246036 200088
rect 245980 155362 246036 155372
rect 245084 66322 245140 66332
rect 243292 37762 243348 37772
rect 243628 31108 243684 31118
rect 233548 4610 233604 4620
rect 233660 24500 233716 24510
rect 232092 480 232260 532
rect 232092 476 232456 480
rect 232092 420 232148 476
rect 231868 364 232148 420
rect 232204 392 232456 476
rect 232232 -960 232456 392
rect 233660 420 233716 24444
rect 238588 12740 238644 12750
rect 236236 7812 236292 7822
rect 233996 480 234164 532
rect 236236 480 236292 7756
rect 238140 6132 238196 6142
rect 238140 480 238196 6076
rect 233996 476 234360 480
rect 233996 420 234052 476
rect 233660 364 234052 420
rect 234108 392 234360 476
rect 234136 -960 234360 392
rect 236040 392 236292 480
rect 237944 392 238196 480
rect 238588 420 238644 12684
rect 241836 2772 241892 2782
rect 239708 480 239876 532
rect 241836 480 241892 2716
rect 243628 480 243684 31052
rect 246876 7588 246932 200088
rect 246876 7522 246932 7532
rect 246988 192388 247044 192398
rect 245756 480 245924 532
rect 239708 476 240072 480
rect 239708 420 239764 476
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 238588 364 239764 420
rect 239820 392 240072 476
rect 239848 -960 240072 392
rect 241752 -960 241976 480
rect 243628 392 243880 480
rect 243656 -960 243880 392
rect 245560 476 245924 480
rect 245560 392 245812 476
rect 245560 -960 245784 392
rect 245868 84 245924 476
rect 246988 420 247044 192332
rect 247772 147028 247828 200088
rect 248668 185668 248724 200088
rect 248668 185602 248724 185612
rect 247772 146962 247828 146972
rect 248668 184212 248724 184222
rect 247324 480 247492 532
rect 247324 476 247688 480
rect 247324 420 247380 476
rect 246988 364 247380 420
rect 247436 392 247688 476
rect 245868 18 245924 28
rect 247464 -960 247688 392
rect 248668 420 248724 184156
rect 249564 17668 249620 200088
rect 249564 17602 249620 17612
rect 250460 4788 250516 200088
rect 251356 175588 251412 200088
rect 251356 175522 251412 175532
rect 252028 189028 252084 189038
rect 250460 4722 250516 4732
rect 251468 4228 251524 4238
rect 249228 480 249396 532
rect 251468 480 251524 4172
rect 249228 476 249592 480
rect 249228 420 249284 476
rect 248668 364 249284 420
rect 249340 392 249592 476
rect 249368 -960 249592 392
rect 251272 392 251524 480
rect 252028 420 252084 188972
rect 252252 183988 252308 200088
rect 252252 183922 252308 183932
rect 253148 32900 253204 200088
rect 254044 197428 254100 200088
rect 254044 197362 254100 197372
rect 254492 197428 254548 197438
rect 253708 196644 253764 196654
rect 253708 192500 253764 196588
rect 253708 192434 253764 192444
rect 254492 184100 254548 197372
rect 254492 184034 254548 184044
rect 253148 32834 253204 32844
rect 252812 32788 252868 32798
rect 252812 4228 252868 32732
rect 252812 4162 252868 4172
rect 253820 17668 253876 17678
rect 253036 480 253204 532
rect 253036 476 253400 480
rect 253036 420 253092 476
rect 251272 -960 251496 392
rect 252028 364 253092 420
rect 253148 392 253400 476
rect 253176 -960 253400 392
rect 253820 420 253876 17612
rect 254940 6020 254996 200088
rect 255836 185780 255892 200088
rect 256732 196644 256788 200088
rect 256732 196578 256788 196588
rect 257068 197204 257124 197214
rect 257068 194180 257124 197148
rect 257068 194114 257124 194124
rect 255836 185714 255892 185724
rect 257628 153748 257684 200088
rect 257628 153682 257684 153692
rect 254940 5954 254996 5964
rect 257180 14532 257236 14542
rect 254940 480 255108 532
rect 257180 480 257236 14476
rect 258524 10948 258580 200088
rect 259420 197204 259476 200088
rect 260316 197428 260372 200088
rect 260316 197362 260372 197372
rect 260428 200060 261240 200116
rect 259420 197138 259476 197148
rect 260428 148708 260484 200060
rect 260428 148642 260484 148652
rect 261212 194068 261268 194078
rect 258524 10882 258580 10892
rect 260988 9268 261044 9278
rect 259084 4228 259140 4238
rect 259084 480 259140 4172
rect 260988 480 261044 9212
rect 261212 4228 261268 194012
rect 262108 173908 262164 200088
rect 262108 173842 262164 173852
rect 263004 24388 263060 200088
rect 263004 24322 263060 24332
rect 263788 200060 263928 200116
rect 261212 4162 261268 4172
rect 262108 14644 262164 14654
rect 254940 476 255304 480
rect 254940 420 254996 476
rect 253820 364 254996 420
rect 255052 392 255304 476
rect 255080 -960 255304 392
rect 256984 392 257236 480
rect 258888 392 259140 480
rect 260792 392 261044 480
rect 262108 420 262164 14588
rect 263788 2548 263844 200060
rect 264572 197428 264628 197438
rect 264572 187460 264628 197372
rect 264572 187394 264628 187404
rect 264796 172228 264852 200088
rect 265692 182420 265748 200088
rect 265692 182354 265748 182364
rect 264796 172162 264852 172172
rect 266588 42980 266644 200088
rect 267484 170548 267540 200088
rect 267484 170482 267540 170492
rect 266588 42914 266644 42924
rect 266252 42868 266308 42878
rect 265468 21252 265524 21262
rect 263788 2482 263844 2492
rect 264796 4228 264852 4238
rect 262556 480 262724 532
rect 264796 480 264852 4172
rect 262556 476 262920 480
rect 262556 420 262612 476
rect 256984 -960 257208 392
rect 258888 -960 259112 392
rect 260792 -960 261016 392
rect 262108 364 262612 420
rect 262668 392 262920 476
rect 262696 -960 262920 392
rect 264600 392 264852 480
rect 265468 420 265524 21196
rect 266252 4228 266308 42812
rect 268380 15988 268436 200088
rect 269276 19348 269332 200088
rect 270172 168868 270228 200088
rect 270172 168802 270228 168812
rect 271068 152068 271124 200088
rect 271068 152002 271124 152012
rect 271964 21028 272020 200088
rect 272860 195972 272916 200088
rect 273756 197428 273812 200088
rect 273756 197362 273812 197372
rect 273868 200060 274680 200116
rect 272860 195906 272916 195916
rect 273868 177268 273924 200060
rect 273868 177202 273924 177212
rect 274652 197428 274708 197438
rect 271964 20962 272020 20972
rect 269276 19282 269332 19292
rect 268380 15922 268436 15932
rect 266252 4162 266308 4172
rect 267148 14420 267204 14430
rect 266364 480 266532 532
rect 266364 476 266728 480
rect 266364 420 266420 476
rect 264600 -960 264824 392
rect 265468 364 266420 420
rect 266476 392 266728 476
rect 266504 -960 266728 392
rect 267148 420 267204 14364
rect 274316 9492 274372 9502
rect 270396 6804 270452 6814
rect 268268 480 268436 532
rect 270396 480 270452 6748
rect 272412 4228 272468 4238
rect 272412 480 272468 4172
rect 274316 480 274372 9436
rect 274652 6804 274708 197372
rect 275548 196588 275604 200088
rect 275436 196532 275604 196588
rect 275436 194292 275492 196532
rect 275436 194226 275492 194236
rect 276444 182532 276500 200088
rect 276444 182466 276500 182476
rect 277340 179060 277396 200088
rect 278236 199220 278292 200088
rect 278236 199154 278292 199164
rect 277340 178994 277396 179004
rect 279132 174020 279188 200088
rect 279132 173954 279188 173964
rect 274652 6738 274708 6748
rect 274764 32900 274820 32910
rect 274764 4228 274820 32844
rect 279020 22820 279076 22830
rect 277228 12852 277284 12862
rect 274764 4162 274820 4172
rect 276220 7588 276276 7598
rect 276220 480 276276 7532
rect 268268 476 268632 480
rect 268268 420 268324 476
rect 267148 364 268324 420
rect 268380 392 268632 476
rect 268408 -960 268632 392
rect 270312 -960 270536 480
rect 272216 392 272468 480
rect 274120 392 274372 480
rect 276024 392 276276 480
rect 277228 420 277284 12796
rect 277788 480 277956 532
rect 277788 476 278152 480
rect 277788 420 277844 476
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277228 364 277844 420
rect 277900 392 278152 476
rect 277928 -960 278152 392
rect 279020 420 279076 22764
rect 280028 17780 280084 200088
rect 280924 167300 280980 200088
rect 280924 167234 280980 167244
rect 281820 29428 281876 200088
rect 281820 29362 281876 29372
rect 280028 17714 280084 17724
rect 281932 10948 281988 10958
rect 279692 480 279860 532
rect 281932 480 281988 10892
rect 282716 9380 282772 200088
rect 283052 196756 283108 196766
rect 283052 93268 283108 196700
rect 283612 190820 283668 200088
rect 283612 190754 283668 190764
rect 284508 150388 284564 200088
rect 284508 150322 284564 150332
rect 283052 93202 283108 93212
rect 285404 12628 285460 200088
rect 285404 12562 285460 12572
rect 285628 180964 285684 180974
rect 282716 9314 282772 9324
rect 283836 6020 283892 6030
rect 283836 480 283892 5964
rect 285628 480 285684 180908
rect 286300 165620 286356 200088
rect 287196 180740 287252 200088
rect 287196 180674 287252 180684
rect 287308 200060 288120 200116
rect 286300 165554 286356 165564
rect 287308 7700 287364 200060
rect 288092 196644 288148 196654
rect 288092 135268 288148 196588
rect 288988 162148 289044 200088
rect 288988 162082 289044 162092
rect 288092 135202 288148 135212
rect 289884 49588 289940 200088
rect 290780 196756 290836 200088
rect 290780 196690 290836 196700
rect 291676 196644 291732 200088
rect 291676 196578 291732 196588
rect 292348 198212 292404 198222
rect 292348 189252 292404 198156
rect 292348 189186 292404 189196
rect 292572 177380 292628 200088
rect 292572 177314 292628 177324
rect 289884 49522 289940 49532
rect 293468 22708 293524 200088
rect 294364 198212 294420 200088
rect 294588 200060 295288 200116
rect 294588 198324 294644 200060
rect 294588 198258 294644 198268
rect 294364 198146 294420 198156
rect 293468 22642 293524 22652
rect 296156 21140 296212 200088
rect 297052 175700 297108 200088
rect 297052 175634 297108 175644
rect 297948 172340 298004 200088
rect 297948 172274 298004 172284
rect 296156 21074 296212 21084
rect 297500 24388 297556 24398
rect 292348 19348 292404 19358
rect 287308 7634 287364 7644
rect 287420 16212 287476 16222
rect 287420 480 287476 16156
rect 289548 11284 289604 11294
rect 289548 480 289604 11228
rect 291452 7700 291508 7710
rect 291452 480 291508 7644
rect 279692 476 280056 480
rect 279692 420 279748 476
rect 279020 364 279748 420
rect 279804 392 280056 476
rect 279832 -960 280056 392
rect 281736 392 281988 480
rect 283640 392 283892 480
rect 281736 -960 281960 392
rect 283640 -960 283864 392
rect 285544 -960 285768 480
rect 287420 392 287672 480
rect 287448 -960 287672 392
rect 289352 392 289604 480
rect 291256 392 291508 480
rect 292348 420 292404 19292
rect 295708 12628 295764 12638
rect 295260 2548 295316 2558
rect 293020 480 293188 532
rect 295260 480 295316 2492
rect 293020 476 293384 480
rect 293020 420 293076 476
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 292348 364 293076 420
rect 293132 392 293384 476
rect 293160 -960 293384 392
rect 295064 392 295316 480
rect 295708 420 295764 12572
rect 296828 480 296996 532
rect 296828 476 297192 480
rect 296828 420 296884 476
rect 295064 -960 295288 392
rect 295708 364 296884 420
rect 296940 392 297192 476
rect 296968 -960 297192 392
rect 297500 420 297556 24332
rect 298844 16100 298900 200088
rect 299740 192612 299796 200088
rect 299740 192546 299796 192556
rect 300636 47908 300692 200088
rect 300636 47842 300692 47852
rect 300748 200060 301560 200116
rect 300748 37940 300804 200060
rect 300860 197988 300916 197998
rect 300860 196084 300916 197932
rect 300860 196018 300916 196028
rect 302428 179172 302484 200088
rect 302428 179106 302484 179116
rect 300748 37874 300804 37884
rect 298844 16034 298900 16044
rect 300972 37828 301028 37838
rect 298732 480 298900 532
rect 300972 480 301028 37772
rect 303324 36148 303380 200088
rect 303324 36082 303380 36092
rect 304220 31220 304276 200088
rect 305116 187572 305172 200088
rect 305116 187506 305172 187516
rect 306012 185892 306068 200088
rect 306012 185826 306068 185836
rect 306908 51268 306964 200088
rect 307804 190932 307860 200088
rect 307804 190866 307860 190876
rect 308252 197876 308308 197886
rect 306908 51202 306964 51212
rect 304220 31154 304276 31164
rect 305788 36148 305844 36158
rect 302428 29652 302484 29662
rect 302428 20188 302484 29596
rect 302428 20132 302708 20188
rect 298732 476 299096 480
rect 298732 420 298788 476
rect 297500 364 298788 420
rect 298844 392 299096 476
rect 298872 -960 299096 392
rect 300776 392 301028 480
rect 302652 480 302708 20132
rect 304108 17780 304164 17790
rect 302652 392 302904 480
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304108 420 304164 17724
rect 304444 480 304612 532
rect 304444 476 304808 480
rect 304444 420 304500 476
rect 304108 364 304500 420
rect 304556 392 304808 476
rect 304584 -960 304808 392
rect 305788 420 305844 36092
rect 308252 16212 308308 197820
rect 308700 39508 308756 200088
rect 309596 197540 309652 200088
rect 310492 197988 310548 200088
rect 310492 197922 310548 197932
rect 311388 197652 311444 200088
rect 311388 197586 311444 197596
rect 309596 197474 309652 197484
rect 311612 197540 311668 197550
rect 308700 39442 308756 39452
rect 308252 16146 308308 16156
rect 307468 15988 307524 15998
rect 306348 480 306516 532
rect 306348 476 306712 480
rect 306348 420 306404 476
rect 305788 364 306404 420
rect 306460 392 306712 476
rect 306488 -960 306712 392
rect 307468 420 307524 15932
rect 311612 11284 311668 197484
rect 311612 11218 311668 11228
rect 310492 6244 310548 6254
rect 308252 480 308420 532
rect 310492 480 310548 6188
rect 312284 5908 312340 200088
rect 313180 197764 313236 200088
rect 313180 197698 313236 197708
rect 314076 195748 314132 200088
rect 314076 195682 314132 195692
rect 314188 200060 315000 200116
rect 312284 5842 312340 5852
rect 312396 11172 312452 11182
rect 312396 480 312452 11116
rect 314188 2660 314244 200060
rect 314972 198212 315028 198222
rect 314188 2594 314244 2604
rect 314300 3556 314356 3566
rect 314300 480 314356 3500
rect 314972 2772 315028 198156
rect 315868 29540 315924 200088
rect 315868 29474 315924 29484
rect 316652 21028 316708 21038
rect 314972 2706 315028 2716
rect 316204 7924 316260 7934
rect 316204 480 316260 7868
rect 316652 3556 316708 20972
rect 316764 11060 316820 200088
rect 317548 200060 317688 200116
rect 317548 19460 317604 200060
rect 318556 44548 318612 200088
rect 319452 46228 319508 200088
rect 319452 46162 319508 46172
rect 318556 44482 318612 44492
rect 320348 24500 320404 200088
rect 320348 24434 320404 24444
rect 317548 19394 317604 19404
rect 317884 19460 317940 19470
rect 316764 10994 316820 11004
rect 316652 3490 316708 3500
rect 308252 476 308616 480
rect 308252 420 308308 476
rect 307468 364 308308 420
rect 308364 392 308616 476
rect 308392 -960 308616 392
rect 310296 392 310548 480
rect 312200 392 312452 480
rect 314104 392 314356 480
rect 316008 392 316260 480
rect 317884 480 317940 19404
rect 321244 7812 321300 200088
rect 321244 7746 321300 7756
rect 322140 6132 322196 200088
rect 322140 6066 322196 6076
rect 322700 16100 322756 16110
rect 321916 5908 321972 5918
rect 320012 4228 320068 4238
rect 320012 480 320068 4172
rect 321916 480 321972 5852
rect 317884 392 318136 480
rect 310296 -960 310520 392
rect 312200 -960 312424 392
rect 314104 -960 314328 392
rect 316008 -960 316232 392
rect 317912 -960 318136 392
rect 319816 392 320068 480
rect 321720 392 321972 480
rect 322700 420 322756 16044
rect 323036 12740 323092 200088
rect 323932 198212 323988 200088
rect 323932 198146 323988 198156
rect 324268 198322 324324 198334
rect 324268 198270 324270 198322
rect 324322 198270 324324 198322
rect 323372 197764 323428 197774
rect 323372 14532 323428 197708
rect 323372 14466 323428 14476
rect 323036 12674 323092 12684
rect 323484 480 323652 532
rect 323484 476 323848 480
rect 323484 420 323540 476
rect 319816 -960 320040 392
rect 321720 -960 321944 392
rect 322700 364 323540 420
rect 323596 392 323848 476
rect 323624 -960 323848 392
rect 324268 84 324324 198270
rect 324380 196644 324436 196654
rect 324380 192388 324436 196588
rect 324380 192322 324436 192332
rect 324828 31108 324884 200088
rect 325052 200060 325752 200116
rect 325052 198322 325108 200060
rect 325052 198270 325054 198322
rect 325106 198270 325108 198322
rect 325052 198258 325108 198270
rect 326620 196644 326676 200088
rect 326620 196578 326676 196588
rect 327516 184212 327572 200088
rect 327516 184146 327572 184156
rect 327628 200060 328440 200116
rect 327628 32788 327684 200060
rect 327628 32722 327684 32732
rect 328412 197652 328468 197662
rect 324828 31042 324884 31052
rect 327516 5124 327572 5134
rect 325724 5012 325780 5022
rect 325724 480 325780 4956
rect 327516 480 327572 5068
rect 328412 5124 328468 197596
rect 329308 189028 329364 200088
rect 329308 188962 329364 188972
rect 329532 195748 329588 195758
rect 328412 5058 328468 5068
rect 329532 480 329588 195692
rect 330204 17668 330260 200088
rect 331100 197764 331156 200088
rect 331100 197698 331156 197708
rect 331996 194068 332052 200088
rect 331996 194002 332052 194012
rect 330204 17602 330260 17612
rect 332892 9268 332948 200088
rect 333788 14644 333844 200088
rect 334684 42868 334740 200088
rect 334684 42802 334740 42812
rect 333788 14578 333844 14588
rect 334460 29428 334516 29438
rect 332892 9202 332948 9212
rect 333116 14308 333172 14318
rect 331436 4452 331492 4462
rect 331436 480 331492 4396
rect 324268 18 324324 28
rect 325528 392 325780 480
rect 325528 -960 325752 392
rect 327432 -960 327656 480
rect 329336 392 329588 480
rect 331240 392 331492 480
rect 333116 480 333172 14252
rect 333116 392 333368 480
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 334460 420 334516 29372
rect 335580 21252 335636 200088
rect 335580 21186 335636 21196
rect 336476 14420 336532 200088
rect 336812 197764 336868 197774
rect 336812 29652 336868 197708
rect 337372 197428 337428 200088
rect 337372 197362 337428 197372
rect 338268 32900 338324 200088
rect 338268 32834 338324 32844
rect 336812 29586 336868 29596
rect 336476 14354 336532 14364
rect 339052 11060 339108 11070
rect 337148 4564 337204 4574
rect 334908 480 335076 532
rect 337148 480 337204 4508
rect 339052 480 339108 11004
rect 339164 9492 339220 200088
rect 340060 197428 340116 200088
rect 340060 197362 340116 197372
rect 340172 198100 340228 198110
rect 339164 9426 339220 9436
rect 339500 32788 339556 32798
rect 334908 476 335272 480
rect 334908 420 334964 476
rect 334460 364 334964 420
rect 335020 392 335272 476
rect 335048 -960 335272 392
rect 336952 392 337204 480
rect 338856 392 339108 480
rect 339500 420 339556 32732
rect 340172 2548 340228 198044
rect 340956 12852 341012 200088
rect 341068 200060 341880 200116
rect 341068 22820 341124 200060
rect 341068 22754 341124 22764
rect 341852 198212 341908 198222
rect 340956 12786 341012 12796
rect 341852 10948 341908 198156
rect 342748 198212 342804 200088
rect 342748 198146 342804 198156
rect 343532 197092 343588 197102
rect 343532 19348 343588 197036
rect 343532 19282 343588 19292
rect 341852 10882 341908 10892
rect 343644 6020 343700 200088
rect 343756 198212 343812 198222
rect 343756 180964 343812 198156
rect 344540 198212 344596 200088
rect 344540 198146 344596 198156
rect 345436 197876 345492 200088
rect 345436 197810 345492 197820
rect 346332 197540 346388 200088
rect 346332 197474 346388 197484
rect 343756 180898 343812 180908
rect 346108 195860 346164 195870
rect 343644 5954 343700 5964
rect 344764 6020 344820 6030
rect 340172 2482 340228 2492
rect 342860 4676 342916 4686
rect 340620 480 340788 532
rect 342860 480 342916 4620
rect 344764 480 344820 5964
rect 340620 476 340984 480
rect 340620 420 340676 476
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 339500 364 340676 420
rect 340732 392 340984 476
rect 340760 -960 340984 392
rect 342664 392 342916 480
rect 344568 392 344820 480
rect 346108 420 346164 195804
rect 347228 7700 347284 200088
rect 348124 197092 348180 200088
rect 349020 198100 349076 200088
rect 349020 198034 349076 198044
rect 348124 197026 348180 197036
rect 347228 7634 347284 7644
rect 349580 19348 349636 19358
rect 348572 4788 348628 4798
rect 346332 480 346500 532
rect 348572 480 348628 4732
rect 346332 476 346696 480
rect 346332 420 346388 476
rect 342664 -960 342888 392
rect 344568 -960 344792 392
rect 346108 364 346388 420
rect 346444 392 346696 476
rect 346472 -960 346696 392
rect 348376 392 348628 480
rect 349580 420 349636 19292
rect 349916 12628 349972 200088
rect 350812 24388 350868 200088
rect 351708 37828 351764 200088
rect 351708 37762 351764 37772
rect 351932 197988 351988 197998
rect 350812 24322 350868 24332
rect 351148 31108 351204 31118
rect 349916 12562 349972 12572
rect 350140 480 350308 532
rect 350140 476 350504 480
rect 350140 420 350196 476
rect 348376 -960 348600 392
rect 349580 364 350196 420
rect 350252 392 350504 476
rect 350280 -960 350504 392
rect 351148 420 351204 31052
rect 351932 15988 351988 197932
rect 352604 197764 352660 200088
rect 352604 197698 352660 197708
rect 353500 17780 353556 200088
rect 354396 36148 354452 200088
rect 354620 200060 355320 200116
rect 354620 197988 354676 200060
rect 354620 197922 354676 197932
rect 355292 198212 355348 198222
rect 354396 36082 354452 36092
rect 354508 197428 354564 197438
rect 353500 17714 353556 17724
rect 351932 15922 351988 15932
rect 354508 7588 354564 197372
rect 354508 7522 354564 7532
rect 355292 6244 355348 198156
rect 356188 198212 356244 200088
rect 356188 198146 356244 198156
rect 356972 197092 357028 197102
rect 356972 7924 357028 197036
rect 357084 11172 357140 200088
rect 357084 11106 357140 11116
rect 357868 195972 357924 195982
rect 356972 7858 357028 7868
rect 355292 6178 355348 6188
rect 356076 7588 356132 7598
rect 354284 4900 354340 4910
rect 352044 480 352212 532
rect 354284 480 354340 4844
rect 356076 480 356132 7532
rect 357868 480 357924 195916
rect 357980 21028 358036 200088
rect 358876 197092 358932 200088
rect 358876 197026 358932 197036
rect 359548 197428 359604 197438
rect 357980 20962 358036 20972
rect 359548 8428 359604 197372
rect 359772 19460 359828 200088
rect 359772 19394 359828 19404
rect 359548 8372 359828 8428
rect 359772 480 359828 8372
rect 360668 4228 360724 200088
rect 361228 200060 361592 200116
rect 361228 5908 361284 200060
rect 362460 16100 362516 200088
rect 362460 16034 362516 16044
rect 361228 5842 361284 5852
rect 361676 15988 361732 15998
rect 360668 4162 360724 4172
rect 361676 480 361732 15932
rect 363356 5012 363412 200088
rect 364252 197652 364308 200088
rect 364252 197586 364308 197596
rect 365148 195748 365204 200088
rect 365148 195682 365204 195692
rect 365372 197764 365428 197774
rect 365372 32788 365428 197708
rect 365372 32722 365428 32732
rect 363356 4946 363412 4956
rect 365708 8484 365764 8494
rect 363804 4340 363860 4350
rect 363804 480 363860 4284
rect 365708 480 365764 8428
rect 366044 4452 366100 200088
rect 366968 200060 367668 200116
rect 367612 196588 367668 200060
rect 367836 198212 367892 200088
rect 367836 198146 367892 198156
rect 367612 196532 368116 196588
rect 368060 14308 368116 196532
rect 368060 14242 368116 14252
rect 368732 4564 368788 200088
rect 369628 11060 369684 200088
rect 370524 197764 370580 200088
rect 370524 197698 370580 197708
rect 371308 200060 371448 200116
rect 369628 10994 369684 11004
rect 370412 197316 370468 197326
rect 370412 6020 370468 197260
rect 370412 5954 370468 5964
rect 371308 4676 371364 200060
rect 371420 198212 371476 198222
rect 371420 29428 371476 198156
rect 372316 197316 372372 200088
rect 372316 197250 372372 197260
rect 373212 195860 373268 200088
rect 373212 195794 373268 195804
rect 373772 198212 373828 198222
rect 373772 31108 373828 198156
rect 373772 31042 373828 31052
rect 371420 29362 371476 29372
rect 371308 4610 371364 4620
rect 373324 6804 373380 6814
rect 368732 4498 368788 4508
rect 371420 4564 371476 4574
rect 366044 4386 366100 4396
rect 369516 4452 369572 4462
rect 367612 4228 367668 4238
rect 367612 480 367668 4172
rect 369516 480 369572 4396
rect 371420 480 371476 4508
rect 373324 480 373380 6748
rect 374108 4788 374164 200088
rect 375004 19348 375060 200088
rect 375900 198212 375956 200088
rect 375900 198146 375956 198156
rect 375004 19282 375060 19292
rect 375452 198100 375508 198110
rect 374108 4722 374164 4732
rect 375228 8820 375284 8830
rect 375228 480 375284 8764
rect 375452 8484 375508 198044
rect 375452 8418 375508 8428
rect 376796 4900 376852 200088
rect 377692 7588 377748 200088
rect 378588 195972 378644 200088
rect 378588 195906 378644 195916
rect 378812 198212 378868 198222
rect 377692 7522 377748 7532
rect 378028 195748 378084 195758
rect 376796 4834 376852 4844
rect 377132 5012 377188 5022
rect 377132 480 377188 4956
rect 352044 476 352408 480
rect 352044 420 352100 476
rect 351148 364 352100 420
rect 352156 392 352408 476
rect 352184 -960 352408 392
rect 354088 392 354340 480
rect 354088 -960 354312 392
rect 355992 -960 356216 480
rect 357868 392 358120 480
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 392 363860 480
rect 365512 392 365764 480
rect 367416 392 367668 480
rect 369320 392 369572 480
rect 371224 392 371476 480
rect 373128 392 373380 480
rect 375032 392 375284 480
rect 376936 392 377188 480
rect 378028 420 378084 195692
rect 378812 15988 378868 198156
rect 379484 197428 379540 200088
rect 379708 200060 380408 200116
rect 380492 200060 381304 200116
rect 379708 198212 379764 200060
rect 380492 198324 380548 200060
rect 379708 198146 379764 198156
rect 379820 198268 380548 198324
rect 379484 197362 379540 197372
rect 378812 15922 378868 15932
rect 379820 4340 379876 198268
rect 382172 198100 382228 200088
rect 382172 198034 382228 198044
rect 380492 196756 380548 196766
rect 380492 8820 380548 196700
rect 380492 8754 380548 8764
rect 379820 4274 379876 4284
rect 380940 4788 380996 4798
rect 378700 480 378868 532
rect 380940 480 380996 4732
rect 382844 4340 382900 4350
rect 382844 480 382900 4284
rect 383068 4228 383124 200088
rect 383852 196644 383908 196654
rect 383068 4162 383124 4172
rect 383292 12628 383348 12638
rect 378700 476 379064 480
rect 378700 420 378756 476
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 369320 -960 369544 392
rect 371224 -960 371448 392
rect 373128 -960 373352 392
rect 375032 -960 375256 392
rect 376936 -960 377160 392
rect 378028 364 378756 420
rect 378812 392 379064 476
rect 378840 -960 379064 392
rect 380744 392 380996 480
rect 382648 392 382900 480
rect 383292 420 383348 12572
rect 383852 6804 383908 196588
rect 383852 6738 383908 6748
rect 383964 4452 384020 200088
rect 384860 4564 384916 200088
rect 385756 196644 385812 200088
rect 386652 196756 386708 200088
rect 386652 196690 386708 196700
rect 385756 196578 385812 196588
rect 384860 4498 384916 4508
rect 386540 52164 386596 52174
rect 383964 4386 384020 4396
rect 384412 480 384580 532
rect 386540 480 386596 52108
rect 387548 5012 387604 200088
rect 388444 195748 388500 200088
rect 388444 195682 388500 195692
rect 387548 4946 387604 4956
rect 389340 4788 389396 200088
rect 390236 20188 390292 200088
rect 390572 198212 390628 198222
rect 390572 52164 390628 198156
rect 390572 52098 390628 52108
rect 390236 20132 390404 20188
rect 389340 4722 389396 4732
rect 390236 12964 390292 12974
rect 388556 4228 388612 4238
rect 388556 480 388612 4172
rect 384412 476 384776 480
rect 384412 420 384468 476
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 383292 364 384468 420
rect 384524 392 384776 476
rect 384552 -960 384776 392
rect 386456 -960 386680 480
rect 388360 392 388612 480
rect 390236 480 390292 12908
rect 390348 4340 390404 20132
rect 391132 12628 391188 200088
rect 392028 198212 392084 200088
rect 392028 198146 392084 198156
rect 392252 198212 392308 198222
rect 392252 12964 392308 198156
rect 392252 12898 392308 12908
rect 391132 12562 391188 12572
rect 390348 4274 390404 4284
rect 392364 4340 392420 4350
rect 392364 480 392420 4284
rect 392924 4228 392980 200088
rect 393820 198212 393876 200088
rect 393820 198146 393876 198156
rect 394716 4340 394772 200088
rect 394716 4274 394772 4284
rect 394828 196644 394884 196654
rect 392924 4162 392980 4172
rect 394268 4228 394324 4238
rect 394268 480 394324 4172
rect 390236 392 390488 480
rect 388360 -960 388584 392
rect 390264 -960 390488 392
rect 392168 392 392420 480
rect 394072 392 394324 480
rect 394828 420 394884 196588
rect 395612 4228 395668 200088
rect 396508 196644 396564 200088
rect 396508 196578 396564 196588
rect 395612 4162 395668 4172
rect 395836 480 396004 532
rect 395836 476 396200 480
rect 395836 420 395892 476
rect 392168 -960 392392 392
rect 394072 -960 394296 392
rect 394828 364 395892 420
rect 395948 392 396200 476
rect 395976 -960 396200 392
rect 397404 420 397460 200088
rect 398300 197428 398356 200088
rect 399196 198212 399252 200088
rect 399196 198146 399252 198156
rect 398300 197362 398356 197372
rect 399868 197428 399924 197438
rect 397740 480 397908 532
rect 399868 480 399924 197372
rect 400092 197316 400148 200088
rect 400092 197250 400148 197260
rect 400652 198212 400708 198222
rect 400652 4228 400708 198156
rect 400988 198212 401044 200088
rect 400988 198146 401044 198156
rect 400652 4162 400708 4172
rect 401660 4228 401716 4238
rect 401660 480 401716 4172
rect 401884 4116 401940 200088
rect 402332 197316 402388 197326
rect 402332 4228 402388 197260
rect 402780 4788 402836 200088
rect 402780 4722 402836 4732
rect 402332 4162 402388 4172
rect 403564 4228 403620 4238
rect 401884 4050 401940 4060
rect 403564 480 403620 4172
rect 403676 4004 403732 200088
rect 404012 198212 404068 198222
rect 404012 4452 404068 198156
rect 404572 197092 404628 200088
rect 405468 197428 405524 200088
rect 405468 197362 405524 197372
rect 404572 197026 404628 197036
rect 405692 197092 405748 197102
rect 405692 5908 405748 197036
rect 405692 5842 405748 5852
rect 404012 4386 404068 4396
rect 405468 4452 405524 4462
rect 403676 3938 403732 3948
rect 405468 480 405524 4396
rect 406364 4452 406420 200088
rect 406364 4386 406420 4396
rect 407260 4340 407316 200088
rect 408156 4676 408212 200088
rect 408156 4610 408212 4620
rect 407260 4274 407316 4284
rect 409052 4228 409108 200088
rect 409948 8036 410004 200088
rect 409948 7970 410004 7980
rect 409052 4162 409108 4172
rect 409276 4788 409332 4798
rect 407372 4116 407428 4126
rect 407372 480 407428 4060
rect 409276 480 409332 4732
rect 410844 4564 410900 200088
rect 411740 198100 411796 200088
rect 411740 198034 411796 198044
rect 412412 197428 412468 197438
rect 412412 5796 412468 197372
rect 412636 196756 412692 200088
rect 413532 196980 413588 200088
rect 413532 196914 413588 196924
rect 414092 198100 414148 198110
rect 412636 196690 412692 196700
rect 414092 6020 414148 198044
rect 414428 12628 414484 200088
rect 414428 12562 414484 12572
rect 414092 5954 414148 5964
rect 412412 5730 412468 5740
rect 413084 5908 413140 5918
rect 410844 4498 410900 4508
rect 411180 4004 411236 4014
rect 411180 480 411236 3948
rect 413084 480 413140 5852
rect 415324 5908 415380 200088
rect 416220 197652 416276 200088
rect 416220 197586 416276 197596
rect 415772 196980 415828 196990
rect 415772 7588 415828 196924
rect 415772 7522 415828 7532
rect 415324 5842 415380 5852
rect 414988 5796 415044 5806
rect 414988 480 415044 5740
rect 416892 4452 416948 4462
rect 416892 480 416948 4396
rect 417116 4452 417172 200088
rect 418012 196644 418068 200088
rect 418012 196578 418068 196588
rect 418908 15988 418964 200088
rect 418908 15922 418964 15932
rect 417116 4386 417172 4396
rect 418796 4340 418852 4350
rect 418796 480 418852 4284
rect 419804 4340 419860 200088
rect 420700 197540 420756 200088
rect 420700 197474 420756 197484
rect 421596 196588 421652 200088
rect 422492 198100 422548 200088
rect 422492 198034 422548 198044
rect 422492 196756 422548 196766
rect 421596 196532 421764 196588
rect 421708 195860 421764 196532
rect 421708 195794 421764 195804
rect 422492 6132 422548 196700
rect 422716 196644 422772 196654
rect 422716 9380 422772 196588
rect 422716 9314 422772 9324
rect 423388 7812 423444 200088
rect 424284 197876 424340 200088
rect 424284 197810 424340 197820
rect 423388 7746 423444 7756
rect 424508 8036 424564 8046
rect 422492 6066 422548 6076
rect 419804 4274 419860 4284
rect 420700 4676 420756 4686
rect 420700 480 420756 4620
rect 422604 4228 422660 4238
rect 422604 480 422660 4172
rect 424508 480 424564 7980
rect 425180 4228 425236 200088
rect 426076 9268 426132 200088
rect 426972 21028 427028 200088
rect 426972 20962 427028 20972
rect 427868 11060 427924 200088
rect 427868 10994 427924 11004
rect 428764 10948 428820 200088
rect 429660 37828 429716 200088
rect 430556 61348 430612 200088
rect 430556 61282 430612 61292
rect 430892 198100 430948 198110
rect 429660 37762 429716 37772
rect 428764 10882 428820 10892
rect 426076 9202 426132 9212
rect 430220 6132 430276 6142
rect 428428 6020 428484 6030
rect 425180 4162 425236 4172
rect 426412 4564 426468 4574
rect 426412 480 426468 4508
rect 428428 480 428484 5964
rect 430220 480 430276 6076
rect 430892 6020 430948 198044
rect 431452 197428 431508 200088
rect 431452 197362 431508 197372
rect 432348 51268 432404 200088
rect 432348 51202 432404 51212
rect 430892 5954 430948 5964
rect 432124 7588 432180 7598
rect 432124 480 432180 7532
rect 433244 6132 433300 200088
rect 434140 14308 434196 200088
rect 434140 14242 434196 14252
rect 433244 6066 433300 6076
rect 433468 12628 433524 12638
rect 397740 476 398104 480
rect 397740 420 397796 476
rect 397404 364 397796 420
rect 397852 392 398104 476
rect 397880 -960 398104 392
rect 399784 -960 400008 480
rect 401660 392 401912 480
rect 403564 392 403816 480
rect 405468 392 405720 480
rect 407372 392 407624 480
rect 409276 392 409528 480
rect 411180 392 411432 480
rect 413084 392 413336 480
rect 414988 392 415240 480
rect 416892 392 417144 480
rect 418796 392 419048 480
rect 420700 392 420952 480
rect 422604 392 422856 480
rect 424508 392 424760 480
rect 426412 392 426664 480
rect 401688 -960 401912 392
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 407400 -960 407624 392
rect 409304 -960 409528 392
rect 411208 -960 411432 392
rect 413112 -960 413336 392
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418824 -960 419048 392
rect 420728 -960 420952 392
rect 422632 -960 422856 392
rect 424536 -960 424760 392
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430220 392 430472 480
rect 432124 392 432376 480
rect 430248 -960 430472 392
rect 432152 -960 432376 392
rect 433468 420 433524 12572
rect 435036 12628 435092 200088
rect 435932 198212 435988 200088
rect 436856 200060 437556 200116
rect 435932 198146 435988 198156
rect 437500 197764 437556 200060
rect 437500 197698 437556 197708
rect 435036 12562 435092 12572
rect 436828 197652 436884 197662
rect 435932 5908 435988 5918
rect 433916 480 434084 532
rect 435932 480 435988 5852
rect 433916 476 434280 480
rect 433916 420 433972 476
rect 433468 364 433972 420
rect 434028 392 434280 476
rect 435932 392 436184 480
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 436828 420 436884 197596
rect 437724 120148 437780 200088
rect 438396 198212 438452 198222
rect 438396 189028 438452 198156
rect 438620 198100 438676 200088
rect 439544 200060 440132 200116
rect 438620 198034 438676 198044
rect 440076 196588 440132 200060
rect 440076 196532 440244 196588
rect 440188 195748 440244 196532
rect 440188 195682 440244 195692
rect 438396 188962 438452 188972
rect 437724 120082 437780 120092
rect 440412 7700 440468 200088
rect 441308 24388 441364 200088
rect 442204 187460 442260 200088
rect 442204 187394 442260 187404
rect 441308 24322 441364 24332
rect 443100 22708 443156 200088
rect 443996 192612 444052 200088
rect 443996 192546 444052 192556
rect 444332 197876 444388 197886
rect 443100 22642 443156 22652
rect 444332 17556 444388 197820
rect 444892 135268 444948 200088
rect 445788 165508 445844 200088
rect 446684 197652 446740 200088
rect 447580 197988 447636 200088
rect 447580 197922 447636 197932
rect 446684 197586 446740 197596
rect 445788 165442 445844 165452
rect 446012 197540 446068 197550
rect 444892 135202 444948 135212
rect 444332 17490 444388 17500
rect 443548 15988 443604 15998
rect 440412 7634 440468 7644
rect 441644 9380 441700 9390
rect 439740 4452 439796 4462
rect 437724 480 437892 532
rect 439740 480 439796 4396
rect 441644 480 441700 9324
rect 443548 480 443604 15932
rect 446012 6804 446068 197484
rect 448476 7588 448532 200088
rect 448476 7522 448532 7532
rect 448588 195860 448644 195870
rect 446012 6738 446068 6748
rect 447356 6804 447412 6814
rect 445452 4340 445508 4350
rect 445452 480 445508 4284
rect 447356 480 447412 6748
rect 437724 476 438088 480
rect 437724 420 437780 476
rect 436828 364 437780 420
rect 437836 392 438088 476
rect 439740 392 439992 480
rect 441644 392 441896 480
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 447356 392 447608 480
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 447384 -960 447608 392
rect 448588 420 448644 195804
rect 449372 123508 449428 200088
rect 450268 197876 450324 200088
rect 450268 197810 450324 197820
rect 449372 123442 449428 123452
rect 451164 20188 451220 200088
rect 452060 195972 452116 200088
rect 452956 197540 453012 200088
rect 452956 197474 453012 197484
rect 452060 195906 452116 195916
rect 451164 20132 451444 20188
rect 451164 6020 451220 6030
rect 449148 480 449316 532
rect 451164 480 451220 5964
rect 451388 6020 451444 20132
rect 453852 19348 453908 200088
rect 453852 19282 453908 19292
rect 454412 198100 454468 198110
rect 454412 17668 454468 198044
rect 454748 196980 454804 200088
rect 454748 196914 454804 196924
rect 455644 192500 455700 200088
rect 455644 192434 455700 192444
rect 456092 196980 456148 196990
rect 454412 17602 454468 17612
rect 453628 17556 453684 17566
rect 451388 5954 451444 5964
rect 453068 7812 453124 7822
rect 453068 480 453124 7756
rect 449148 476 449512 480
rect 449148 420 449204 476
rect 448588 364 449204 420
rect 449260 392 449512 476
rect 451164 392 451416 480
rect 453068 392 453320 480
rect 449288 -960 449512 392
rect 451192 -960 451416 392
rect 453096 -960 453320 392
rect 453628 420 453684 17500
rect 456092 5908 456148 196924
rect 456540 190820 456596 200088
rect 456540 190754 456596 190764
rect 457436 178948 457492 200088
rect 458332 194180 458388 200088
rect 458332 194114 458388 194124
rect 457436 178882 457492 178892
rect 456092 5842 456148 5852
rect 458780 9268 458836 9278
rect 456988 4228 457044 4238
rect 454860 480 455028 532
rect 456988 480 457044 4172
rect 458780 480 458836 9212
rect 459228 9268 459284 200088
rect 460124 177268 460180 200088
rect 461020 185668 461076 200088
rect 461020 185602 461076 185612
rect 460124 177202 460180 177212
rect 459228 9202 459284 9212
rect 460348 21028 460404 21038
rect 454860 476 455224 480
rect 454860 420 454916 476
rect 453628 364 454916 420
rect 454972 392 455224 476
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 458808 -960 459032 392
rect 460348 420 460404 20972
rect 461916 15988 461972 200088
rect 461916 15922 461972 15932
rect 462588 11060 462644 11070
rect 460572 480 460740 532
rect 462588 480 462644 11004
rect 462812 4676 462868 200088
rect 463708 183988 463764 200088
rect 463708 183922 463764 183932
rect 464604 21028 464660 200088
rect 464604 20962 464660 20972
rect 465388 37828 465444 37838
rect 462812 4610 462868 4620
rect 464492 10948 464548 10958
rect 464492 480 464548 10892
rect 460572 476 460936 480
rect 460572 420 460628 476
rect 460348 364 460628 420
rect 460684 392 460936 476
rect 462588 392 462840 480
rect 464492 392 464744 480
rect 460712 -960 460936 392
rect 462616 -960 462840 392
rect 464520 -960 464744 392
rect 465388 420 465444 37772
rect 465500 4564 465556 200088
rect 466396 187348 466452 200088
rect 466396 187282 466452 187292
rect 467292 180628 467348 200088
rect 467292 180562 467348 180572
rect 467852 197652 467908 197662
rect 467852 10948 467908 197596
rect 467852 10882 467908 10892
rect 465500 4498 465556 4508
rect 468188 4452 468244 200088
rect 469084 195860 469140 200088
rect 469084 195794 469140 195804
rect 468860 61348 468916 61358
rect 468748 29428 468804 29438
rect 468748 7028 468804 29372
rect 468748 6962 468804 6972
rect 468188 4386 468244 4396
rect 468860 3780 468916 61292
rect 469980 54628 470036 200088
rect 470876 197092 470932 200088
rect 471772 198212 471828 200088
rect 471772 198146 471828 198156
rect 470876 197026 470932 197036
rect 472668 194068 472724 200088
rect 472668 194002 472724 194012
rect 472892 198212 472948 198222
rect 472892 182308 472948 198156
rect 472892 182242 472948 182252
rect 469980 54562 470036 54572
rect 472108 51268 472164 51278
rect 468524 3724 468916 3780
rect 469532 7028 469588 7038
rect 466284 480 466452 532
rect 468524 480 468580 3724
rect 466284 476 466648 480
rect 466284 420 466340 476
rect 465388 364 466340 420
rect 466396 392 466648 476
rect 466424 -960 466648 392
rect 468328 392 468580 480
rect 469532 420 469588 6972
rect 470092 480 470260 532
rect 472108 480 472164 51212
rect 473564 4340 473620 200088
rect 474460 199220 474516 200088
rect 474460 199154 474516 199164
rect 475356 199108 475412 200088
rect 475356 199042 475412 199052
rect 475468 14308 475524 14318
rect 473564 4274 473620 4284
rect 474012 6132 474068 6142
rect 474012 480 474068 6076
rect 470092 476 470456 480
rect 470092 420 470148 476
rect 468328 -960 468552 392
rect 469532 364 470148 420
rect 470204 392 470456 476
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475468 420 475524 14252
rect 476252 4228 476308 200088
rect 477148 192388 477204 200088
rect 477148 192322 477204 192332
rect 478044 14308 478100 200088
rect 478940 198212 478996 200088
rect 478940 198146 478996 198156
rect 478940 197428 478996 197438
rect 478044 14242 478100 14252
rect 478828 189028 478884 189038
rect 476252 4162 476308 4172
rect 477148 12628 477204 12638
rect 475804 480 475972 532
rect 475804 476 476168 480
rect 475804 420 475860 476
rect 475468 364 475860 420
rect 475916 392 476168 476
rect 475944 -960 476168 392
rect 477148 420 477204 12572
rect 477708 480 477876 532
rect 477708 476 478072 480
rect 477708 420 477764 476
rect 477148 364 477764 420
rect 477820 392 478072 476
rect 477848 -960 478072 392
rect 478828 420 478884 188972
rect 478940 29428 478996 197372
rect 479052 197092 479108 197102
rect 479052 189140 479108 197036
rect 479836 190708 479892 200088
rect 479836 190642 479892 190652
rect 479052 189074 479108 189084
rect 480732 189028 480788 200088
rect 480732 188962 480788 188972
rect 478940 29362 478996 29372
rect 481628 12628 481684 200088
rect 482524 197652 482580 200088
rect 482524 197586 482580 197596
rect 481628 12562 481684 12572
rect 482188 120148 482244 120158
rect 481852 11620 481908 11630
rect 479612 480 479780 532
rect 481852 480 481908 11564
rect 479612 476 479976 480
rect 479612 420 479668 476
rect 478828 364 479668 420
rect 479724 392 479976 476
rect 479752 -960 479976 392
rect 481656 392 481908 480
rect 482188 420 482244 120092
rect 483420 29428 483476 200088
rect 483420 29362 483476 29372
rect 483868 197764 483924 197774
rect 483868 11620 483924 197708
rect 484316 197428 484372 200088
rect 488012 198212 488068 198222
rect 484316 197362 484372 197372
rect 486332 197988 486388 197998
rect 486332 36148 486388 197932
rect 486332 36082 486388 36092
rect 487228 195748 487284 195758
rect 487228 20188 487284 195692
rect 488012 195748 488068 198156
rect 488012 195682 488068 195692
rect 494732 197876 494788 197886
rect 491372 187460 491428 187470
rect 490588 24388 490644 24398
rect 487228 20132 487396 20188
rect 483868 11554 483924 11564
rect 485548 17668 485604 17678
rect 483420 480 483588 532
rect 485548 480 485604 17612
rect 487340 480 487396 20132
rect 489244 7700 489300 7710
rect 489244 480 489300 7644
rect 483420 476 483784 480
rect 483420 420 483476 476
rect 481656 -960 481880 392
rect 482188 364 483476 420
rect 483532 392 483784 476
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487340 392 487592 480
rect 489244 392 489496 480
rect 487368 -960 487592 392
rect 489272 -960 489496 392
rect 490588 420 490644 24332
rect 491372 4788 491428 187404
rect 493948 22708 494004 22718
rect 491372 4722 491428 4732
rect 493052 4788 493108 4798
rect 491036 480 491204 532
rect 493052 480 493108 4732
rect 491036 476 491400 480
rect 491036 420 491092 476
rect 490588 364 491092 420
rect 491148 392 491400 476
rect 493052 392 493304 480
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 493948 420 494004 22652
rect 494732 22708 494788 197820
rect 494732 22642 494788 22652
rect 495628 192612 495684 192622
rect 494844 480 495012 532
rect 494844 476 495208 480
rect 494844 420 494900 476
rect 493948 364 494900 420
rect 494956 392 495208 476
rect 494984 -960 495208 392
rect 495628 420 495684 192556
rect 498988 163044 499044 498988
rect 499100 495684 499156 501116
rect 499100 495618 499156 495628
rect 498988 162978 499044 162988
rect 499772 165508 499828 165518
rect 497308 135268 497364 135278
rect 496748 480 496916 532
rect 496748 476 497112 480
rect 496748 420 496804 476
rect 495628 364 496804 420
rect 496860 392 497112 476
rect 496888 -960 497112 392
rect 497308 420 497364 135212
rect 499772 4116 499828 165452
rect 500668 121044 500724 502572
rect 504028 502404 504084 502414
rect 502348 501060 502404 501070
rect 500668 120978 500724 120988
rect 501452 123508 501508 123518
rect 501452 4788 501508 123452
rect 502348 79044 502404 501004
rect 502348 78978 502404 78988
rect 504028 41188 504084 502348
rect 506492 362964 506548 506156
rect 512428 502964 512484 502974
rect 506492 362898 506548 362908
rect 509068 502516 509124 502526
rect 504028 41122 504084 41132
rect 506492 197540 506548 197550
rect 504028 36148 504084 36158
rect 501452 4722 501508 4732
rect 502572 10948 502628 10958
rect 499772 4050 499828 4060
rect 500668 4116 500724 4126
rect 498652 480 498820 532
rect 500668 480 500724 4060
rect 502572 480 502628 10892
rect 498652 476 499016 480
rect 498652 420 498708 476
rect 497308 364 498708 420
rect 498764 392 499016 476
rect 500668 392 500920 480
rect 502572 392 502824 480
rect 498792 -960 499016 392
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504028 420 504084 36092
rect 506492 32676 506548 197484
rect 509068 94948 509124 502460
rect 509068 94882 509124 94892
rect 506492 32610 506548 32620
rect 512428 27748 512484 502908
rect 514108 502740 514164 502750
rect 513212 499268 513268 499278
rect 513212 430164 513268 499212
rect 513212 430098 513268 430108
rect 512428 27682 512484 27692
rect 514108 26068 514164 502684
rect 514892 500948 514948 500958
rect 514892 468804 514948 500892
rect 514892 468738 514948 468748
rect 516572 112644 516628 509180
rect 518252 151284 518308 512540
rect 519932 231924 519988 521052
rect 521612 509348 521668 509358
rect 521612 270564 521668 509292
rect 523292 310884 523348 525980
rect 539308 519988 539364 595644
rect 540428 595476 540484 595644
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584696 595672 584920 597000
rect 584696 595560 584948 595672
rect 540540 595476 540596 595560
rect 540428 595420 540596 595476
rect 560252 591220 560308 591230
rect 560252 538468 560308 591164
rect 562604 591220 562660 595560
rect 562604 591154 562660 591164
rect 584892 590212 584948 595560
rect 584892 590146 584948 590156
rect 593180 590212 593236 590222
rect 560252 538402 560308 538412
rect 593068 588644 593124 588654
rect 593068 535108 593124 588588
rect 593068 535042 593124 535052
rect 539308 519922 539364 519932
rect 593068 525924 593124 525934
rect 536732 519428 536788 519438
rect 526652 514500 526708 514510
rect 526652 349524 526708 514444
rect 533372 512708 533428 512718
rect 531692 505876 531748 505886
rect 531692 389844 531748 505820
rect 533372 416724 533428 512652
rect 535052 504420 535108 504430
rect 535052 455364 535108 504364
rect 535052 455298 535108 455308
rect 533372 416658 533428 416668
rect 531692 389778 531748 389788
rect 526652 349458 526708 349468
rect 523292 310818 523348 310828
rect 521612 270498 521668 270508
rect 519932 231858 519988 231868
rect 536732 218484 536788 519372
rect 540092 519316 540148 519326
rect 536732 218418 536788 218428
rect 538412 516068 538468 516078
rect 531692 197652 531748 197662
rect 519148 195972 519204 195982
rect 518252 151218 518308 151228
rect 518364 178948 518420 178958
rect 516572 112578 516628 112588
rect 514108 26002 514164 26012
rect 515788 32676 515844 32686
rect 509068 22708 509124 22718
rect 506380 7588 506436 7598
rect 504364 480 504532 532
rect 506380 480 506436 7532
rect 508284 4788 508340 4798
rect 508284 480 508340 4732
rect 504364 476 504728 480
rect 504364 420 504420 476
rect 504028 364 504420 420
rect 504476 392 504728 476
rect 506380 392 506632 480
rect 508284 392 508536 480
rect 504504 -960 504728 392
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 509068 420 509124 22652
rect 515788 20188 515844 32620
rect 515788 20132 515956 20188
rect 512092 6020 512148 6030
rect 510076 480 510244 532
rect 512092 480 512148 5964
rect 514220 3668 514276 3678
rect 514220 480 514276 3612
rect 510076 476 510440 480
rect 510076 420 510132 476
rect 509068 364 510132 420
rect 510188 392 510440 476
rect 512092 392 512344 480
rect 510216 -960 510440 392
rect 512120 -960 512344 392
rect 514024 392 514276 480
rect 515900 480 515956 20132
rect 517468 19348 517524 19358
rect 515900 392 516152 480
rect 514024 -960 514248 392
rect 515928 -960 516152 392
rect 517468 420 517524 19292
rect 518364 4116 518420 178892
rect 518364 4050 518420 4060
rect 519148 3668 519204 195916
rect 525868 194180 525924 194190
rect 520828 192500 520884 192510
rect 519148 3602 519204 3612
rect 519708 5908 519764 5918
rect 517692 480 517860 532
rect 519708 480 519764 5852
rect 517692 476 518056 480
rect 517692 420 517748 476
rect 517468 364 517748 420
rect 517804 392 518056 476
rect 519708 392 519960 480
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 520828 420 520884 192444
rect 522508 190820 522564 190830
rect 521500 480 521668 532
rect 521500 476 521864 480
rect 521500 420 521556 476
rect 520828 364 521556 420
rect 521612 392 521864 476
rect 521640 -960 521864 392
rect 522508 420 522564 190764
rect 525420 4116 525476 4126
rect 523404 480 523572 532
rect 525420 480 525476 4060
rect 523404 476 523768 480
rect 523404 420 523460 476
rect 522508 364 523460 420
rect 523516 392 523768 476
rect 525420 392 525672 480
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 525868 420 525924 194124
rect 531692 26068 531748 197596
rect 531692 26002 531748 26012
rect 532588 185668 532644 185678
rect 529228 9268 529284 9278
rect 527212 480 527380 532
rect 529228 480 529284 9212
rect 531356 4116 531412 4126
rect 531356 480 531412 4060
rect 527212 476 527576 480
rect 527212 420 527268 476
rect 525868 364 527268 420
rect 527324 392 527576 476
rect 529228 392 529480 480
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 392 531412 480
rect 532588 420 532644 185612
rect 536732 183988 536788 183998
rect 534268 177268 534324 177278
rect 534268 4116 534324 177212
rect 534268 4050 534324 4060
rect 534380 15988 534436 15998
rect 532924 480 533092 532
rect 532924 476 533288 480
rect 532924 420 532980 476
rect 531160 -960 531384 392
rect 532588 364 532980 420
rect 533036 392 533288 476
rect 533064 -960 533288 392
rect 534380 420 534436 15932
rect 536732 5012 536788 183932
rect 538412 99204 538468 516012
rect 540092 137844 540148 519260
rect 550172 517860 550228 517870
rect 541772 510916 541828 510926
rect 541772 178164 541828 510860
rect 548492 502852 548548 502862
rect 545132 500836 545188 500846
rect 545132 297444 545188 500780
rect 548492 336084 548548 502796
rect 550172 376404 550228 517804
rect 550172 376338 550228 376348
rect 588812 517524 588868 517534
rect 548492 336018 548548 336028
rect 545132 297378 545188 297388
rect 588812 258468 588868 517468
rect 588812 258402 588868 258412
rect 590492 515844 590548 515854
rect 560252 199220 560308 199230
rect 549388 195860 549444 195870
rect 544348 187348 544404 187358
rect 541772 178098 541828 178108
rect 541884 180628 541940 180638
rect 540092 137778 540148 137788
rect 538412 99138 538468 99148
rect 539308 21028 539364 21038
rect 536732 4946 536788 4956
rect 538748 5012 538804 5022
rect 536844 4676 536900 4686
rect 534828 480 534996 532
rect 536844 480 536900 4620
rect 538748 480 538804 4956
rect 534828 476 535192 480
rect 534828 420 534884 476
rect 534380 364 534884 420
rect 534940 392 535192 476
rect 536844 392 537096 480
rect 538748 392 539000 480
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 538776 -960 539000 392
rect 539308 420 539364 20972
rect 540204 4452 540260 4462
rect 540204 4116 540260 4396
rect 541884 4452 541940 180572
rect 544348 20188 544404 187292
rect 544348 20132 544516 20188
rect 541884 4386 541940 4396
rect 542668 4564 542724 4574
rect 540204 4050 540260 4060
rect 540540 480 540708 532
rect 542668 480 542724 4508
rect 544460 480 544516 20132
rect 546364 4452 546420 4462
rect 546364 480 546420 4396
rect 548268 4116 548324 4126
rect 548268 480 548324 4060
rect 540540 476 540904 480
rect 540540 420 540596 476
rect 539308 364 540596 420
rect 540652 392 540904 476
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 549388 420 549444 195804
rect 557788 194068 557844 194078
rect 552748 189140 552804 189150
rect 551068 54628 551124 54638
rect 550060 480 550228 532
rect 550060 476 550424 480
rect 550060 420 550116 476
rect 549388 364 550116 420
rect 550172 392 550424 476
rect 550200 -960 550424 392
rect 551068 420 551124 54572
rect 551964 480 552132 532
rect 551964 476 552328 480
rect 551964 420 552020 476
rect 551068 364 552020 420
rect 552076 392 552328 476
rect 552104 -960 552328 392
rect 552748 420 552804 189084
rect 554428 182308 554484 182318
rect 553868 480 554036 532
rect 553868 476 554232 480
rect 553868 420 553924 476
rect 552748 364 553924 420
rect 553980 392 554232 476
rect 554008 -960 554232 392
rect 554428 420 554484 182252
rect 555772 480 555940 532
rect 557788 480 557844 194012
rect 560252 5012 560308 199164
rect 570332 197428 570388 197438
rect 567868 14308 567924 14318
rect 560252 4946 560308 4956
rect 561596 5012 561652 5022
rect 559692 4340 559748 4350
rect 559692 480 559748 4284
rect 561596 480 561652 4956
rect 563724 4340 563780 4350
rect 563724 480 563780 4284
rect 555772 476 556136 480
rect 555772 420 555828 476
rect 554428 364 555828 420
rect 555884 392 556136 476
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 563528 392 563780 480
rect 565404 4228 565460 4238
rect 565404 480 565460 4172
rect 567532 4228 567588 4238
rect 567532 480 567588 4172
rect 565404 392 565656 480
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 567336 392 567588 480
rect 567868 420 567924 14252
rect 570332 4452 570388 197372
rect 570332 4386 570388 4396
rect 571228 195748 571284 195758
rect 569100 480 569268 532
rect 571228 480 571284 195692
rect 590492 192388 590548 515788
rect 593068 205604 593124 525868
rect 593180 525028 593236 590156
rect 593180 524962 593236 524972
rect 593292 529396 593348 529406
rect 593068 205538 593124 205548
rect 593180 520996 593236 521006
rect 590492 192322 590548 192332
rect 593068 199108 593124 199118
rect 572908 190708 572964 190718
rect 572908 20188 572964 190652
rect 574588 189028 574644 189038
rect 572908 20132 573076 20188
rect 573020 480 573076 20132
rect 569100 476 569464 480
rect 569100 420 569156 476
rect 567336 -960 567560 392
rect 567868 364 569156 420
rect 569212 392 569464 476
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 573048 -960 573272 392
rect 574588 420 574644 188972
rect 590492 34468 590548 34478
rect 581308 29428 581364 29438
rect 579628 26068 579684 26078
rect 576268 12628 576324 12638
rect 574812 480 574980 532
rect 574812 476 575176 480
rect 574812 420 574868 476
rect 574588 364 574868 420
rect 574924 392 575176 476
rect 574952 -960 575176 392
rect 576268 420 576324 12572
rect 576716 480 576884 532
rect 576716 476 577080 480
rect 576716 420 576772 476
rect 576268 364 576772 420
rect 576828 392 577080 476
rect 576856 -960 577080 392
rect 578760 -960 578984 480
rect 579628 420 579684 26012
rect 580524 480 580692 532
rect 580524 476 580888 480
rect 580524 420 580580 476
rect 579628 364 580580 420
rect 580636 392 580888 476
rect 580664 -960 580888 392
rect 581308 420 581364 29372
rect 590492 20580 590548 34412
rect 590492 20514 590548 20524
rect 584444 4452 584500 4462
rect 582428 480 582596 532
rect 584444 480 584500 4396
rect 593068 4340 593124 199052
rect 593180 7364 593236 520940
rect 593292 33796 593348 529340
rect 593852 527716 593908 527726
rect 593516 524244 593572 524254
rect 593404 504196 593460 504206
rect 593404 47012 593460 504140
rect 593516 73444 593572 524188
rect 593628 514276 593684 514286
rect 593628 86660 593684 514220
rect 593740 500724 593796 500734
rect 593740 126308 593796 500668
rect 593852 165956 593908 527660
rect 593964 522788 594020 522798
rect 593964 245252 594020 522732
rect 594524 511028 594580 511038
rect 594412 507668 594468 507678
rect 594300 505764 594356 505774
rect 594076 504308 594132 504318
rect 594076 284900 594132 504252
rect 594188 499156 594244 499166
rect 594188 324548 594244 499100
rect 594300 403844 594356 505708
rect 594412 443492 594468 507612
rect 594524 483140 594580 510972
rect 594524 483074 594580 483084
rect 594412 443426 594468 443436
rect 594300 403778 594356 403788
rect 594188 324482 594244 324492
rect 594076 284834 594132 284844
rect 593964 245186 594020 245196
rect 593852 165890 593908 165900
rect 593964 192276 594020 192286
rect 593740 126242 593796 126252
rect 593628 86594 593684 86604
rect 593516 73378 593572 73388
rect 593404 46946 593460 46956
rect 593292 33730 593348 33740
rect 593180 7298 593236 7308
rect 593068 4274 593124 4284
rect 593964 4228 594020 192220
rect 593964 4162 594020 4172
rect 582428 476 582792 480
rect 582428 420 582484 476
rect 581308 364 582484 420
rect 582540 392 582792 476
rect 584444 392 584696 480
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 9212 520828 9268 520884
rect 4172 516572 4228 516628
rect 4172 503132 4228 503188
rect 5852 502460 5908 502516
rect 5852 501452 5908 501508
rect 14252 586348 14308 586404
rect 55356 593068 55412 593124
rect 31948 583772 32004 583828
rect 14252 565292 14308 565348
rect 27692 530908 27748 530964
rect 10108 503244 10164 503300
rect 12572 527548 12628 527604
rect 22652 519148 22708 519204
rect 19292 514108 19348 514164
rect 12572 275548 12628 275604
rect 14252 510748 14308 510804
rect 17612 504028 17668 504084
rect 15932 498988 15988 499044
rect 17612 473788 17668 473844
rect 15932 458668 15988 458724
rect 22652 361228 22708 361284
rect 19292 317548 19348 317604
rect 14252 262108 14308 262164
rect 9212 206332 9268 206388
rect 10108 195692 10164 195748
rect 4172 94892 4228 94948
rect 4172 93436 4228 93492
rect 4172 41132 4228 41188
rect 4172 36876 4228 36932
rect 4284 27692 4340 27748
rect 4172 26012 4228 26068
rect 4284 22876 4340 22932
rect 4172 8764 4228 8820
rect 22652 192332 22708 192388
rect 11788 31052 11844 31108
rect 18508 12572 18564 12628
rect 17276 6188 17332 6244
rect 15372 4956 15428 5012
rect 187740 593180 187796 593236
rect 165676 590156 165732 590212
rect 167132 590156 167188 590212
rect 143612 585452 143668 585508
rect 99148 550172 99204 550228
rect 77308 526652 77364 526708
rect 167132 551852 167188 551908
rect 120988 525084 121044 525140
rect 206668 529340 206724 529396
rect 44492 522508 44548 522564
rect 203308 520940 203364 520996
rect 158732 517692 158788 517748
rect 155372 517580 155428 517636
rect 98252 507500 98308 507556
rect 98252 487228 98308 487284
rect 44492 233548 44548 233604
rect 144508 199164 144564 199220
rect 65548 199052 65604 199108
rect 57036 195804 57092 195860
rect 27692 191548 27748 191604
rect 29372 194012 29428 194068
rect 27692 190652 27748 190708
rect 22652 4956 22708 5012
rect 24892 9212 24948 9268
rect 22988 4284 23044 4340
rect 21084 4060 21140 4116
rect 27692 4284 27748 4340
rect 28700 4284 28756 4340
rect 26796 4172 26852 4228
rect 36988 189084 37044 189140
rect 31948 188972 32004 189028
rect 30268 44492 30324 44548
rect 29372 4172 29428 4228
rect 33628 14252 33684 14308
rect 36316 4396 36372 4452
rect 45388 187292 45444 187348
rect 41132 178892 41188 178948
rect 40124 4060 40180 4116
rect 44492 56252 44548 56308
rect 41132 4060 41188 4116
rect 41916 4956 41972 5012
rect 47068 180572 47124 180628
rect 44492 4956 44548 5012
rect 43932 4508 43988 4564
rect 52108 160412 52164 160468
rect 48748 52892 48804 52948
rect 51548 4620 51604 4676
rect 53788 54572 53844 54628
rect 62972 165452 63028 165508
rect 58828 158732 58884 158788
rect 62860 4732 62916 4788
rect 61068 4060 61124 4116
rect 62972 4060 63028 4116
rect 63868 157052 63924 157108
rect 113372 197484 113428 197540
rect 94892 197372 94948 197428
rect 80668 185612 80724 185668
rect 72268 182252 72324 182308
rect 71372 167132 71428 167188
rect 68012 61292 68068 61348
rect 68012 4732 68068 4788
rect 68908 37772 68964 37828
rect 68684 4060 68740 4116
rect 71372 4060 71428 4116
rect 75628 155372 75684 155428
rect 74396 4060 74452 4116
rect 78092 66332 78148 66388
rect 78092 4060 78148 4116
rect 78204 7532 78260 7588
rect 80108 4060 80164 4116
rect 89068 183932 89124 183988
rect 87388 175532 87444 175588
rect 84812 146972 84868 147028
rect 82348 17612 82404 17668
rect 84812 4060 84868 4116
rect 85820 4732 85876 4788
rect 90748 32844 90804 32900
rect 93436 5068 93492 5124
rect 104188 194124 104244 194180
rect 97468 192444 97524 192500
rect 94892 5068 94948 5124
rect 95340 5964 95396 6020
rect 97244 4060 97300 4116
rect 99932 185724 99988 185780
rect 99932 4060 99988 4116
rect 100828 153692 100884 153748
rect 102956 10892 103012 10948
rect 105868 184044 105924 184100
rect 109228 173852 109284 173908
rect 107548 148652 107604 148708
rect 132636 195916 132692 195972
rect 117628 182364 117684 182420
rect 115948 172172 116004 172228
rect 113372 12572 113428 12628
rect 113484 24332 113540 24388
rect 112476 4060 112532 4116
rect 113484 4060 113540 4116
rect 114380 2492 114436 2548
rect 120988 170492 121044 170548
rect 119308 42924 119364 42980
rect 126028 168812 126084 168868
rect 124348 19292 124404 19348
rect 122668 15932 122724 15988
rect 129276 152012 129332 152068
rect 131068 20972 131124 21028
rect 137788 194236 137844 194292
rect 134428 187404 134484 187460
rect 136108 177212 136164 177268
rect 139468 182476 139524 182532
rect 142828 179004 142884 179060
rect 142716 173964 142772 174020
rect 142716 4060 142772 4116
rect 154476 190764 154532 190820
rect 149436 167244 149492 167300
rect 147868 17724 147924 17780
rect 146524 4060 146580 4116
rect 151228 29372 151284 29428
rect 149436 4956 149492 5012
rect 150332 4956 150388 5012
rect 154364 9324 154420 9380
rect 157052 515900 157108 515956
rect 157052 105868 157108 105924
rect 157948 150332 158004 150388
rect 155372 63868 155428 63924
rect 154476 4060 154532 4116
rect 156044 4060 156100 4116
rect 163772 516124 163828 516180
rect 185612 514332 185668 514388
rect 173852 512428 173908 512484
rect 167132 509404 167188 509460
rect 167132 445228 167188 445284
rect 170492 507388 170548 507444
rect 163772 403228 163828 403284
rect 162988 180684 163044 180740
rect 158732 149548 158788 149604
rect 161308 165564 161364 165620
rect 159852 12572 159908 12628
rect 166348 162092 166404 162148
rect 165788 7644 165844 7700
rect 173068 135212 173124 135268
rect 170492 50428 170548 50484
rect 171388 93212 171444 93268
rect 170492 49532 170548 49588
rect 169596 4060 169652 4116
rect 170492 4060 170548 4116
rect 178892 507724 178948 507780
rect 178108 189196 178164 189252
rect 173852 134428 173908 134484
rect 174748 177324 174804 177380
rect 176428 22652 176484 22708
rect 182252 506044 182308 506100
rect 180572 505932 180628 505988
rect 182252 388108 182308 388164
rect 180572 346108 180628 346164
rect 190652 512764 190708 512820
rect 188972 502460 189028 502516
rect 192332 511084 192388 511140
rect 190652 431788 190708 431844
rect 191436 500668 191492 500724
rect 188972 304108 189028 304164
rect 185612 220108 185668 220164
rect 178892 176428 178948 176484
rect 179788 198268 179844 198324
rect 182252 197820 182308 197876
rect 181468 21084 181524 21140
rect 182252 9212 182308 9268
rect 185612 175644 185668 175700
rect 184716 4956 184772 5012
rect 188972 172284 189028 172340
rect 185612 4956 185668 5012
rect 188412 16044 188468 16100
rect 186732 4060 186788 4116
rect 197372 509516 197428 509572
rect 194012 507836 194068 507892
rect 195692 504476 195748 504532
rect 195692 374668 195748 374724
rect 194012 332668 194068 332724
rect 199836 502348 199892 502404
rect 199052 501004 199108 501060
rect 199052 416668 199108 416724
rect 197372 290668 197428 290724
rect 192332 246988 192388 247044
rect 197372 197932 197428 197988
rect 191436 58828 191492 58884
rect 194012 192556 194068 192612
rect 191548 47852 191604 47908
rect 188972 4060 189028 4116
rect 190540 4060 190596 4116
rect 193228 37884 193284 37940
rect 194012 4060 194068 4116
rect 194908 179116 194964 179172
rect 197372 44492 197428 44548
rect 196588 36092 196644 36148
rect 208348 523292 208404 523348
rect 213388 524188 213444 524244
rect 223468 516012 223524 516068
rect 218428 514220 218484 514276
rect 212156 504140 212212 504196
rect 209580 502348 209636 502404
rect 217308 500668 217364 500724
rect 221788 509180 221844 509236
rect 253932 591276 253988 591332
rect 257852 591276 257908 591332
rect 275996 591276 276052 591332
rect 279692 591276 279748 591332
rect 319228 578732 319284 578788
rect 297388 543452 297444 543508
rect 314972 561148 315028 561204
rect 279692 536732 279748 536788
rect 257852 535164 257908 535220
rect 311612 535948 311668 536004
rect 307468 531804 307524 531860
rect 235228 527660 235284 527716
rect 231868 519260 231924 519316
rect 230188 503468 230244 503524
rect 230300 512540 230356 512596
rect 227612 500668 227668 500724
rect 260428 525980 260484 526036
rect 241948 525868 242004 525924
rect 239372 515788 239428 515844
rect 237916 503916 237972 503972
rect 250348 522732 250404 522788
rect 245308 521052 245364 521108
rect 239372 503916 239428 503972
rect 240268 510860 240324 510916
rect 246988 519372 247044 519428
rect 255388 517468 255444 517524
rect 252588 509292 252644 509348
rect 258524 504252 258580 504308
rect 304108 522620 304164 522676
rect 278908 517804 278964 517860
rect 268828 514444 268884 514500
rect 263676 500780 263732 500836
rect 273868 506156 273924 506212
rect 271404 502796 271460 502852
rect 275772 505820 275828 505876
rect 286076 512652 286132 512708
rect 280924 505708 280980 505764
rect 296380 510972 296436 511028
rect 288988 507612 289044 507668
rect 294588 504364 294644 504420
rect 292012 500892 292068 500948
rect 299068 509068 299124 509124
rect 302316 501116 302372 501172
rect 310044 503916 310100 503972
rect 314188 535052 314244 535108
rect 311612 503916 311668 503972
rect 312620 504588 312676 504644
rect 333452 547708 333508 547764
rect 324268 538412 324324 538468
rect 314972 504588 315028 504644
rect 317548 528332 317604 528388
rect 319228 524972 319284 525028
rect 322588 519932 322644 519988
rect 327628 533372 327684 533428
rect 339388 541772 339444 541828
rect 333452 531804 333508 531860
rect 334348 540092 334404 540148
rect 332668 531692 332724 531748
rect 330652 503356 330708 503412
rect 362012 590492 362068 590548
rect 351148 578732 351204 578788
rect 343532 574588 343588 574644
rect 341068 521276 341124 521332
rect 342748 528444 342804 528500
rect 338380 503580 338436 503636
rect 343532 528332 343588 528388
rect 346108 521276 346164 521332
rect 348684 503692 348740 503748
rect 356188 543452 356244 543508
rect 352828 536732 352884 536788
rect 357868 535164 357924 535220
rect 362012 528444 362068 528500
rect 361228 523292 361284 523348
rect 365372 593180 365428 593236
rect 380492 593068 380548 593124
rect 367948 585452 368004 585508
rect 371308 551852 371364 551908
rect 365372 503916 365428 503972
rect 366716 503916 366772 503972
rect 362908 503692 362964 503748
rect 364140 503468 364196 503524
rect 378028 550172 378084 550228
rect 376348 526652 376404 526708
rect 372988 525084 373044 525140
rect 386092 590492 386148 590548
rect 386428 583772 386484 583828
rect 394828 572908 394884 572964
rect 389788 565292 389844 565348
rect 380492 503916 380548 503972
rect 382172 503916 382228 503972
rect 384748 503244 384804 503300
rect 391468 557788 391524 557844
rect 393932 529228 393988 529284
rect 393932 514892 393988 514948
rect 396508 544348 396564 544404
rect 401548 514892 401604 514948
rect 400204 503132 400260 503188
rect 407932 504028 407988 504084
rect 405356 501452 405412 501508
rect 451052 590156 451108 590212
rect 430108 541772 430164 541828
rect 452284 590156 452340 590212
rect 451052 540092 451108 540148
rect 463708 530908 463764 530964
rect 448588 527548 448644 527604
rect 433468 519148 433524 519204
rect 425068 516124 425124 516180
rect 414988 512764 415044 512820
rect 408268 503580 408324 503636
rect 409948 507500 410004 507556
rect 417452 509404 417508 509460
rect 423388 506044 423444 506100
rect 420812 501004 420868 501060
rect 430332 505932 430388 505988
rect 428540 504476 428596 504532
rect 440188 514108 440244 514164
rect 435484 507836 435540 507892
rect 438844 502460 438900 502516
rect 445788 510748 445844 510804
rect 443548 509516 443604 509572
rect 455308 522508 455364 522564
rect 453628 514332 453684 514388
rect 450940 511084 450996 511140
rect 458668 520828 458724 520884
rect 472108 517692 472164 517748
rect 462028 507724 462084 507780
rect 468972 512428 469028 512484
rect 517468 533372 517524 533428
rect 495628 531692 495684 531748
rect 523292 525980 523348 526036
rect 519932 521052 519988 521108
rect 487228 517580 487284 517636
rect 478828 515900 478884 515956
rect 473788 503356 473844 503412
rect 474908 502572 474964 502628
rect 477484 502460 477540 502516
rect 484428 507388 484484 507444
rect 482636 501004 482692 501060
rect 518252 512540 518308 512596
rect 516572 509180 516628 509236
rect 506492 506156 506548 506212
rect 495516 502908 495572 502964
rect 492940 502684 492996 502740
rect 490364 502348 490420 502404
rect 500668 502572 500724 502628
rect 499100 501116 499156 501172
rect 467180 499324 467236 499380
rect 266252 499212 266308 499268
rect 284284 499212 284340 499268
rect 413084 499212 413140 499268
rect 498988 498988 499044 499044
rect 212828 198156 212884 198212
rect 209916 197596 209972 197652
rect 206668 190876 206724 190932
rect 199836 34412 199892 34468
rect 201628 187516 201684 187572
rect 199836 31164 199892 31220
rect 203308 185836 203364 185892
rect 205772 4060 205828 4116
rect 207452 51212 207508 51268
rect 207452 4060 207508 4116
rect 208348 39452 208404 39508
rect 211708 196028 211764 196084
rect 209916 25116 209972 25172
rect 210028 194348 210084 194404
rect 215516 198156 215572 198212
rect 212828 195692 212884 195748
rect 214956 197260 215012 197316
rect 217308 192332 217364 192388
rect 216412 31052 216468 31108
rect 214956 5068 215012 5124
rect 215068 25116 215124 25172
rect 219100 197484 219156 197540
rect 218204 6188 218260 6244
rect 217196 5740 217252 5796
rect 218876 5068 218932 5124
rect 219996 4172 220052 4228
rect 220108 195692 220164 195748
rect 221788 197708 221844 197764
rect 222684 194012 222740 194068
rect 220892 190652 220948 190708
rect 224476 197932 224532 197988
rect 223692 197708 223748 197764
rect 223692 197260 223748 197316
rect 224252 197484 224308 197540
rect 225372 188972 225428 189028
rect 224252 157052 224308 157108
rect 223580 4284 223636 4340
rect 225932 29484 225988 29540
rect 224812 4172 224868 4228
rect 222908 2604 222964 2660
rect 226268 14252 226324 14308
rect 225932 4172 225988 4228
rect 226716 11004 226772 11060
rect 228060 189084 228116 189140
rect 228956 178892 229012 178948
rect 229852 56252 229908 56308
rect 230300 44492 230356 44548
rect 227164 4396 227220 4452
rect 228508 19404 228564 19460
rect 231644 187292 231700 187348
rect 232540 180572 232596 180628
rect 233436 52892 233492 52948
rect 230748 4508 230804 4564
rect 231868 46172 231924 46228
rect 234332 198156 234388 198212
rect 235228 160412 235284 160468
rect 234332 158732 234388 158788
rect 237916 198156 237972 198212
rect 237020 195804 237076 195860
rect 238812 165452 238868 165508
rect 241500 199052 241556 199108
rect 240604 197484 240660 197540
rect 241948 197484 242004 197540
rect 241948 194348 242004 194404
rect 242396 167132 242452 167188
rect 239708 61292 239764 61348
rect 236124 54572 236180 54628
rect 244188 182252 244244 182308
rect 245980 155372 246036 155428
rect 245084 66332 245140 66388
rect 243292 37772 243348 37828
rect 243628 31052 243684 31108
rect 233548 4620 233604 4676
rect 233660 24444 233716 24500
rect 238588 12684 238644 12740
rect 236236 7756 236292 7812
rect 238140 6076 238196 6132
rect 241836 2716 241892 2772
rect 246876 7532 246932 7588
rect 246988 192332 247044 192388
rect 248668 185612 248724 185668
rect 247772 146972 247828 147028
rect 248668 184156 248724 184212
rect 245868 28 245924 84
rect 249564 17612 249620 17668
rect 251356 175532 251412 175588
rect 252028 188972 252084 189028
rect 250460 4732 250516 4788
rect 251468 4172 251524 4228
rect 252252 183932 252308 183988
rect 254044 197372 254100 197428
rect 254492 197372 254548 197428
rect 253708 196588 253764 196644
rect 253708 192444 253764 192500
rect 254492 184044 254548 184100
rect 253148 32844 253204 32900
rect 252812 32732 252868 32788
rect 252812 4172 252868 4228
rect 253820 17612 253876 17668
rect 256732 196588 256788 196644
rect 257068 197148 257124 197204
rect 257068 194124 257124 194180
rect 255836 185724 255892 185780
rect 257628 153692 257684 153748
rect 254940 5964 254996 6020
rect 257180 14476 257236 14532
rect 260316 197372 260372 197428
rect 259420 197148 259476 197204
rect 260428 148652 260484 148708
rect 261212 194012 261268 194068
rect 258524 10892 258580 10948
rect 260988 9212 261044 9268
rect 259084 4172 259140 4228
rect 262108 173852 262164 173908
rect 263004 24332 263060 24388
rect 261212 4172 261268 4228
rect 262108 14588 262164 14644
rect 264572 197372 264628 197428
rect 264572 187404 264628 187460
rect 265692 182364 265748 182420
rect 264796 172172 264852 172228
rect 267484 170492 267540 170548
rect 266588 42924 266644 42980
rect 266252 42812 266308 42868
rect 265468 21196 265524 21252
rect 263788 2492 263844 2548
rect 264796 4172 264852 4228
rect 270172 168812 270228 168868
rect 271068 152012 271124 152068
rect 273756 197372 273812 197428
rect 272860 195916 272916 195972
rect 273868 177212 273924 177268
rect 274652 197372 274708 197428
rect 271964 20972 272020 21028
rect 269276 19292 269332 19348
rect 268380 15932 268436 15988
rect 266252 4172 266308 4228
rect 267148 14364 267204 14420
rect 274316 9436 274372 9492
rect 270396 6748 270452 6804
rect 272412 4172 272468 4228
rect 275436 194236 275492 194292
rect 276444 182476 276500 182532
rect 278236 199164 278292 199220
rect 277340 179004 277396 179060
rect 279132 173964 279188 174020
rect 274652 6748 274708 6804
rect 274764 32844 274820 32900
rect 279020 22764 279076 22820
rect 277228 12796 277284 12852
rect 274764 4172 274820 4228
rect 276220 7532 276276 7588
rect 280924 167244 280980 167300
rect 281820 29372 281876 29428
rect 280028 17724 280084 17780
rect 281932 10892 281988 10948
rect 283052 196700 283108 196756
rect 283612 190764 283668 190820
rect 284508 150332 284564 150388
rect 283052 93212 283108 93268
rect 285404 12572 285460 12628
rect 285628 180908 285684 180964
rect 282716 9324 282772 9380
rect 283836 5964 283892 6020
rect 287196 180684 287252 180740
rect 286300 165564 286356 165620
rect 288092 196588 288148 196644
rect 288988 162092 289044 162148
rect 288092 135212 288148 135268
rect 290780 196700 290836 196756
rect 291676 196588 291732 196644
rect 292348 198156 292404 198212
rect 292348 189196 292404 189252
rect 292572 177324 292628 177380
rect 289884 49532 289940 49588
rect 294588 198268 294644 198324
rect 294364 198156 294420 198212
rect 293468 22652 293524 22708
rect 297052 175644 297108 175700
rect 297948 172284 298004 172340
rect 296156 21084 296212 21140
rect 297500 24332 297556 24388
rect 292348 19292 292404 19348
rect 287308 7644 287364 7700
rect 287420 16156 287476 16212
rect 289548 11228 289604 11284
rect 291452 7644 291508 7700
rect 295708 12572 295764 12628
rect 295260 2492 295316 2548
rect 299740 192556 299796 192612
rect 300636 47852 300692 47908
rect 300860 197932 300916 197988
rect 300860 196028 300916 196084
rect 302428 179116 302484 179172
rect 300748 37884 300804 37940
rect 298844 16044 298900 16100
rect 300972 37772 301028 37828
rect 303324 36092 303380 36148
rect 305116 187516 305172 187572
rect 306012 185836 306068 185892
rect 307804 190876 307860 190932
rect 308252 197820 308308 197876
rect 306908 51212 306964 51268
rect 304220 31164 304276 31220
rect 305788 36092 305844 36148
rect 302428 29596 302484 29652
rect 304108 17724 304164 17780
rect 310492 197932 310548 197988
rect 311388 197596 311444 197652
rect 309596 197484 309652 197540
rect 311612 197484 311668 197540
rect 308700 39452 308756 39508
rect 308252 16156 308308 16212
rect 307468 15932 307524 15988
rect 311612 11228 311668 11284
rect 310492 6188 310548 6244
rect 313180 197708 313236 197764
rect 314076 195692 314132 195748
rect 312284 5852 312340 5908
rect 312396 11116 312452 11172
rect 314972 198156 315028 198212
rect 314188 2604 314244 2660
rect 314300 3500 314356 3556
rect 315868 29484 315924 29540
rect 316652 20972 316708 21028
rect 314972 2716 315028 2772
rect 316204 7868 316260 7924
rect 319452 46172 319508 46228
rect 318556 44492 318612 44548
rect 320348 24444 320404 24500
rect 317548 19404 317604 19460
rect 317884 19404 317940 19460
rect 316764 11004 316820 11060
rect 316652 3500 316708 3556
rect 321244 7756 321300 7812
rect 322140 6076 322196 6132
rect 322700 16044 322756 16100
rect 321916 5852 321972 5908
rect 320012 4172 320068 4228
rect 323932 198156 323988 198212
rect 323372 197708 323428 197764
rect 323372 14476 323428 14532
rect 323036 12684 323092 12740
rect 324380 196588 324436 196644
rect 324380 192332 324436 192388
rect 326620 196588 326676 196644
rect 327516 184156 327572 184212
rect 327628 32732 327684 32788
rect 328412 197596 328468 197652
rect 324828 31052 324884 31108
rect 327516 5068 327572 5124
rect 325724 4956 325780 5012
rect 329308 188972 329364 189028
rect 329532 195692 329588 195748
rect 328412 5068 328468 5124
rect 331100 197708 331156 197764
rect 331996 194012 332052 194068
rect 330204 17612 330260 17668
rect 334684 42812 334740 42868
rect 333788 14588 333844 14644
rect 334460 29372 334516 29428
rect 332892 9212 332948 9268
rect 333116 14252 333172 14308
rect 331436 4396 331492 4452
rect 324268 28 324324 84
rect 335580 21196 335636 21252
rect 336812 197708 336868 197764
rect 337372 197372 337428 197428
rect 338268 32844 338324 32900
rect 336812 29596 336868 29652
rect 336476 14364 336532 14420
rect 339052 11004 339108 11060
rect 337148 4508 337204 4564
rect 340060 197372 340116 197428
rect 340172 198044 340228 198100
rect 339164 9436 339220 9492
rect 339500 32732 339556 32788
rect 341068 22764 341124 22820
rect 341852 198156 341908 198212
rect 340956 12796 341012 12852
rect 342748 198156 342804 198212
rect 343532 197036 343588 197092
rect 343532 19292 343588 19348
rect 341852 10892 341908 10948
rect 343756 198156 343812 198212
rect 344540 198156 344596 198212
rect 345436 197820 345492 197876
rect 346332 197484 346388 197540
rect 343756 180908 343812 180964
rect 346108 195804 346164 195860
rect 343644 5964 343700 6020
rect 344764 5964 344820 6020
rect 340172 2492 340228 2548
rect 342860 4620 342916 4676
rect 349020 198044 349076 198100
rect 348124 197036 348180 197092
rect 347228 7644 347284 7700
rect 349580 19292 349636 19348
rect 348572 4732 348628 4788
rect 351708 37772 351764 37828
rect 351932 197932 351988 197988
rect 350812 24332 350868 24388
rect 351148 31052 351204 31108
rect 349916 12572 349972 12628
rect 352604 197708 352660 197764
rect 354620 197932 354676 197988
rect 355292 198156 355348 198212
rect 354396 36092 354452 36148
rect 354508 197372 354564 197428
rect 353500 17724 353556 17780
rect 351932 15932 351988 15988
rect 354508 7532 354564 7588
rect 356188 198156 356244 198212
rect 356972 197036 357028 197092
rect 357084 11116 357140 11172
rect 357868 195916 357924 195972
rect 356972 7868 357028 7924
rect 355292 6188 355348 6244
rect 356076 7532 356132 7588
rect 354284 4844 354340 4900
rect 358876 197036 358932 197092
rect 359548 197372 359604 197428
rect 357980 20972 358036 21028
rect 359772 19404 359828 19460
rect 362460 16044 362516 16100
rect 361228 5852 361284 5908
rect 361676 15932 361732 15988
rect 360668 4172 360724 4228
rect 364252 197596 364308 197652
rect 365148 195692 365204 195748
rect 365372 197708 365428 197764
rect 365372 32732 365428 32788
rect 363356 4956 363412 5012
rect 365708 8428 365764 8484
rect 363804 4284 363860 4340
rect 367836 198156 367892 198212
rect 368060 14252 368116 14308
rect 370524 197708 370580 197764
rect 369628 11004 369684 11060
rect 370412 197260 370468 197316
rect 370412 5964 370468 6020
rect 371420 198156 371476 198212
rect 372316 197260 372372 197316
rect 373212 195804 373268 195860
rect 373772 198156 373828 198212
rect 373772 31052 373828 31108
rect 371420 29372 371476 29428
rect 371308 4620 371364 4676
rect 373324 6748 373380 6804
rect 368732 4508 368788 4564
rect 371420 4508 371476 4564
rect 366044 4396 366100 4452
rect 369516 4396 369572 4452
rect 367612 4172 367668 4228
rect 375900 198156 375956 198212
rect 375004 19292 375060 19348
rect 375452 198044 375508 198100
rect 374108 4732 374164 4788
rect 375228 8764 375284 8820
rect 375452 8428 375508 8484
rect 378588 195916 378644 195972
rect 378812 198156 378868 198212
rect 377692 7532 377748 7588
rect 378028 195692 378084 195748
rect 376796 4844 376852 4900
rect 377132 4956 377188 5012
rect 379708 198156 379764 198212
rect 379484 197372 379540 197428
rect 378812 15932 378868 15988
rect 382172 198044 382228 198100
rect 380492 196700 380548 196756
rect 380492 8764 380548 8820
rect 379820 4284 379876 4340
rect 380940 4732 380996 4788
rect 382844 4284 382900 4340
rect 383852 196588 383908 196644
rect 383068 4172 383124 4228
rect 383292 12572 383348 12628
rect 383852 6748 383908 6804
rect 386652 196700 386708 196756
rect 385756 196588 385812 196644
rect 384860 4508 384916 4564
rect 386540 52108 386596 52164
rect 383964 4396 384020 4452
rect 388444 195692 388500 195748
rect 387548 4956 387604 5012
rect 390572 198156 390628 198212
rect 390572 52108 390628 52164
rect 389340 4732 389396 4788
rect 390236 12908 390292 12964
rect 388556 4172 388612 4228
rect 392028 198156 392084 198212
rect 392252 198156 392308 198212
rect 392252 12908 392308 12964
rect 391132 12572 391188 12628
rect 390348 4284 390404 4340
rect 392364 4284 392420 4340
rect 393820 198156 393876 198212
rect 394716 4284 394772 4340
rect 394828 196588 394884 196644
rect 392924 4172 392980 4228
rect 394268 4172 394324 4228
rect 396508 196588 396564 196644
rect 395612 4172 395668 4228
rect 399196 198156 399252 198212
rect 398300 197372 398356 197428
rect 399868 197372 399924 197428
rect 400092 197260 400148 197316
rect 400652 198156 400708 198212
rect 400988 198156 401044 198212
rect 400652 4172 400708 4228
rect 401660 4172 401716 4228
rect 402332 197260 402388 197316
rect 402780 4732 402836 4788
rect 402332 4172 402388 4228
rect 403564 4172 403620 4228
rect 401884 4060 401940 4116
rect 404012 198156 404068 198212
rect 405468 197372 405524 197428
rect 404572 197036 404628 197092
rect 405692 197036 405748 197092
rect 405692 5852 405748 5908
rect 404012 4396 404068 4452
rect 405468 4396 405524 4452
rect 403676 3948 403732 4004
rect 406364 4396 406420 4452
rect 408156 4620 408212 4676
rect 407260 4284 407316 4340
rect 409948 7980 410004 8036
rect 409052 4172 409108 4228
rect 409276 4732 409332 4788
rect 407372 4060 407428 4116
rect 411740 198044 411796 198100
rect 412412 197372 412468 197428
rect 413532 196924 413588 196980
rect 414092 198044 414148 198100
rect 412636 196700 412692 196756
rect 414428 12572 414484 12628
rect 414092 5964 414148 6020
rect 412412 5740 412468 5796
rect 413084 5852 413140 5908
rect 410844 4508 410900 4564
rect 411180 3948 411236 4004
rect 416220 197596 416276 197652
rect 415772 196924 415828 196980
rect 415772 7532 415828 7588
rect 415324 5852 415380 5908
rect 414988 5740 415044 5796
rect 416892 4396 416948 4452
rect 418012 196588 418068 196644
rect 418908 15932 418964 15988
rect 417116 4396 417172 4452
rect 418796 4284 418852 4340
rect 420700 197484 420756 197540
rect 422492 198044 422548 198100
rect 422492 196700 422548 196756
rect 421708 195804 421764 195860
rect 422716 196588 422772 196644
rect 422716 9324 422772 9380
rect 424284 197820 424340 197876
rect 423388 7756 423444 7812
rect 424508 7980 424564 8036
rect 422492 6076 422548 6132
rect 419804 4284 419860 4340
rect 420700 4620 420756 4676
rect 422604 4172 422660 4228
rect 426972 20972 427028 21028
rect 427868 11004 427924 11060
rect 430556 61292 430612 61348
rect 430892 198044 430948 198100
rect 429660 37772 429716 37828
rect 428764 10892 428820 10948
rect 426076 9212 426132 9268
rect 430220 6076 430276 6132
rect 428428 5964 428484 6020
rect 425180 4172 425236 4228
rect 426412 4508 426468 4564
rect 431452 197372 431508 197428
rect 432348 51212 432404 51268
rect 430892 5964 430948 6020
rect 432124 7532 432180 7588
rect 434140 14252 434196 14308
rect 433244 6076 433300 6132
rect 433468 12572 433524 12628
rect 435932 198156 435988 198212
rect 437500 197708 437556 197764
rect 435036 12572 435092 12628
rect 436828 197596 436884 197652
rect 435932 5852 435988 5908
rect 438396 198156 438452 198212
rect 438620 198044 438676 198100
rect 440188 195692 440244 195748
rect 438396 188972 438452 189028
rect 437724 120092 437780 120148
rect 442204 187404 442260 187460
rect 441308 24332 441364 24388
rect 443996 192556 444052 192612
rect 444332 197820 444388 197876
rect 443100 22652 443156 22708
rect 447580 197932 447636 197988
rect 446684 197596 446740 197652
rect 445788 165452 445844 165508
rect 446012 197484 446068 197540
rect 444892 135212 444948 135268
rect 444332 17500 444388 17556
rect 443548 15932 443604 15988
rect 440412 7644 440468 7700
rect 441644 9324 441700 9380
rect 439740 4396 439796 4452
rect 448476 7532 448532 7588
rect 448588 195804 448644 195860
rect 446012 6748 446068 6804
rect 447356 6748 447412 6804
rect 445452 4284 445508 4340
rect 450268 197820 450324 197876
rect 449372 123452 449428 123508
rect 452956 197484 453012 197540
rect 452060 195916 452116 195972
rect 451164 5964 451220 6020
rect 453852 19292 453908 19348
rect 454412 198044 454468 198100
rect 454748 196924 454804 196980
rect 455644 192444 455700 192500
rect 456092 196924 456148 196980
rect 454412 17612 454468 17668
rect 453628 17500 453684 17556
rect 451388 5964 451444 6020
rect 453068 7756 453124 7812
rect 456540 190764 456596 190820
rect 458332 194124 458388 194180
rect 457436 178892 457492 178948
rect 456092 5852 456148 5908
rect 458780 9212 458836 9268
rect 456988 4172 457044 4228
rect 461020 185612 461076 185668
rect 460124 177212 460180 177268
rect 459228 9212 459284 9268
rect 460348 20972 460404 21028
rect 461916 15932 461972 15988
rect 462588 11004 462644 11060
rect 463708 183932 463764 183988
rect 464604 20972 464660 21028
rect 465388 37772 465444 37828
rect 462812 4620 462868 4676
rect 464492 10892 464548 10948
rect 466396 187292 466452 187348
rect 467292 180572 467348 180628
rect 467852 197596 467908 197652
rect 467852 10892 467908 10948
rect 465500 4508 465556 4564
rect 469084 195804 469140 195860
rect 468860 61292 468916 61348
rect 468748 29372 468804 29428
rect 468748 6972 468804 7028
rect 468188 4396 468244 4452
rect 471772 198156 471828 198212
rect 470876 197036 470932 197092
rect 472668 194012 472724 194068
rect 472892 198156 472948 198212
rect 472892 182252 472948 182308
rect 469980 54572 470036 54628
rect 472108 51212 472164 51268
rect 469532 6972 469588 7028
rect 474460 199164 474516 199220
rect 475356 199052 475412 199108
rect 475468 14252 475524 14308
rect 473564 4284 473620 4340
rect 474012 6076 474068 6132
rect 477148 192332 477204 192388
rect 478940 198156 478996 198212
rect 478940 197372 478996 197428
rect 478044 14252 478100 14308
rect 478828 188972 478884 189028
rect 476252 4172 476308 4228
rect 477148 12572 477204 12628
rect 479052 197036 479108 197092
rect 479836 190652 479892 190708
rect 479052 189084 479108 189140
rect 480732 188972 480788 189028
rect 478940 29372 478996 29428
rect 482524 197596 482580 197652
rect 481628 12572 481684 12628
rect 482188 120092 482244 120148
rect 481852 11564 481908 11620
rect 483420 29372 483476 29428
rect 483868 197708 483924 197764
rect 488012 198156 488068 198212
rect 484316 197372 484372 197428
rect 486332 197932 486388 197988
rect 486332 36092 486388 36148
rect 487228 195692 487284 195748
rect 488012 195692 488068 195748
rect 494732 197820 494788 197876
rect 491372 187404 491428 187460
rect 490588 24332 490644 24388
rect 483868 11564 483924 11620
rect 485548 17612 485604 17668
rect 489244 7644 489300 7700
rect 493948 22652 494004 22708
rect 491372 4732 491428 4788
rect 493052 4732 493108 4788
rect 494732 22652 494788 22708
rect 495628 192556 495684 192612
rect 499100 495628 499156 495684
rect 498988 162988 499044 163044
rect 499772 165452 499828 165508
rect 497308 135212 497364 135268
rect 504028 502348 504084 502404
rect 502348 501004 502404 501060
rect 500668 120988 500724 121044
rect 501452 123452 501508 123508
rect 502348 78988 502404 79044
rect 512428 502908 512484 502964
rect 506492 362908 506548 362964
rect 509068 502460 509124 502516
rect 504028 41132 504084 41188
rect 506492 197484 506548 197540
rect 504028 36092 504084 36148
rect 501452 4732 501508 4788
rect 502572 10892 502628 10948
rect 499772 4060 499828 4116
rect 500668 4060 500724 4116
rect 509068 94892 509124 94948
rect 506492 32620 506548 32676
rect 514108 502684 514164 502740
rect 513212 499212 513268 499268
rect 513212 430108 513268 430164
rect 512428 27692 512484 27748
rect 514892 500892 514948 500948
rect 514892 468748 514948 468804
rect 521612 509292 521668 509348
rect 560252 591164 560308 591220
rect 562604 591164 562660 591220
rect 584892 590156 584948 590212
rect 593180 590156 593236 590212
rect 560252 538412 560308 538468
rect 593068 588588 593124 588644
rect 593068 535052 593124 535108
rect 539308 519932 539364 519988
rect 593068 525868 593124 525924
rect 536732 519372 536788 519428
rect 526652 514444 526708 514500
rect 533372 512652 533428 512708
rect 531692 505820 531748 505876
rect 535052 504364 535108 504420
rect 535052 455308 535108 455364
rect 533372 416668 533428 416724
rect 531692 389788 531748 389844
rect 526652 349468 526708 349524
rect 523292 310828 523348 310884
rect 521612 270508 521668 270564
rect 519932 231868 519988 231924
rect 540092 519260 540148 519316
rect 536732 218428 536788 218484
rect 538412 516012 538468 516068
rect 531692 197596 531748 197652
rect 519148 195916 519204 195972
rect 518252 151228 518308 151284
rect 518364 178892 518420 178948
rect 516572 112588 516628 112644
rect 514108 26012 514164 26068
rect 515788 32620 515844 32676
rect 509068 22652 509124 22708
rect 506380 7532 506436 7588
rect 508284 4732 508340 4788
rect 512092 5964 512148 6020
rect 514220 3612 514276 3668
rect 517468 19292 517524 19348
rect 518364 4060 518420 4116
rect 525868 194124 525924 194180
rect 520828 192444 520884 192500
rect 519148 3612 519204 3668
rect 519708 5852 519764 5908
rect 522508 190764 522564 190820
rect 525420 4060 525476 4116
rect 531692 26012 531748 26068
rect 532588 185612 532644 185668
rect 529228 9212 529284 9268
rect 531356 4060 531412 4116
rect 536732 183932 536788 183988
rect 534268 177212 534324 177268
rect 534268 4060 534324 4116
rect 534380 15932 534436 15988
rect 550172 517804 550228 517860
rect 541772 510860 541828 510916
rect 548492 502796 548548 502852
rect 545132 500780 545188 500836
rect 550172 376348 550228 376404
rect 588812 517468 588868 517524
rect 548492 336028 548548 336084
rect 545132 297388 545188 297444
rect 588812 258412 588868 258468
rect 590492 515788 590548 515844
rect 560252 199164 560308 199220
rect 549388 195804 549444 195860
rect 544348 187292 544404 187348
rect 541772 178108 541828 178164
rect 541884 180572 541940 180628
rect 540092 137788 540148 137844
rect 538412 99148 538468 99204
rect 539308 20972 539364 21028
rect 536732 4956 536788 5012
rect 538748 4956 538804 5012
rect 536844 4620 536900 4676
rect 540204 4396 540260 4452
rect 541884 4396 541940 4452
rect 542668 4508 542724 4564
rect 540204 4060 540260 4116
rect 546364 4396 546420 4452
rect 548268 4060 548324 4116
rect 557788 194012 557844 194068
rect 552748 189084 552804 189140
rect 551068 54572 551124 54628
rect 554428 182252 554484 182308
rect 570332 197372 570388 197428
rect 567868 14252 567924 14308
rect 560252 4956 560308 5012
rect 561596 4956 561652 5012
rect 559692 4284 559748 4340
rect 563724 4284 563780 4340
rect 565404 4172 565460 4228
rect 567532 4172 567588 4228
rect 570332 4396 570388 4452
rect 571228 195692 571284 195748
rect 593180 524972 593236 525028
rect 593292 529340 593348 529396
rect 593068 205548 593124 205604
rect 593180 520940 593236 520996
rect 590492 192332 590548 192388
rect 593068 199052 593124 199108
rect 572908 190652 572964 190708
rect 574588 188972 574644 189028
rect 590492 34412 590548 34468
rect 581308 29372 581364 29428
rect 579628 26012 579684 26068
rect 576268 12572 576324 12628
rect 590492 20524 590548 20580
rect 584444 4396 584500 4452
rect 593852 527660 593908 527716
rect 593516 524188 593572 524244
rect 593404 504140 593460 504196
rect 593628 514220 593684 514276
rect 593740 500668 593796 500724
rect 593964 522732 594020 522788
rect 594524 510972 594580 511028
rect 594412 507612 594468 507668
rect 594300 505708 594356 505764
rect 594076 504252 594132 504308
rect 594188 499100 594244 499156
rect 594524 483084 594580 483140
rect 594412 443436 594468 443492
rect 594300 403788 594356 403844
rect 594188 324492 594244 324548
rect 594076 284844 594132 284900
rect 593964 245196 594020 245252
rect 593852 165900 593908 165956
rect 593964 192220 594020 192276
rect 593740 126252 593796 126308
rect 593628 86604 593684 86660
rect 593516 73388 593572 73444
rect 593404 46956 593460 47012
rect 593292 33740 593348 33796
rect 593180 7308 593236 7364
rect 593068 4284 593124 4340
rect 593964 4172 594020 4228
<< metal3 >>
rect 187730 593180 187740 593236
rect 187796 593180 365372 593236
rect 365428 593180 365438 593236
rect 55346 593068 55356 593124
rect 55412 593068 380492 593124
rect 380548 593068 380558 593124
rect 253922 591276 253932 591332
rect 253988 591276 257852 591332
rect 257908 591276 257918 591332
rect 275986 591276 275996 591332
rect 276052 591276 279692 591332
rect 279748 591276 279758 591332
rect 560242 591164 560252 591220
rect 560308 591164 562604 591220
rect 562660 591164 562670 591220
rect 362002 590492 362012 590548
rect 362068 590492 386092 590548
rect 386148 590492 386158 590548
rect 165666 590156 165676 590212
rect 165732 590156 167132 590212
rect 167188 590156 167198 590212
rect 451042 590156 451052 590212
rect 451108 590156 452284 590212
rect 452340 590156 452350 590212
rect 584882 590156 584892 590212
rect 584948 590156 593180 590212
rect 593236 590156 593246 590212
rect 595560 588644 597000 588840
rect 593058 588588 593068 588644
rect 593124 588616 597000 588644
rect 593124 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 532 587188
rect 392 587132 532 587160
rect 476 587076 532 587132
rect 364 587020 532 587076
rect 364 586404 420 587020
rect 364 586348 14252 586404
rect 14308 586348 14318 586404
rect 143602 585452 143612 585508
rect 143668 585452 367948 585508
rect 368004 585452 368014 585508
rect 31938 583772 31948 583828
rect 32004 583772 386428 583828
rect 386484 583772 386494 583828
rect 319218 578732 319228 578788
rect 319284 578732 351148 578788
rect 351204 578732 351214 578788
rect 595560 575428 597000 575624
rect 595420 575400 597000 575428
rect 595420 575372 595672 575400
rect 595420 575316 595476 575372
rect 595420 575260 595700 575316
rect 595644 574644 595700 575260
rect 343522 574588 343532 574644
rect 343588 574588 595700 574644
rect -960 573076 480 573272
rect -960 573048 8428 573076
rect 392 573020 8428 573048
rect 8372 572964 8428 573020
rect 8372 572908 394828 572964
rect 394884 572908 394894 572964
rect 14242 565292 14252 565348
rect 14308 565292 389788 565348
rect 389844 565292 389854 565348
rect 595560 562212 597000 562408
rect 595420 562184 597000 562212
rect 595420 562156 595672 562184
rect 595420 562100 595476 562156
rect 595420 562044 595700 562100
rect 595644 561204 595700 562044
rect 314962 561148 314972 561204
rect 315028 561148 595700 561204
rect -960 558964 480 559160
rect -960 558936 532 558964
rect 392 558908 532 558936
rect 476 558852 532 558908
rect 364 558796 532 558852
rect 364 557844 420 558796
rect 364 557788 391468 557844
rect 391524 557788 391534 557844
rect 167122 551852 167132 551908
rect 167188 551852 371308 551908
rect 371364 551852 371374 551908
rect 99138 550172 99148 550228
rect 99204 550172 378028 550228
rect 378084 550172 378094 550228
rect 595560 548996 597000 549192
rect 595420 548968 597000 548996
rect 595420 548940 595672 548968
rect 595420 548884 595476 548940
rect 595420 548828 595700 548884
rect 595644 547764 595700 548828
rect 333442 547708 333452 547764
rect 333508 547708 595700 547764
rect -960 544852 480 545048
rect -960 544824 532 544852
rect 392 544796 532 544824
rect 476 544740 532 544796
rect 364 544684 532 544740
rect 364 544404 420 544684
rect 364 544348 396508 544404
rect 396564 544348 396574 544404
rect 297378 543452 297388 543508
rect 297444 543452 356188 543508
rect 356244 543452 356254 543508
rect 339378 541772 339388 541828
rect 339444 541772 430108 541828
rect 430164 541772 430174 541828
rect 334338 540092 334348 540148
rect 334404 540092 451052 540148
rect 451108 540092 451118 540148
rect 324258 538412 324268 538468
rect 324324 538412 560252 538468
rect 560308 538412 560318 538468
rect 279682 536732 279692 536788
rect 279748 536732 352828 536788
rect 352884 536732 352894 536788
rect 311602 535948 311612 536004
rect 311668 535948 590212 536004
rect 590156 535892 590212 535948
rect 595560 535892 597000 535976
rect 590156 535836 597000 535892
rect 595560 535752 597000 535836
rect 257842 535164 257852 535220
rect 257908 535164 357868 535220
rect 357924 535164 357934 535220
rect 314178 535052 314188 535108
rect 314244 535052 593068 535108
rect 593124 535052 593134 535108
rect 327618 533372 327628 533428
rect 327684 533372 517468 533428
rect 517524 533372 517534 533428
rect 307458 531804 307468 531860
rect 307524 531804 333452 531860
rect 333508 531804 333518 531860
rect 332658 531692 332668 531748
rect 332724 531692 495628 531748
rect 495684 531692 495694 531748
rect -960 530740 480 530936
rect 27682 530908 27692 530964
rect 27748 530908 463708 530964
rect 463764 530908 463774 530964
rect -960 530712 532 530740
rect 392 530684 532 530712
rect 476 530628 532 530684
rect 364 530572 532 530628
rect 364 529284 420 530572
rect 206658 529340 206668 529396
rect 206724 529340 593292 529396
rect 593348 529340 593358 529396
rect 364 529228 393932 529284
rect 393988 529228 393998 529284
rect 342738 528444 342748 528500
rect 342804 528444 362012 528500
rect 362068 528444 362078 528500
rect 317538 528332 317548 528388
rect 317604 528332 343532 528388
rect 343588 528332 343598 528388
rect 235218 527660 235228 527716
rect 235284 527660 593852 527716
rect 593908 527660 593918 527716
rect 12562 527548 12572 527604
rect 12628 527548 448588 527604
rect 448644 527548 448654 527604
rect 77298 526652 77308 526708
rect 77364 526652 376348 526708
rect 376404 526652 376414 526708
rect 260418 525980 260428 526036
rect 260484 525980 523292 526036
rect 523348 525980 523358 526036
rect 241938 525868 241948 525924
rect 242004 525868 593068 525924
rect 593124 525868 593134 525924
rect 120978 525084 120988 525140
rect 121044 525084 372988 525140
rect 373044 525084 373054 525140
rect 319218 524972 319228 525028
rect 319284 524972 593180 525028
rect 593236 524972 593246 525028
rect 213378 524188 213388 524244
rect 213444 524188 593516 524244
rect 593572 524188 593582 524244
rect 208338 523292 208348 523348
rect 208404 523292 361228 523348
rect 361284 523292 361294 523348
rect 250338 522732 250348 522788
rect 250404 522732 593964 522788
rect 594020 522732 594030 522788
rect 595560 522676 597000 522760
rect 304098 522620 304108 522676
rect 304164 522620 597000 522676
rect 44482 522508 44492 522564
rect 44548 522508 455308 522564
rect 455364 522508 455374 522564
rect 595560 522536 597000 522620
rect 341058 521276 341068 521332
rect 341124 521276 346108 521332
rect 346164 521276 346174 521332
rect 245298 521052 245308 521108
rect 245364 521052 519932 521108
rect 519988 521052 519998 521108
rect 203298 520940 203308 520996
rect 203364 520940 593180 520996
rect 593236 520940 593246 520996
rect 9202 520828 9212 520884
rect 9268 520828 458668 520884
rect 458724 520828 458734 520884
rect 322578 519932 322588 519988
rect 322644 519932 539308 519988
rect 539364 519932 539374 519988
rect 246978 519372 246988 519428
rect 247044 519372 536732 519428
rect 536788 519372 536798 519428
rect 231858 519260 231868 519316
rect 231924 519260 540092 519316
rect 540148 519260 540158 519316
rect 22642 519148 22652 519204
rect 22708 519148 433468 519204
rect 433524 519148 433534 519204
rect 278898 517804 278908 517860
rect 278964 517804 550172 517860
rect 550228 517804 550238 517860
rect 158722 517692 158732 517748
rect 158788 517692 472108 517748
rect 472164 517692 472174 517748
rect 155362 517580 155372 517636
rect 155428 517580 487228 517636
rect 487284 517580 487294 517636
rect 255378 517468 255388 517524
rect 255444 517468 588812 517524
rect 588868 517468 588878 517524
rect -960 516628 480 516824
rect -960 516600 4172 516628
rect 392 516572 4172 516600
rect 4228 516572 4238 516628
rect 163762 516124 163772 516180
rect 163828 516124 425068 516180
rect 425124 516124 425134 516180
rect 223458 516012 223468 516068
rect 223524 516012 538412 516068
rect 538468 516012 538478 516068
rect 157042 515900 157052 515956
rect 157108 515900 478828 515956
rect 478884 515900 478894 515956
rect 239362 515788 239372 515844
rect 239428 515788 590492 515844
rect 590548 515788 590558 515844
rect 393922 514892 393932 514948
rect 393988 514892 401548 514948
rect 401604 514892 401614 514948
rect 268818 514444 268828 514500
rect 268884 514444 526652 514500
rect 526708 514444 526718 514500
rect 185602 514332 185612 514388
rect 185668 514332 453628 514388
rect 453684 514332 453694 514388
rect 218418 514220 218428 514276
rect 218484 514220 593628 514276
rect 593684 514220 593694 514276
rect 19282 514108 19292 514164
rect 19348 514108 440188 514164
rect 440244 514108 440254 514164
rect 190642 512764 190652 512820
rect 190708 512764 414988 512820
rect 415044 512764 415054 512820
rect 286066 512652 286076 512708
rect 286132 512652 533372 512708
rect 533428 512652 533438 512708
rect 230290 512540 230300 512596
rect 230356 512540 518252 512596
rect 518308 512540 518318 512596
rect 173842 512428 173852 512484
rect 173908 512428 468972 512484
rect 469028 512428 469038 512484
rect 192322 511084 192332 511140
rect 192388 511084 450940 511140
rect 450996 511084 451006 511140
rect 296370 510972 296380 511028
rect 296436 510972 594524 511028
rect 594580 510972 594590 511028
rect 240258 510860 240268 510916
rect 240324 510860 541772 510916
rect 541828 510860 541838 510916
rect 14242 510748 14252 510804
rect 14308 510748 445788 510804
rect 445844 510748 445854 510804
rect 197362 509516 197372 509572
rect 197428 509516 443548 509572
rect 443604 509516 443614 509572
rect 167122 509404 167132 509460
rect 167188 509404 417452 509460
rect 417508 509404 417518 509460
rect 595560 509348 597000 509544
rect 252578 509292 252588 509348
rect 252644 509292 521612 509348
rect 521668 509292 521678 509348
rect 572852 509320 597000 509348
rect 572852 509292 595672 509320
rect 221778 509180 221788 509236
rect 221844 509180 516572 509236
rect 516628 509180 516638 509236
rect 572852 509124 572908 509292
rect 299058 509068 299068 509124
rect 299124 509068 572908 509124
rect 194002 507836 194012 507892
rect 194068 507836 435484 507892
rect 435540 507836 435550 507892
rect 178882 507724 178892 507780
rect 178948 507724 462028 507780
rect 462084 507724 462094 507780
rect 288978 507612 288988 507668
rect 289044 507612 594412 507668
rect 594468 507612 594478 507668
rect 98242 507500 98252 507556
rect 98308 507500 409948 507556
rect 410004 507500 410014 507556
rect 170482 507388 170492 507444
rect 170548 507388 484428 507444
rect 484484 507388 484494 507444
rect 273858 506156 273868 506212
rect 273924 506156 506492 506212
rect 506548 506156 506558 506212
rect 182242 506044 182252 506100
rect 182308 506044 423388 506100
rect 423444 506044 423454 506100
rect 180562 505932 180572 505988
rect 180628 505932 430332 505988
rect 430388 505932 430398 505988
rect 275762 505820 275772 505876
rect 275828 505820 531692 505876
rect 531748 505820 531758 505876
rect 280914 505708 280924 505764
rect 280980 505708 594300 505764
rect 594356 505708 594366 505764
rect 312610 504588 312620 504644
rect 312676 504588 314972 504644
rect 315028 504588 315038 504644
rect 195682 504476 195692 504532
rect 195748 504476 428540 504532
rect 428596 504476 428606 504532
rect 294578 504364 294588 504420
rect 294644 504364 535052 504420
rect 535108 504364 535118 504420
rect 258514 504252 258524 504308
rect 258580 504252 594076 504308
rect 594132 504252 594142 504308
rect 212146 504140 212156 504196
rect 212212 504140 593404 504196
rect 593460 504140 593470 504196
rect 17602 504028 17612 504084
rect 17668 504028 407932 504084
rect 407988 504028 407998 504084
rect 237906 503916 237916 503972
rect 237972 503916 239372 503972
rect 239428 503916 239438 503972
rect 310034 503916 310044 503972
rect 310100 503916 311612 503972
rect 311668 503916 311678 503972
rect 365362 503916 365372 503972
rect 365428 503916 366716 503972
rect 366772 503916 366782 503972
rect 380482 503916 380492 503972
rect 380548 503916 382172 503972
rect 382228 503916 382238 503972
rect 348674 503692 348684 503748
rect 348740 503692 362908 503748
rect 362964 503692 362974 503748
rect 338370 503580 338380 503636
rect 338436 503580 408268 503636
rect 408324 503580 408334 503636
rect 230178 503468 230188 503524
rect 230244 503468 364140 503524
rect 364196 503468 364206 503524
rect 330642 503356 330652 503412
rect 330708 503356 473788 503412
rect 473844 503356 473854 503412
rect 10098 503244 10108 503300
rect 10164 503244 384748 503300
rect 384804 503244 384814 503300
rect 4162 503132 4172 503188
rect 4228 503132 400204 503188
rect 400260 503132 400270 503188
rect 495506 502908 495516 502964
rect 495572 502908 512428 502964
rect 512484 502908 512494 502964
rect 271394 502796 271404 502852
rect 271460 502796 548492 502852
rect 548548 502796 548558 502852
rect -960 502516 480 502712
rect 492930 502684 492940 502740
rect 492996 502684 514108 502740
rect 514164 502684 514174 502740
rect 474898 502572 474908 502628
rect 474964 502572 500668 502628
rect 500724 502572 500734 502628
rect -960 502488 5852 502516
rect 392 502460 5852 502488
rect 5908 502460 5918 502516
rect 188962 502460 188972 502516
rect 189028 502460 438844 502516
rect 438900 502460 438910 502516
rect 477474 502460 477484 502516
rect 477540 502460 509068 502516
rect 509124 502460 509134 502516
rect 199826 502348 199836 502404
rect 199892 502348 209580 502404
rect 209636 502348 209646 502404
rect 490354 502348 490364 502404
rect 490420 502348 504028 502404
rect 504084 502348 504094 502404
rect 5842 501452 5852 501508
rect 5908 501452 405356 501508
rect 405412 501452 405422 501508
rect 302306 501116 302316 501172
rect 302372 501116 499100 501172
rect 499156 501116 499166 501172
rect 199042 501004 199052 501060
rect 199108 501004 420812 501060
rect 420868 501004 420878 501060
rect 482626 501004 482636 501060
rect 482692 501004 502348 501060
rect 502404 501004 502414 501060
rect 292002 500892 292012 500948
rect 292068 500892 514892 500948
rect 514948 500892 514958 500948
rect 263666 500780 263676 500836
rect 263732 500780 545132 500836
rect 545188 500780 545198 500836
rect 191426 500668 191436 500724
rect 191492 500668 217308 500724
rect 217364 500668 217374 500724
rect 227602 500668 227612 500724
rect 227668 500668 593740 500724
rect 593796 500668 593806 500724
rect 408212 499324 420028 499380
rect 467170 499324 467180 499380
rect 467236 499324 467274 499380
rect 408212 499268 408268 499324
rect 419972 499268 420028 499324
rect 266242 499212 266252 499268
rect 266308 499212 267148 499268
rect 284274 499212 284284 499268
rect 284340 499212 408268 499268
rect 413074 499212 413084 499268
rect 413140 499212 413150 499268
rect 419972 499212 513212 499268
rect 513268 499212 513278 499268
rect 267092 499156 267148 499212
rect 267092 499100 412860 499156
rect 412916 499100 412926 499156
rect 413084 499044 413140 499212
rect 413298 499100 413308 499156
rect 413364 499100 594188 499156
rect 594244 499100 594254 499156
rect 15922 498988 15932 499044
rect 15988 498988 413140 499044
rect 467170 498988 467180 499044
rect 467236 498988 498988 499044
rect 499044 498988 499054 499044
rect 595560 496132 597000 496328
rect 595420 496104 597000 496132
rect 595420 496076 595672 496104
rect 595420 496020 595476 496076
rect 595420 495964 595700 496020
rect 595644 495684 595700 495964
rect 499090 495628 499100 495684
rect 499156 495628 595700 495684
rect -960 488404 480 488600
rect -960 488376 532 488404
rect 392 488348 532 488376
rect 476 488292 532 488348
rect 364 488236 532 488292
rect 364 487284 420 488236
rect 364 487228 98252 487284
rect 98308 487228 98318 487284
rect 594514 483084 594524 483140
rect 594580 483112 595672 483140
rect 594580 483084 597000 483112
rect 595560 482888 597000 483084
rect -960 474292 480 474488
rect -960 474264 532 474292
rect 392 474236 532 474264
rect 476 474180 532 474236
rect 364 474124 532 474180
rect 364 473844 420 474124
rect 364 473788 17612 473844
rect 17668 473788 17678 473844
rect 595560 469700 597000 469896
rect 595420 469672 597000 469700
rect 595420 469644 595672 469672
rect 595420 469588 595476 469644
rect 595420 469532 595700 469588
rect 595644 468804 595700 469532
rect 514882 468748 514892 468804
rect 514948 468748 595700 468804
rect -960 460180 480 460376
rect -960 460152 532 460180
rect 392 460124 532 460152
rect 476 460068 532 460124
rect 364 460012 532 460068
rect 364 458724 420 460012
rect 364 458668 15932 458724
rect 15988 458668 15998 458724
rect 595560 456484 597000 456680
rect 595420 456456 597000 456484
rect 595420 456428 595672 456456
rect 595420 456372 595476 456428
rect 595420 456316 595700 456372
rect 595644 455364 595700 456316
rect 535042 455308 535052 455364
rect 535108 455308 595700 455364
rect -960 446068 480 446264
rect -960 446040 532 446068
rect 392 446012 532 446040
rect 476 445956 532 446012
rect 364 445900 532 445956
rect 364 445284 420 445900
rect 364 445228 167132 445284
rect 167188 445228 167198 445284
rect 594402 443436 594412 443492
rect 594468 443464 595672 443492
rect 594468 443436 597000 443464
rect 595560 443240 597000 443436
rect -960 431956 480 432152
rect -960 431928 8428 431956
rect 392 431900 8428 431928
rect 8372 431844 8428 431900
rect 8372 431788 190652 431844
rect 190708 431788 190718 431844
rect 595560 430164 597000 430248
rect 513202 430108 513212 430164
rect 513268 430108 597000 430164
rect 595560 430024 597000 430108
rect -960 417844 480 418040
rect -960 417816 532 417844
rect 392 417788 532 417816
rect 476 417732 532 417788
rect 364 417676 532 417732
rect 364 416724 420 417676
rect 595560 416836 597000 417032
rect 572852 416808 597000 416836
rect 572852 416780 595672 416808
rect 572852 416724 572908 416780
rect 364 416668 199052 416724
rect 199108 416668 199118 416724
rect 533362 416668 533372 416724
rect 533428 416668 572908 416724
rect -960 403732 480 403928
rect 594290 403788 594300 403844
rect 594356 403816 595672 403844
rect 594356 403788 597000 403816
rect -960 403704 532 403732
rect 392 403676 532 403704
rect 476 403620 532 403676
rect 364 403564 532 403620
rect 595560 403592 597000 403788
rect 364 403284 420 403564
rect 364 403228 163772 403284
rect 163828 403228 163838 403284
rect 595560 390404 597000 390600
rect 595420 390376 597000 390404
rect 595420 390348 595672 390376
rect 595420 390292 595476 390348
rect 595420 390236 595700 390292
rect 595644 389844 595700 390236
rect -960 389620 480 389816
rect 531682 389788 531692 389844
rect 531748 389788 595700 389844
rect -960 389592 532 389620
rect 392 389564 532 389592
rect 476 389508 532 389564
rect 364 389452 532 389508
rect 364 388164 420 389452
rect 364 388108 182252 388164
rect 182308 388108 182318 388164
rect 595560 377188 597000 377384
rect 595420 377160 597000 377188
rect 595420 377132 595672 377160
rect 595420 377076 595476 377132
rect 595420 377020 595700 377076
rect 595644 376404 595700 377020
rect 550162 376348 550172 376404
rect 550228 376348 595700 376404
rect -960 375508 480 375704
rect -960 375480 532 375508
rect 392 375452 532 375480
rect 476 375396 532 375452
rect 364 375340 532 375396
rect 364 374724 420 375340
rect 364 374668 195692 374724
rect 195748 374668 195758 374724
rect 595560 363972 597000 364168
rect 595420 363944 597000 363972
rect 595420 363916 595672 363944
rect 595420 363860 595476 363916
rect 595420 363804 595700 363860
rect 595644 362964 595700 363804
rect 506482 362908 506492 362964
rect 506548 362908 595700 362964
rect -960 361396 480 361592
rect -960 361368 8428 361396
rect 392 361340 8428 361368
rect 8372 361284 8428 361340
rect 8372 361228 22652 361284
rect 22708 361228 22718 361284
rect 595560 350756 597000 350952
rect 595420 350728 597000 350756
rect 595420 350700 595672 350728
rect 595420 350644 595476 350700
rect 595420 350588 595700 350644
rect 595644 349524 595700 350588
rect 526642 349468 526652 349524
rect 526708 349468 595700 349524
rect -960 347284 480 347480
rect -960 347256 532 347284
rect 392 347228 532 347256
rect 476 347172 532 347228
rect 364 347116 532 347172
rect 364 346164 420 347116
rect 364 346108 180572 346164
rect 180628 346108 180638 346164
rect 595560 337540 597000 337736
rect 595420 337512 597000 337540
rect 595420 337484 595672 337512
rect 595420 337428 595476 337484
rect 595420 337372 595700 337428
rect 595644 336084 595700 337372
rect 548482 336028 548492 336084
rect 548548 336028 595700 336084
rect -960 333172 480 333368
rect -960 333144 532 333172
rect 392 333116 532 333144
rect 476 333060 532 333116
rect 364 333004 532 333060
rect 364 332724 420 333004
rect 364 332668 194012 332724
rect 194068 332668 194078 332724
rect 594178 324492 594188 324548
rect 594244 324520 595672 324548
rect 594244 324492 597000 324520
rect 595560 324296 597000 324492
rect -960 319060 480 319256
rect -960 319032 532 319060
rect 392 319004 532 319032
rect 476 318948 532 319004
rect 364 318892 532 318948
rect 364 317604 420 318892
rect 364 317548 19292 317604
rect 19348 317548 19358 317604
rect 595560 311108 597000 311304
rect 572852 311080 597000 311108
rect 572852 311052 595672 311080
rect 572852 310884 572908 311052
rect 523282 310828 523292 310884
rect 523348 310828 572908 310884
rect -960 304948 480 305144
rect -960 304920 532 304948
rect 392 304892 532 304920
rect 476 304836 532 304892
rect 364 304780 532 304836
rect 364 304164 420 304780
rect 364 304108 188972 304164
rect 189028 304108 189038 304164
rect 595560 297892 597000 298088
rect 595420 297864 597000 297892
rect 595420 297836 595672 297864
rect 595420 297780 595476 297836
rect 595420 297724 595700 297780
rect 595644 297444 595700 297724
rect 545122 297388 545132 297444
rect 545188 297388 595700 297444
rect -960 290836 480 291032
rect -960 290808 8428 290836
rect 392 290780 8428 290808
rect 8372 290724 8428 290780
rect 8372 290668 197372 290724
rect 197428 290668 197438 290724
rect 594066 284844 594076 284900
rect 594132 284872 595672 284900
rect 594132 284844 597000 284872
rect 595560 284648 597000 284844
rect -960 276724 480 276920
rect -960 276696 532 276724
rect 392 276668 532 276696
rect 476 276612 532 276668
rect 364 276556 532 276612
rect 364 275604 420 276556
rect 364 275548 12572 275604
rect 12628 275548 12638 275604
rect 595560 271460 597000 271656
rect 595420 271432 597000 271460
rect 595420 271404 595672 271432
rect 595420 271348 595476 271404
rect 595420 271292 595700 271348
rect 595644 270564 595700 271292
rect 521602 270508 521612 270564
rect 521668 270508 595700 270564
rect -960 262612 480 262808
rect -960 262584 532 262612
rect 392 262556 532 262584
rect 476 262500 532 262556
rect 364 262444 532 262500
rect 364 262164 420 262444
rect 364 262108 14252 262164
rect 14308 262108 14318 262164
rect 588802 258412 588812 258468
rect 588868 258440 595672 258468
rect 588868 258412 597000 258440
rect 595560 258216 597000 258412
rect -960 248500 480 248696
rect -960 248472 532 248500
rect 392 248444 532 248472
rect 476 248388 532 248444
rect 364 248332 532 248388
rect 364 247044 420 248332
rect 364 246988 192332 247044
rect 192388 246988 192398 247044
rect 593954 245196 593964 245252
rect 594020 245224 595672 245252
rect 594020 245196 597000 245224
rect 595560 245000 597000 245196
rect -960 234388 480 234584
rect -960 234360 532 234388
rect 392 234332 532 234360
rect 476 234276 532 234332
rect 364 234220 532 234276
rect 364 233604 420 234220
rect 364 233548 44492 233604
rect 44548 233548 44558 233604
rect 595560 231924 597000 232008
rect 519922 231868 519932 231924
rect 519988 231868 597000 231924
rect 595560 231784 597000 231868
rect -960 220276 480 220472
rect -960 220248 8428 220276
rect 392 220220 8428 220248
rect 8372 220164 8428 220220
rect 8372 220108 185612 220164
rect 185668 220108 185678 220164
rect 595560 218596 597000 218792
rect 572852 218568 597000 218596
rect 572852 218540 595672 218568
rect 572852 218484 572908 218540
rect 536722 218428 536732 218484
rect 536788 218428 572908 218484
rect 392 206360 9212 206388
rect -960 206332 9212 206360
rect 9268 206332 9278 206388
rect -960 206136 480 206332
rect 593058 205548 593068 205604
rect 593124 205576 595672 205604
rect 593124 205548 597000 205576
rect 595560 205352 597000 205548
rect 144498 199164 144508 199220
rect 144564 199164 278236 199220
rect 278292 199164 278302 199220
rect 474450 199164 474460 199220
rect 474516 199164 560252 199220
rect 560308 199164 560318 199220
rect 65538 199052 65548 199108
rect 65604 199052 241500 199108
rect 241556 199052 241566 199108
rect 475346 199052 475356 199108
rect 475412 199052 593068 199108
rect 593124 199052 593134 199108
rect 179778 198268 179788 198324
rect 179844 198268 294588 198324
rect 294644 198268 294654 198324
rect 212818 198156 212828 198212
rect 212884 198156 215516 198212
rect 215572 198156 215582 198212
rect 234322 198156 234332 198212
rect 234388 198156 237916 198212
rect 237972 198156 237982 198212
rect 292338 198156 292348 198212
rect 292404 198156 294364 198212
rect 294420 198156 294430 198212
rect 314962 198156 314972 198212
rect 315028 198156 323932 198212
rect 323988 198156 323998 198212
rect 341842 198156 341852 198212
rect 341908 198156 342748 198212
rect 342804 198156 342814 198212
rect 343746 198156 343756 198212
rect 343812 198156 344540 198212
rect 344596 198156 344606 198212
rect 355282 198156 355292 198212
rect 355348 198156 356188 198212
rect 356244 198156 356254 198212
rect 367826 198156 367836 198212
rect 367892 198156 371420 198212
rect 371476 198156 371486 198212
rect 373762 198156 373772 198212
rect 373828 198156 375900 198212
rect 375956 198156 375966 198212
rect 378802 198156 378812 198212
rect 378868 198156 379708 198212
rect 379764 198156 379774 198212
rect 390562 198156 390572 198212
rect 390628 198156 392028 198212
rect 392084 198156 392094 198212
rect 392242 198156 392252 198212
rect 392308 198156 393820 198212
rect 393876 198156 393886 198212
rect 399186 198156 399196 198212
rect 399252 198156 400652 198212
rect 400708 198156 400718 198212
rect 400978 198156 400988 198212
rect 401044 198156 404012 198212
rect 404068 198156 404078 198212
rect 435922 198156 435932 198212
rect 435988 198156 438396 198212
rect 438452 198156 438462 198212
rect 471762 198156 471772 198212
rect 471828 198156 472892 198212
rect 472948 198156 472958 198212
rect 478930 198156 478940 198212
rect 478996 198156 488012 198212
rect 488068 198156 488078 198212
rect 340162 198044 340172 198100
rect 340228 198044 349020 198100
rect 349076 198044 349086 198100
rect 375442 198044 375452 198100
rect 375508 198044 382172 198100
rect 382228 198044 382238 198100
rect 411730 198044 411740 198100
rect 411796 198044 414092 198100
rect 414148 198044 414158 198100
rect 422482 198044 422492 198100
rect 422548 198044 430892 198100
rect 430948 198044 430958 198100
rect 438610 198044 438620 198100
rect 438676 198044 454412 198100
rect 454468 198044 454478 198100
rect 197362 197932 197372 197988
rect 197428 197932 224476 197988
rect 224532 197932 224542 197988
rect 300850 197932 300860 197988
rect 300916 197932 310492 197988
rect 310548 197932 310558 197988
rect 351922 197932 351932 197988
rect 351988 197932 354620 197988
rect 354676 197932 354686 197988
rect 447570 197932 447580 197988
rect 447636 197932 486332 197988
rect 486388 197932 486398 197988
rect 182242 197820 182252 197876
rect 182308 197820 196588 197876
rect 308242 197820 308252 197876
rect 308308 197820 345436 197876
rect 345492 197820 345502 197876
rect 424274 197820 424284 197876
rect 424340 197820 444332 197876
rect 444388 197820 444398 197876
rect 450258 197820 450268 197876
rect 450324 197820 494732 197876
rect 494788 197820 494798 197876
rect 196532 197764 196588 197820
rect 196532 197708 221788 197764
rect 221844 197708 221854 197764
rect 223682 197708 223692 197764
rect 223748 197708 313180 197764
rect 313236 197708 313246 197764
rect 323362 197708 323372 197764
rect 323428 197708 331100 197764
rect 331156 197708 331166 197764
rect 336802 197708 336812 197764
rect 336868 197708 352604 197764
rect 352660 197708 352670 197764
rect 365362 197708 365372 197764
rect 365428 197708 370524 197764
rect 370580 197708 370590 197764
rect 437490 197708 437500 197764
rect 437556 197708 483868 197764
rect 483924 197708 483934 197764
rect 209906 197596 209916 197652
rect 209972 197596 311388 197652
rect 311444 197596 311454 197652
rect 328402 197596 328412 197652
rect 328468 197596 364252 197652
rect 364308 197596 364318 197652
rect 416210 197596 416220 197652
rect 416276 197596 436828 197652
rect 436884 197596 436894 197652
rect 446674 197596 446684 197652
rect 446740 197596 467852 197652
rect 467908 197596 467918 197652
rect 482514 197596 482524 197652
rect 482580 197596 531692 197652
rect 531748 197596 531758 197652
rect 113362 197484 113372 197540
rect 113428 197484 219100 197540
rect 219156 197484 219166 197540
rect 224242 197484 224252 197540
rect 224308 197484 240604 197540
rect 240660 197484 240670 197540
rect 241938 197484 241948 197540
rect 242004 197484 309596 197540
rect 309652 197484 309662 197540
rect 311602 197484 311612 197540
rect 311668 197484 346332 197540
rect 346388 197484 346398 197540
rect 420690 197484 420700 197540
rect 420756 197484 446012 197540
rect 446068 197484 446078 197540
rect 452946 197484 452956 197540
rect 453012 197484 506492 197540
rect 506548 197484 506558 197540
rect 94882 197372 94892 197428
rect 94948 197372 254044 197428
rect 254100 197372 254110 197428
rect 254482 197372 254492 197428
rect 254548 197372 260316 197428
rect 260372 197372 260382 197428
rect 264562 197372 264572 197428
rect 264628 197372 273756 197428
rect 273812 197372 273822 197428
rect 274642 197372 274652 197428
rect 274708 197372 337372 197428
rect 337428 197372 337438 197428
rect 340050 197372 340060 197428
rect 340116 197372 354508 197428
rect 354564 197372 354574 197428
rect 359538 197372 359548 197428
rect 359604 197372 379484 197428
rect 379540 197372 379550 197428
rect 398290 197372 398300 197428
rect 398356 197372 399868 197428
rect 399924 197372 399934 197428
rect 405458 197372 405468 197428
rect 405524 197372 412412 197428
rect 412468 197372 412478 197428
rect 431442 197372 431452 197428
rect 431508 197372 478940 197428
rect 478996 197372 479006 197428
rect 484306 197372 484316 197428
rect 484372 197372 570332 197428
rect 570388 197372 570398 197428
rect 214946 197260 214956 197316
rect 215012 197260 223692 197316
rect 223748 197260 223758 197316
rect 370402 197260 370412 197316
rect 370468 197260 372316 197316
rect 372372 197260 372382 197316
rect 400082 197260 400092 197316
rect 400148 197260 402332 197316
rect 402388 197260 402398 197316
rect 257058 197148 257068 197204
rect 257124 197148 259420 197204
rect 259476 197148 259486 197204
rect 343522 197036 343532 197092
rect 343588 197036 348124 197092
rect 348180 197036 348190 197092
rect 356962 197036 356972 197092
rect 357028 197036 358876 197092
rect 358932 197036 358942 197092
rect 404562 197036 404572 197092
rect 404628 197036 405692 197092
rect 405748 197036 405758 197092
rect 470866 197036 470876 197092
rect 470932 197036 479052 197092
rect 479108 197036 479118 197092
rect 413522 196924 413532 196980
rect 413588 196924 415772 196980
rect 415828 196924 415838 196980
rect 454738 196924 454748 196980
rect 454804 196924 456092 196980
rect 456148 196924 456158 196980
rect 283042 196700 283052 196756
rect 283108 196700 290780 196756
rect 290836 196700 290846 196756
rect 380482 196700 380492 196756
rect 380548 196700 386652 196756
rect 386708 196700 386718 196756
rect 412626 196700 412636 196756
rect 412692 196700 422492 196756
rect 422548 196700 422558 196756
rect 253698 196588 253708 196644
rect 253764 196588 256732 196644
rect 256788 196588 256798 196644
rect 288082 196588 288092 196644
rect 288148 196588 291676 196644
rect 291732 196588 291742 196644
rect 324370 196588 324380 196644
rect 324436 196588 326620 196644
rect 326676 196588 326686 196644
rect 383842 196588 383852 196644
rect 383908 196588 385756 196644
rect 385812 196588 385822 196644
rect 394818 196588 394828 196644
rect 394884 196588 396508 196644
rect 396564 196588 396574 196644
rect 418002 196588 418012 196644
rect 418068 196588 422716 196644
rect 422772 196588 422782 196644
rect 211698 196028 211708 196084
rect 211764 196028 300860 196084
rect 300916 196028 300926 196084
rect 132626 195916 132636 195972
rect 132692 195916 272860 195972
rect 272916 195916 272926 195972
rect 357858 195916 357868 195972
rect 357924 195916 378588 195972
rect 378644 195916 378654 195972
rect 452050 195916 452060 195972
rect 452116 195916 519148 195972
rect 519204 195916 519214 195972
rect 57026 195804 57036 195860
rect 57092 195804 237020 195860
rect 237076 195804 237086 195860
rect 346098 195804 346108 195860
rect 346164 195804 373212 195860
rect 373268 195804 373278 195860
rect 421698 195804 421708 195860
rect 421764 195804 448588 195860
rect 448644 195804 448654 195860
rect 469074 195804 469084 195860
rect 469140 195804 549388 195860
rect 549444 195804 549454 195860
rect 10098 195692 10108 195748
rect 10164 195692 212828 195748
rect 212884 195692 212894 195748
rect 220098 195692 220108 195748
rect 220164 195692 314076 195748
rect 314132 195692 314142 195748
rect 329522 195692 329532 195748
rect 329588 195692 365148 195748
rect 365204 195692 365214 195748
rect 378018 195692 378028 195748
rect 378084 195692 388444 195748
rect 388500 195692 388510 195748
rect 440178 195692 440188 195748
rect 440244 195692 487228 195748
rect 487284 195692 487294 195748
rect 488002 195692 488012 195748
rect 488068 195692 571228 195748
rect 571284 195692 571294 195748
rect 210018 194348 210028 194404
rect 210084 194348 241948 194404
rect 242004 194348 242014 194404
rect 137778 194236 137788 194292
rect 137844 194236 275436 194292
rect 275492 194236 275502 194292
rect 104178 194124 104188 194180
rect 104244 194124 257068 194180
rect 257124 194124 257134 194180
rect 458322 194124 458332 194180
rect 458388 194124 525868 194180
rect 525924 194124 525934 194180
rect 29362 194012 29372 194068
rect 29428 194012 222684 194068
rect 222740 194012 222750 194068
rect 261202 194012 261212 194068
rect 261268 194012 331996 194068
rect 332052 194012 332062 194068
rect 472658 194012 472668 194068
rect 472724 194012 557788 194068
rect 557844 194012 557854 194068
rect 194002 192556 194012 192612
rect 194068 192556 299740 192612
rect 299796 192556 299806 192612
rect 443986 192556 443996 192612
rect 444052 192556 495628 192612
rect 495684 192556 495694 192612
rect 97458 192444 97468 192500
rect 97524 192444 253708 192500
rect 253764 192444 253774 192500
rect 455634 192444 455644 192500
rect 455700 192444 520828 192500
rect 520884 192444 520894 192500
rect 22642 192332 22652 192388
rect 22708 192332 217308 192388
rect 217364 192332 217374 192388
rect 246978 192332 246988 192388
rect 247044 192332 324380 192388
rect 324436 192332 324446 192388
rect 477138 192332 477148 192388
rect 477204 192332 572908 192388
rect 590482 192332 590492 192388
rect 590548 192360 595672 192388
rect 590548 192332 597000 192360
rect 572852 192276 572908 192332
rect -960 192052 480 192248
rect 572852 192220 593964 192276
rect 594020 192220 594030 192276
rect 595560 192136 597000 192332
rect -960 192024 532 192052
rect 392 191996 532 192024
rect 476 191940 532 191996
rect 364 191884 532 191940
rect 364 191604 420 191884
rect 364 191548 27692 191604
rect 27748 191548 27758 191604
rect 206658 190876 206668 190932
rect 206724 190876 307804 190932
rect 307860 190876 307870 190932
rect 154466 190764 154476 190820
rect 154532 190764 283612 190820
rect 283668 190764 283678 190820
rect 456530 190764 456540 190820
rect 456596 190764 522508 190820
rect 522564 190764 522574 190820
rect 27682 190652 27692 190708
rect 27748 190652 220892 190708
rect 220948 190652 220958 190708
rect 479826 190652 479836 190708
rect 479892 190652 572908 190708
rect 572964 190652 572974 190708
rect 178098 189196 178108 189252
rect 178164 189196 292348 189252
rect 292404 189196 292414 189252
rect 36978 189084 36988 189140
rect 37044 189084 228060 189140
rect 228116 189084 228126 189140
rect 479042 189084 479052 189140
rect 479108 189084 552748 189140
rect 552804 189084 552814 189140
rect 31938 188972 31948 189028
rect 32004 188972 225372 189028
rect 225428 188972 225438 189028
rect 252018 188972 252028 189028
rect 252084 188972 329308 189028
rect 329364 188972 329374 189028
rect 438386 188972 438396 189028
rect 438452 188972 478828 189028
rect 478884 188972 478894 189028
rect 480722 188972 480732 189028
rect 480788 188972 574588 189028
rect 574644 188972 574654 189028
rect 201618 187516 201628 187572
rect 201684 187516 305116 187572
rect 305172 187516 305182 187572
rect 134418 187404 134428 187460
rect 134484 187404 264572 187460
rect 264628 187404 264638 187460
rect 442194 187404 442204 187460
rect 442260 187404 491372 187460
rect 491428 187404 491438 187460
rect 45378 187292 45388 187348
rect 45444 187292 231644 187348
rect 231700 187292 231710 187348
rect 466386 187292 466396 187348
rect 466452 187292 544348 187348
rect 544404 187292 544414 187348
rect 203298 185836 203308 185892
rect 203364 185836 306012 185892
rect 306068 185836 306078 185892
rect 99922 185724 99932 185780
rect 99988 185724 255836 185780
rect 255892 185724 255902 185780
rect 80658 185612 80668 185668
rect 80724 185612 248668 185668
rect 248724 185612 248734 185668
rect 461010 185612 461020 185668
rect 461076 185612 532588 185668
rect 532644 185612 532654 185668
rect 248658 184156 248668 184212
rect 248724 184156 327516 184212
rect 327572 184156 327582 184212
rect 105858 184044 105868 184100
rect 105924 184044 254492 184100
rect 254548 184044 254558 184100
rect 89058 183932 89068 183988
rect 89124 183932 252252 183988
rect 252308 183932 252318 183988
rect 463698 183932 463708 183988
rect 463764 183932 536732 183988
rect 536788 183932 536798 183988
rect 139458 182476 139468 182532
rect 139524 182476 276444 182532
rect 276500 182476 276510 182532
rect 117618 182364 117628 182420
rect 117684 182364 265692 182420
rect 265748 182364 265758 182420
rect 72258 182252 72268 182308
rect 72324 182252 244188 182308
rect 244244 182252 244254 182308
rect 472882 182252 472892 182308
rect 472948 182252 554428 182308
rect 554484 182252 554494 182308
rect 285618 180908 285628 180964
rect 285684 180908 343756 180964
rect 343812 180908 343822 180964
rect 162978 180684 162988 180740
rect 163044 180684 287196 180740
rect 287252 180684 287262 180740
rect 47058 180572 47068 180628
rect 47124 180572 232540 180628
rect 232596 180572 232606 180628
rect 467282 180572 467292 180628
rect 467348 180572 541884 180628
rect 541940 180572 541950 180628
rect 194898 179116 194908 179172
rect 194964 179116 302428 179172
rect 302484 179116 302494 179172
rect 142818 179004 142828 179060
rect 142884 179004 277340 179060
rect 277396 179004 277406 179060
rect 595560 178948 597000 179144
rect 41122 178892 41132 178948
rect 41188 178892 228956 178948
rect 229012 178892 229022 178948
rect 457426 178892 457436 178948
rect 457492 178892 518364 178948
rect 518420 178892 518430 178948
rect 595420 178920 597000 178948
rect 595420 178892 595672 178920
rect 595420 178836 595476 178892
rect 595420 178780 595700 178836
rect 595644 178164 595700 178780
rect -960 177940 480 178136
rect 541762 178108 541772 178164
rect 541828 178108 595700 178164
rect -960 177912 532 177940
rect 392 177884 532 177912
rect 476 177828 532 177884
rect 364 177772 532 177828
rect 364 176484 420 177772
rect 174738 177324 174748 177380
rect 174804 177324 292572 177380
rect 292628 177324 292638 177380
rect 136098 177212 136108 177268
rect 136164 177212 273868 177268
rect 273924 177212 273934 177268
rect 460114 177212 460124 177268
rect 460180 177212 534268 177268
rect 534324 177212 534334 177268
rect 364 176428 178892 176484
rect 178948 176428 178958 176484
rect 185602 175644 185612 175700
rect 185668 175644 297052 175700
rect 297108 175644 297118 175700
rect 87378 175532 87388 175588
rect 87444 175532 251356 175588
rect 251412 175532 251422 175588
rect 142706 173964 142716 174020
rect 142772 173964 279132 174020
rect 279188 173964 279198 174020
rect 109218 173852 109228 173908
rect 109284 173852 262108 173908
rect 262164 173852 262174 173908
rect 188962 172284 188972 172340
rect 189028 172284 297948 172340
rect 298004 172284 298014 172340
rect 115938 172172 115948 172228
rect 116004 172172 264796 172228
rect 264852 172172 264862 172228
rect 120978 170492 120988 170548
rect 121044 170492 267484 170548
rect 267540 170492 267550 170548
rect 126018 168812 126028 168868
rect 126084 168812 270172 168868
rect 270228 168812 270238 168868
rect 149426 167244 149436 167300
rect 149492 167244 280924 167300
rect 280980 167244 280990 167300
rect 71362 167132 71372 167188
rect 71428 167132 242396 167188
rect 242452 167132 242462 167188
rect 593842 165900 593852 165956
rect 593908 165928 595672 165956
rect 593908 165900 597000 165928
rect 595560 165704 597000 165900
rect 161298 165564 161308 165620
rect 161364 165564 286300 165620
rect 286356 165564 286366 165620
rect 62962 165452 62972 165508
rect 63028 165452 238812 165508
rect 238868 165452 238878 165508
rect 445778 165452 445788 165508
rect 445844 165452 499772 165508
rect 499828 165452 499838 165508
rect -960 163828 480 164024
rect -960 163800 532 163828
rect 392 163772 532 163800
rect 476 163716 532 163772
rect 364 163660 532 163716
rect 364 163044 420 163660
rect 364 162988 498988 163044
rect 499044 162988 499054 163044
rect 166338 162092 166348 162148
rect 166404 162092 288988 162148
rect 289044 162092 289054 162148
rect 52098 160412 52108 160468
rect 52164 160412 235228 160468
rect 235284 160412 235294 160468
rect 58818 158732 58828 158788
rect 58884 158732 234332 158788
rect 234388 158732 234398 158788
rect 63858 157052 63868 157108
rect 63924 157052 224252 157108
rect 224308 157052 224318 157108
rect 75618 155372 75628 155428
rect 75684 155372 245980 155428
rect 246036 155372 246046 155428
rect 100818 153692 100828 153748
rect 100884 153692 257628 153748
rect 257684 153692 257694 153748
rect 595560 152516 597000 152712
rect 595420 152488 597000 152516
rect 595420 152460 595672 152488
rect 595420 152404 595476 152460
rect 595420 152348 595700 152404
rect 129266 152012 129276 152068
rect 129332 152012 271068 152068
rect 271124 152012 271134 152068
rect 595644 151284 595700 152348
rect 518242 151228 518252 151284
rect 518308 151228 595700 151284
rect 157938 150332 157948 150388
rect 158004 150332 284508 150388
rect 284564 150332 284574 150388
rect -960 149716 480 149912
rect -960 149688 8428 149716
rect 392 149660 8428 149688
rect 8372 149604 8428 149660
rect 8372 149548 158732 149604
rect 158788 149548 158798 149604
rect 107538 148652 107548 148708
rect 107604 148652 260428 148708
rect 260484 148652 260494 148708
rect 84802 146972 84812 147028
rect 84868 146972 247772 147028
rect 247828 146972 247838 147028
rect 595560 139300 597000 139496
rect 595420 139272 597000 139300
rect 595420 139244 595672 139272
rect 595420 139188 595476 139244
rect 595420 139132 595700 139188
rect 595644 137844 595700 139132
rect 540082 137788 540092 137844
rect 540148 137788 595700 137844
rect -960 135604 480 135800
rect -960 135576 532 135604
rect 392 135548 532 135576
rect 476 135492 532 135548
rect 364 135436 532 135492
rect 364 134484 420 135436
rect 173058 135212 173068 135268
rect 173124 135212 288092 135268
rect 288148 135212 288158 135268
rect 444882 135212 444892 135268
rect 444948 135212 497308 135268
rect 497364 135212 497374 135268
rect 364 134428 173852 134484
rect 173908 134428 173918 134484
rect 593730 126252 593740 126308
rect 593796 126280 595672 126308
rect 593796 126252 597000 126280
rect 595560 126056 597000 126252
rect 449362 123452 449372 123508
rect 449428 123452 501452 123508
rect 501508 123452 501518 123508
rect -960 121492 480 121688
rect -960 121464 532 121492
rect 392 121436 532 121464
rect 476 121380 532 121436
rect 364 121324 532 121380
rect 364 121044 420 121324
rect 364 120988 500668 121044
rect 500724 120988 500734 121044
rect 437714 120092 437724 120148
rect 437780 120092 482188 120148
rect 482244 120092 482254 120148
rect 595560 112868 597000 113064
rect 572852 112840 597000 112868
rect 572852 112812 595672 112840
rect 572852 112644 572908 112812
rect 516562 112588 516572 112644
rect 516628 112588 572908 112644
rect -960 107380 480 107576
rect -960 107352 532 107380
rect 392 107324 532 107352
rect 476 107268 532 107324
rect 364 107212 532 107268
rect 364 105924 420 107212
rect 364 105868 157052 105924
rect 157108 105868 157118 105924
rect 595560 99652 597000 99848
rect 595420 99624 597000 99652
rect 595420 99596 595672 99624
rect 595420 99540 595476 99596
rect 595420 99484 595700 99540
rect 595644 99204 595700 99484
rect 538402 99148 538412 99204
rect 538468 99148 595700 99204
rect 4162 94892 4172 94948
rect 4228 94892 509068 94948
rect 509124 94892 509134 94948
rect 392 93464 4172 93492
rect -960 93436 4172 93464
rect 4228 93436 4238 93492
rect -960 93240 480 93436
rect 171378 93212 171388 93268
rect 171444 93212 283052 93268
rect 283108 93212 283118 93268
rect 593618 86604 593628 86660
rect 593684 86632 595672 86660
rect 593684 86604 597000 86632
rect 595560 86408 597000 86604
rect -960 79156 480 79352
rect -960 79128 8428 79156
rect 392 79100 8428 79128
rect 8372 79044 8428 79100
rect 8372 78988 502348 79044
rect 502404 78988 502414 79044
rect 593506 73388 593516 73444
rect 593572 73416 595672 73444
rect 593572 73388 597000 73416
rect 595560 73192 597000 73388
rect 78082 66332 78092 66388
rect 78148 66332 245084 66388
rect 245140 66332 245150 66388
rect -960 65044 480 65240
rect -960 65016 532 65044
rect 392 64988 532 65016
rect 476 64932 532 64988
rect 364 64876 532 64932
rect 364 63924 420 64876
rect 364 63868 155372 63924
rect 155428 63868 155438 63924
rect 68002 61292 68012 61348
rect 68068 61292 239708 61348
rect 239764 61292 239774 61348
rect 430546 61292 430556 61348
rect 430612 61292 468860 61348
rect 468916 61292 468926 61348
rect 595560 60004 597000 60200
rect 595420 59976 597000 60004
rect 595420 59948 595672 59976
rect 595420 59892 595476 59948
rect 595420 59836 595700 59892
rect 595644 58884 595700 59836
rect 191426 58828 191436 58884
rect 191492 58828 595700 58884
rect 44482 56252 44492 56308
rect 44548 56252 229852 56308
rect 229908 56252 229918 56308
rect 53778 54572 53788 54628
rect 53844 54572 236124 54628
rect 236180 54572 236190 54628
rect 469970 54572 469980 54628
rect 470036 54572 551068 54628
rect 551124 54572 551134 54628
rect 48738 52892 48748 52948
rect 48804 52892 233436 52948
rect 233492 52892 233502 52948
rect 386530 52108 386540 52164
rect 386596 52108 390572 52164
rect 390628 52108 390638 52164
rect 207442 51212 207452 51268
rect 207508 51212 306908 51268
rect 306964 51212 306974 51268
rect 432338 51212 432348 51268
rect 432404 51212 472108 51268
rect 472164 51212 472174 51268
rect -960 50932 480 51128
rect -960 50904 532 50932
rect 392 50876 532 50904
rect 476 50820 532 50876
rect 364 50764 532 50820
rect 364 50484 420 50764
rect 364 50428 170492 50484
rect 170548 50428 170558 50484
rect 170482 49532 170492 49588
rect 170548 49532 289884 49588
rect 289940 49532 289950 49588
rect 191538 47852 191548 47908
rect 191604 47852 300636 47908
rect 300692 47852 300702 47908
rect 593394 46956 593404 47012
rect 593460 46984 595672 47012
rect 593460 46956 597000 46984
rect 595560 46760 597000 46956
rect 231858 46172 231868 46228
rect 231924 46172 319452 46228
rect 319508 46172 319518 46228
rect 30258 44492 30268 44548
rect 30324 44492 197372 44548
rect 197428 44492 197438 44548
rect 230290 44492 230300 44548
rect 230356 44492 318556 44548
rect 318612 44492 318622 44548
rect 119298 42924 119308 42980
rect 119364 42924 266588 42980
rect 266644 42924 266654 42980
rect 266242 42812 266252 42868
rect 266308 42812 334684 42868
rect 334740 42812 334750 42868
rect 4162 41132 4172 41188
rect 4228 41132 504028 41188
rect 504084 41132 504094 41188
rect 208338 39452 208348 39508
rect 208404 39452 308700 39508
rect 308756 39452 308766 39508
rect 193218 37884 193228 37940
rect 193284 37884 300748 37940
rect 300804 37884 300814 37940
rect 68898 37772 68908 37828
rect 68964 37772 243292 37828
rect 243348 37772 243358 37828
rect 300962 37772 300972 37828
rect 301028 37772 351708 37828
rect 351764 37772 351774 37828
rect 429650 37772 429660 37828
rect 429716 37772 465388 37828
rect 465444 37772 465454 37828
rect -960 36932 480 37016
rect -960 36876 4172 36932
rect 4228 36876 4238 36932
rect -960 36792 480 36876
rect 196578 36092 196588 36148
rect 196644 36092 303324 36148
rect 303380 36092 303390 36148
rect 305778 36092 305788 36148
rect 305844 36092 354396 36148
rect 354452 36092 354462 36148
rect 486322 36092 486332 36148
rect 486388 36092 504028 36148
rect 504084 36092 504094 36148
rect 199826 34412 199836 34468
rect 199892 34412 590492 34468
rect 590548 34412 590558 34468
rect 593282 33740 593292 33796
rect 593348 33768 595672 33796
rect 593348 33740 597000 33768
rect 595560 33544 597000 33740
rect 90738 32844 90748 32900
rect 90804 32844 253148 32900
rect 253204 32844 253214 32900
rect 274754 32844 274764 32900
rect 274820 32844 338268 32900
rect 338324 32844 338334 32900
rect 252802 32732 252812 32788
rect 252868 32732 327628 32788
rect 327684 32732 327694 32788
rect 339490 32732 339500 32788
rect 339556 32732 365372 32788
rect 365428 32732 365438 32788
rect 506482 32620 506492 32676
rect 506548 32620 515788 32676
rect 515844 32620 515854 32676
rect 199826 31164 199836 31220
rect 199892 31164 304220 31220
rect 304276 31164 304286 31220
rect 11778 31052 11788 31108
rect 11844 31052 216412 31108
rect 216468 31052 216478 31108
rect 243618 31052 243628 31108
rect 243684 31052 324828 31108
rect 324884 31052 324894 31108
rect 351138 31052 351148 31108
rect 351204 31052 373772 31108
rect 373828 31052 373838 31108
rect 302418 29596 302428 29652
rect 302484 29596 336812 29652
rect 336868 29596 336878 29652
rect 225922 29484 225932 29540
rect 225988 29484 315868 29540
rect 315924 29484 315934 29540
rect 151218 29372 151228 29428
rect 151284 29372 281820 29428
rect 281876 29372 281886 29428
rect 334450 29372 334460 29428
rect 334516 29372 371420 29428
rect 371476 29372 371486 29428
rect 468738 29372 468748 29428
rect 468804 29372 478940 29428
rect 478996 29372 479006 29428
rect 483410 29372 483420 29428
rect 483476 29372 581308 29428
rect 581364 29372 581374 29428
rect 4274 27692 4284 27748
rect 4340 27692 512428 27748
rect 512484 27692 512494 27748
rect 4162 26012 4172 26068
rect 4228 26012 514108 26068
rect 514164 26012 514174 26068
rect 531682 26012 531692 26068
rect 531748 26012 579628 26068
rect 579684 26012 579694 26068
rect 209906 25116 209916 25172
rect 209972 25116 215068 25172
rect 215124 25116 215134 25172
rect 233650 24444 233660 24500
rect 233716 24444 320348 24500
rect 320404 24444 320414 24500
rect 113474 24332 113484 24388
rect 113540 24332 263004 24388
rect 263060 24332 263070 24388
rect 297490 24332 297500 24388
rect 297556 24332 350812 24388
rect 350868 24332 350878 24388
rect 441298 24332 441308 24388
rect 441364 24332 490588 24388
rect 490644 24332 490654 24388
rect 392 22904 4284 22932
rect -960 22876 4284 22904
rect 4340 22876 4350 22932
rect -960 22680 480 22876
rect 279010 22764 279020 22820
rect 279076 22764 341068 22820
rect 341124 22764 341134 22820
rect 176418 22652 176428 22708
rect 176484 22652 293468 22708
rect 293524 22652 293534 22708
rect 443090 22652 443100 22708
rect 443156 22652 493948 22708
rect 494004 22652 494014 22708
rect 494722 22652 494732 22708
rect 494788 22652 509068 22708
rect 509124 22652 509134 22708
rect 265458 21196 265468 21252
rect 265524 21196 335580 21252
rect 335636 21196 335646 21252
rect 181458 21084 181468 21140
rect 181524 21084 296156 21140
rect 296212 21084 296222 21140
rect 131058 20972 131068 21028
rect 131124 20972 271964 21028
rect 272020 20972 272030 21028
rect 316642 20972 316652 21028
rect 316708 20972 357980 21028
rect 358036 20972 358046 21028
rect 426962 20972 426972 21028
rect 427028 20972 460348 21028
rect 460404 20972 460414 21028
rect 464594 20972 464604 21028
rect 464660 20972 539308 21028
rect 539364 20972 539374 21028
rect 590482 20524 590492 20580
rect 590548 20552 595672 20580
rect 590548 20524 597000 20552
rect 595560 20328 597000 20524
rect 228498 19404 228508 19460
rect 228564 19404 317548 19460
rect 317604 19404 317614 19460
rect 317874 19404 317884 19460
rect 317940 19404 359772 19460
rect 359828 19404 359838 19460
rect 124338 19292 124348 19348
rect 124404 19292 269276 19348
rect 269332 19292 269342 19348
rect 292338 19292 292348 19348
rect 292404 19292 343532 19348
rect 343588 19292 343598 19348
rect 349570 19292 349580 19348
rect 349636 19292 375004 19348
rect 375060 19292 375070 19348
rect 453842 19292 453852 19348
rect 453908 19292 517468 19348
rect 517524 19292 517534 19348
rect 147858 17724 147868 17780
rect 147924 17724 280028 17780
rect 280084 17724 280094 17780
rect 304098 17724 304108 17780
rect 304164 17724 353500 17780
rect 353556 17724 353566 17780
rect 82338 17612 82348 17668
rect 82404 17612 249564 17668
rect 249620 17612 249630 17668
rect 253810 17612 253820 17668
rect 253876 17612 330204 17668
rect 330260 17612 330270 17668
rect 454402 17612 454412 17668
rect 454468 17612 485548 17668
rect 485604 17612 485614 17668
rect 444322 17500 444332 17556
rect 444388 17500 453628 17556
rect 453684 17500 453694 17556
rect 287410 16156 287420 16212
rect 287476 16156 308252 16212
rect 308308 16156 308318 16212
rect 188402 16044 188412 16100
rect 188468 16044 298844 16100
rect 298900 16044 298910 16100
rect 322690 16044 322700 16100
rect 322756 16044 362460 16100
rect 362516 16044 362526 16100
rect 122658 15932 122668 15988
rect 122724 15932 268380 15988
rect 268436 15932 268446 15988
rect 307458 15932 307468 15988
rect 307524 15932 351932 15988
rect 351988 15932 351998 15988
rect 361666 15932 361676 15988
rect 361732 15932 378812 15988
rect 378868 15932 378878 15988
rect 418898 15932 418908 15988
rect 418964 15932 443548 15988
rect 443604 15932 443614 15988
rect 461906 15932 461916 15988
rect 461972 15932 534380 15988
rect 534436 15932 534446 15988
rect 262098 14588 262108 14644
rect 262164 14588 333788 14644
rect 333844 14588 333854 14644
rect 257170 14476 257180 14532
rect 257236 14476 323372 14532
rect 323428 14476 323438 14532
rect 267138 14364 267148 14420
rect 267204 14364 336476 14420
rect 336532 14364 336542 14420
rect 33618 14252 33628 14308
rect 33684 14252 226268 14308
rect 226324 14252 226334 14308
rect 333106 14252 333116 14308
rect 333172 14252 368060 14308
rect 368116 14252 368126 14308
rect 434130 14252 434140 14308
rect 434196 14252 475468 14308
rect 475524 14252 475534 14308
rect 478034 14252 478044 14308
rect 478100 14252 567868 14308
rect 567924 14252 567934 14308
rect 390226 12908 390236 12964
rect 390292 12908 392252 12964
rect 392308 12908 392318 12964
rect 277218 12796 277228 12852
rect 277284 12796 340956 12852
rect 341012 12796 341022 12852
rect 238578 12684 238588 12740
rect 238644 12684 323036 12740
rect 323092 12684 323102 12740
rect 18498 12572 18508 12628
rect 18564 12572 113372 12628
rect 113428 12572 113438 12628
rect 159842 12572 159852 12628
rect 159908 12572 285404 12628
rect 285460 12572 285470 12628
rect 295698 12572 295708 12628
rect 295764 12572 349916 12628
rect 349972 12572 349982 12628
rect 383282 12572 383292 12628
rect 383348 12572 391132 12628
rect 391188 12572 391198 12628
rect 414418 12572 414428 12628
rect 414484 12572 433468 12628
rect 433524 12572 433534 12628
rect 435026 12572 435036 12628
rect 435092 12572 477148 12628
rect 477204 12572 477214 12628
rect 481618 12572 481628 12628
rect 481684 12572 576268 12628
rect 576324 12572 576334 12628
rect 481842 11564 481852 11620
rect 481908 11564 483868 11620
rect 483924 11564 483934 11620
rect 289538 11228 289548 11284
rect 289604 11228 311612 11284
rect 311668 11228 311678 11284
rect 312386 11116 312396 11172
rect 312452 11116 357084 11172
rect 357140 11116 357150 11172
rect 226706 11004 226716 11060
rect 226772 11004 316764 11060
rect 316820 11004 316830 11060
rect 339042 11004 339052 11060
rect 339108 11004 369628 11060
rect 369684 11004 369694 11060
rect 427858 11004 427868 11060
rect 427924 11004 462588 11060
rect 462644 11004 462654 11060
rect 102946 10892 102956 10948
rect 103012 10892 258524 10948
rect 258580 10892 258590 10948
rect 281922 10892 281932 10948
rect 281988 10892 341852 10948
rect 341908 10892 341918 10948
rect 428754 10892 428764 10948
rect 428820 10892 464492 10948
rect 464548 10892 464558 10948
rect 467842 10892 467852 10948
rect 467908 10892 502572 10948
rect 502628 10892 502638 10948
rect 274306 9436 274316 9492
rect 274372 9436 339164 9492
rect 339220 9436 339230 9492
rect 154354 9324 154364 9380
rect 154420 9324 282716 9380
rect 282772 9324 282782 9380
rect 422706 9324 422716 9380
rect 422772 9324 441644 9380
rect 441700 9324 441710 9380
rect 24882 9212 24892 9268
rect 24948 9212 182252 9268
rect 182308 9212 182318 9268
rect 260978 9212 260988 9268
rect 261044 9212 332892 9268
rect 332948 9212 332958 9268
rect 426066 9212 426076 9268
rect 426132 9212 458780 9268
rect 458836 9212 458846 9268
rect 459218 9212 459228 9268
rect 459284 9212 529228 9268
rect 529284 9212 529294 9268
rect 392 8792 4172 8820
rect -960 8764 4172 8792
rect 4228 8764 4238 8820
rect 375218 8764 375228 8820
rect 375284 8764 380492 8820
rect 380548 8764 380558 8820
rect -960 8568 480 8764
rect 365698 8428 365708 8484
rect 365764 8428 375452 8484
rect 375508 8428 375518 8484
rect 409938 7980 409948 8036
rect 410004 7980 424508 8036
rect 424564 7980 424574 8036
rect 316194 7868 316204 7924
rect 316260 7868 356972 7924
rect 357028 7868 357038 7924
rect 236226 7756 236236 7812
rect 236292 7756 321244 7812
rect 321300 7756 321310 7812
rect 423378 7756 423388 7812
rect 423444 7756 453068 7812
rect 453124 7756 453134 7812
rect 165778 7644 165788 7700
rect 165844 7644 287308 7700
rect 287364 7644 287374 7700
rect 291442 7644 291452 7700
rect 291508 7644 347228 7700
rect 347284 7644 347294 7700
rect 440402 7644 440412 7700
rect 440468 7644 489244 7700
rect 489300 7644 489310 7700
rect 78194 7532 78204 7588
rect 78260 7532 246876 7588
rect 246932 7532 246942 7588
rect 276210 7532 276220 7588
rect 276276 7532 354508 7588
rect 354564 7532 354574 7588
rect 356066 7532 356076 7588
rect 356132 7532 377692 7588
rect 377748 7532 377758 7588
rect 415762 7532 415772 7588
rect 415828 7532 432124 7588
rect 432180 7532 432190 7588
rect 448466 7532 448476 7588
rect 448532 7532 506380 7588
rect 506436 7532 506446 7588
rect 593170 7308 593180 7364
rect 593236 7336 595672 7364
rect 593236 7308 597000 7336
rect 595560 7112 597000 7308
rect 468738 6972 468748 7028
rect 468804 6972 469532 7028
rect 469588 6972 469598 7028
rect 270386 6748 270396 6804
rect 270452 6748 274652 6804
rect 274708 6748 274718 6804
rect 373314 6748 373324 6804
rect 373380 6748 383852 6804
rect 383908 6748 383918 6804
rect 446002 6748 446012 6804
rect 446068 6748 447356 6804
rect 447412 6748 447422 6804
rect 17266 6188 17276 6244
rect 17332 6188 218204 6244
rect 218260 6188 218270 6244
rect 310482 6188 310492 6244
rect 310548 6188 355292 6244
rect 355348 6188 355358 6244
rect 238130 6076 238140 6132
rect 238196 6076 322140 6132
rect 322196 6076 322206 6132
rect 422482 6076 422492 6132
rect 422548 6076 430220 6132
rect 430276 6076 430286 6132
rect 433234 6076 433244 6132
rect 433300 6076 474012 6132
rect 474068 6076 474078 6132
rect 95330 5964 95340 6020
rect 95396 5964 254940 6020
rect 254996 5964 255006 6020
rect 283826 5964 283836 6020
rect 283892 5964 343644 6020
rect 343700 5964 343710 6020
rect 344754 5964 344764 6020
rect 344820 5964 370412 6020
rect 370468 5964 370478 6020
rect 414082 5964 414092 6020
rect 414148 5964 428428 6020
rect 428484 5964 428494 6020
rect 430882 5964 430892 6020
rect 430948 5964 451164 6020
rect 451220 5964 451230 6020
rect 451378 5964 451388 6020
rect 451444 5964 512092 6020
rect 512148 5964 512158 6020
rect 220052 5852 312284 5908
rect 312340 5852 312350 5908
rect 321906 5852 321916 5908
rect 321972 5852 361228 5908
rect 361284 5852 361294 5908
rect 405682 5852 405692 5908
rect 405748 5852 413084 5908
rect 413140 5852 413150 5908
rect 415314 5852 415324 5908
rect 415380 5852 435932 5908
rect 435988 5852 435998 5908
rect 456082 5852 456092 5908
rect 456148 5852 519708 5908
rect 519764 5852 519774 5908
rect 220052 5796 220108 5852
rect 217186 5740 217196 5796
rect 217252 5740 220108 5796
rect 412402 5740 412412 5796
rect 412468 5740 414988 5796
rect 415044 5740 415054 5796
rect 93426 5068 93436 5124
rect 93492 5068 94892 5124
rect 94948 5068 94958 5124
rect 214946 5068 214956 5124
rect 215012 5068 218876 5124
rect 218932 5068 218942 5124
rect 327506 5068 327516 5124
rect 327572 5068 328412 5124
rect 328468 5068 328478 5124
rect 15362 4956 15372 5012
rect 15428 4956 22652 5012
rect 22708 4956 22718 5012
rect 41906 4956 41916 5012
rect 41972 4956 44492 5012
rect 44548 4956 44558 5012
rect 149426 4956 149436 5012
rect 149492 4956 150332 5012
rect 150388 4956 150398 5012
rect 184706 4956 184716 5012
rect 184772 4956 185612 5012
rect 185668 4956 185678 5012
rect 325714 4956 325724 5012
rect 325780 4956 363356 5012
rect 363412 4956 363422 5012
rect 377122 4956 377132 5012
rect 377188 4956 387548 5012
rect 387604 4956 387614 5012
rect 536722 4956 536732 5012
rect 536788 4956 538748 5012
rect 538804 4956 538814 5012
rect 560242 4956 560252 5012
rect 560308 4956 561596 5012
rect 561652 4956 561662 5012
rect 354274 4844 354284 4900
rect 354340 4844 376796 4900
rect 376852 4844 376862 4900
rect 62850 4732 62860 4788
rect 62916 4732 68012 4788
rect 68068 4732 68078 4788
rect 85810 4732 85820 4788
rect 85876 4732 250460 4788
rect 250516 4732 250526 4788
rect 348562 4732 348572 4788
rect 348628 4732 374108 4788
rect 374164 4732 374174 4788
rect 380930 4732 380940 4788
rect 380996 4732 389340 4788
rect 389396 4732 389406 4788
rect 402770 4732 402780 4788
rect 402836 4732 409276 4788
rect 409332 4732 409342 4788
rect 491362 4732 491372 4788
rect 491428 4732 493052 4788
rect 493108 4732 493118 4788
rect 501442 4732 501452 4788
rect 501508 4732 508284 4788
rect 508340 4732 508350 4788
rect 51538 4620 51548 4676
rect 51604 4620 233548 4676
rect 233604 4620 233614 4676
rect 342850 4620 342860 4676
rect 342916 4620 371308 4676
rect 371364 4620 371374 4676
rect 408146 4620 408156 4676
rect 408212 4620 420700 4676
rect 420756 4620 420766 4676
rect 462802 4620 462812 4676
rect 462868 4620 536844 4676
rect 536900 4620 536910 4676
rect 43922 4508 43932 4564
rect 43988 4508 230748 4564
rect 230804 4508 230814 4564
rect 337138 4508 337148 4564
rect 337204 4508 368732 4564
rect 368788 4508 368798 4564
rect 371410 4508 371420 4564
rect 371476 4508 384860 4564
rect 384916 4508 384926 4564
rect 410834 4508 410844 4564
rect 410900 4508 426412 4564
rect 426468 4508 426478 4564
rect 465490 4508 465500 4564
rect 465556 4508 542668 4564
rect 542724 4508 542734 4564
rect 36306 4396 36316 4452
rect 36372 4396 227164 4452
rect 227220 4396 227230 4452
rect 331426 4396 331436 4452
rect 331492 4396 366044 4452
rect 366100 4396 366110 4452
rect 369506 4396 369516 4452
rect 369572 4396 383964 4452
rect 384020 4396 384030 4452
rect 404002 4396 404012 4452
rect 404068 4396 405468 4452
rect 405524 4396 405534 4452
rect 406354 4396 406364 4452
rect 406420 4396 416892 4452
rect 416948 4396 416958 4452
rect 417106 4396 417116 4452
rect 417172 4396 439740 4452
rect 439796 4396 439806 4452
rect 468178 4396 468188 4452
rect 468244 4396 540204 4452
rect 540260 4396 540270 4452
rect 541874 4396 541884 4452
rect 541940 4396 546364 4452
rect 546420 4396 546430 4452
rect 570322 4396 570332 4452
rect 570388 4396 584444 4452
rect 584500 4396 584510 4452
rect 22978 4284 22988 4340
rect 23044 4284 27692 4340
rect 27748 4284 27758 4340
rect 28690 4284 28700 4340
rect 28756 4284 223580 4340
rect 223636 4284 223646 4340
rect 363794 4284 363804 4340
rect 363860 4284 379820 4340
rect 379876 4284 379886 4340
rect 382834 4284 382844 4340
rect 382900 4284 390348 4340
rect 390404 4284 390414 4340
rect 392354 4284 392364 4340
rect 392420 4284 394716 4340
rect 394772 4284 394782 4340
rect 407250 4284 407260 4340
rect 407316 4284 418796 4340
rect 418852 4284 418862 4340
rect 419794 4284 419804 4340
rect 419860 4284 445452 4340
rect 445508 4284 445518 4340
rect 473554 4284 473564 4340
rect 473620 4284 559692 4340
rect 559748 4284 559758 4340
rect 563714 4284 563724 4340
rect 563780 4284 593068 4340
rect 593124 4284 593134 4340
rect 26786 4172 26796 4228
rect 26852 4172 29372 4228
rect 29428 4172 29438 4228
rect 31892 4172 219996 4228
rect 220052 4172 220062 4228
rect 224802 4172 224812 4228
rect 224868 4172 225932 4228
rect 225988 4172 225998 4228
rect 251458 4172 251468 4228
rect 251524 4172 252812 4228
rect 252868 4172 252878 4228
rect 259074 4172 259084 4228
rect 259140 4172 261212 4228
rect 261268 4172 261278 4228
rect 264786 4172 264796 4228
rect 264852 4172 266252 4228
rect 266308 4172 266318 4228
rect 272402 4172 272412 4228
rect 272468 4172 274764 4228
rect 274820 4172 274830 4228
rect 320002 4172 320012 4228
rect 320068 4172 360668 4228
rect 360724 4172 360734 4228
rect 367602 4172 367612 4228
rect 367668 4172 383068 4228
rect 383124 4172 383134 4228
rect 388546 4172 388556 4228
rect 388612 4172 392924 4228
rect 392980 4172 392990 4228
rect 394258 4172 394268 4228
rect 394324 4172 395612 4228
rect 395668 4172 395678 4228
rect 400642 4172 400652 4228
rect 400708 4172 401660 4228
rect 401716 4172 401726 4228
rect 402322 4172 402332 4228
rect 402388 4172 403564 4228
rect 403620 4172 403630 4228
rect 409042 4172 409052 4228
rect 409108 4172 422604 4228
rect 422660 4172 422670 4228
rect 425170 4172 425180 4228
rect 425236 4172 456988 4228
rect 457044 4172 457054 4228
rect 476242 4172 476252 4228
rect 476308 4172 565404 4228
rect 565460 4172 565470 4228
rect 567522 4172 567532 4228
rect 567588 4172 593964 4228
rect 594020 4172 594030 4228
rect 31892 4116 31948 4172
rect 21074 4060 21084 4116
rect 21140 4060 31948 4116
rect 40114 4060 40124 4116
rect 40180 4060 41132 4116
rect 41188 4060 41198 4116
rect 61058 4060 61068 4116
rect 61124 4060 62972 4116
rect 63028 4060 63038 4116
rect 68674 4060 68684 4116
rect 68740 4060 71372 4116
rect 71428 4060 71438 4116
rect 74386 4060 74396 4116
rect 74452 4060 78092 4116
rect 78148 4060 78158 4116
rect 80098 4060 80108 4116
rect 80164 4060 84812 4116
rect 84868 4060 84878 4116
rect 97234 4060 97244 4116
rect 97300 4060 99932 4116
rect 99988 4060 99998 4116
rect 112466 4060 112476 4116
rect 112532 4060 113484 4116
rect 113540 4060 113550 4116
rect 142706 4060 142716 4116
rect 142772 4060 146524 4116
rect 146580 4060 146590 4116
rect 154466 4060 154476 4116
rect 154532 4060 156044 4116
rect 156100 4060 156110 4116
rect 169586 4060 169596 4116
rect 169652 4060 170492 4116
rect 170548 4060 170558 4116
rect 186722 4060 186732 4116
rect 186788 4060 188972 4116
rect 189028 4060 189038 4116
rect 190530 4060 190540 4116
rect 190596 4060 194012 4116
rect 194068 4060 194078 4116
rect 205762 4060 205772 4116
rect 205828 4060 207452 4116
rect 207508 4060 207518 4116
rect 401874 4060 401884 4116
rect 401940 4060 407372 4116
rect 407428 4060 407438 4116
rect 499762 4060 499772 4116
rect 499828 4060 500668 4116
rect 500724 4060 500734 4116
rect 518354 4060 518364 4116
rect 518420 4060 525420 4116
rect 525476 4060 525486 4116
rect 531346 4060 531356 4116
rect 531412 4060 534268 4116
rect 534324 4060 534334 4116
rect 540194 4060 540204 4116
rect 540260 4060 548268 4116
rect 548324 4060 548334 4116
rect 403666 3948 403676 4004
rect 403732 3948 411180 4004
rect 411236 3948 411246 4004
rect 514210 3612 514220 3668
rect 514276 3612 519148 3668
rect 519204 3612 519214 3668
rect 314290 3500 314300 3556
rect 314356 3500 316652 3556
rect 316708 3500 316718 3556
rect 241826 2716 241836 2772
rect 241892 2716 314972 2772
rect 315028 2716 315038 2772
rect 222898 2604 222908 2660
rect 222964 2604 314188 2660
rect 314244 2604 314254 2660
rect 114370 2492 114380 2548
rect 114436 2492 263788 2548
rect 263844 2492 263854 2548
rect 295250 2492 295260 2548
rect 295316 2492 340172 2548
rect 340228 2492 340238 2548
rect 245858 28 245868 84
rect 245924 28 324268 84
rect 324324 28 324334 84
<< via3 >>
rect 467180 499324 467236 499380
rect 412860 499100 412916 499156
rect 413308 499100 413364 499156
rect 467180 498988 467236 499044
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 3154 597212 3774 598268
rect 3154 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 3774 597212
rect 3154 597088 3774 597156
rect 3154 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 3774 597088
rect 3154 596964 3774 597032
rect 3154 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 3774 596964
rect 3154 596840 3774 596908
rect 3154 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 3774 596840
rect 3154 580350 3774 596784
rect 3154 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 3774 580350
rect 3154 580226 3774 580294
rect 3154 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 3774 580226
rect 3154 580102 3774 580170
rect 3154 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 3774 580102
rect 3154 579978 3774 580046
rect 3154 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 3774 579978
rect 3154 562350 3774 579922
rect 3154 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 3774 562350
rect 3154 562226 3774 562294
rect 3154 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 3774 562226
rect 3154 562102 3774 562170
rect 3154 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 3774 562102
rect 3154 561978 3774 562046
rect 3154 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 3774 561978
rect 3154 544350 3774 561922
rect 3154 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 3774 544350
rect 3154 544226 3774 544294
rect 3154 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 3774 544226
rect 3154 544102 3774 544170
rect 3154 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 3774 544102
rect 3154 543978 3774 544046
rect 3154 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 3774 543978
rect 3154 526350 3774 543922
rect 3154 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 3774 526350
rect 3154 526226 3774 526294
rect 3154 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 3774 526226
rect 3154 526102 3774 526170
rect 3154 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 3774 526102
rect 3154 525978 3774 526046
rect 3154 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 3774 525978
rect 3154 508350 3774 525922
rect 3154 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 3774 508350
rect 3154 508226 3774 508294
rect 3154 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 3774 508226
rect 3154 508102 3774 508170
rect 3154 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 3774 508102
rect 3154 507978 3774 508046
rect 3154 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 3774 507978
rect 3154 490350 3774 507922
rect 3154 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 3774 490350
rect 3154 490226 3774 490294
rect 3154 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 3774 490226
rect 3154 490102 3774 490170
rect 3154 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 3774 490102
rect 3154 489978 3774 490046
rect 3154 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 3774 489978
rect 3154 472350 3774 489922
rect 3154 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 3774 472350
rect 3154 472226 3774 472294
rect 3154 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 3774 472226
rect 3154 472102 3774 472170
rect 3154 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 3774 472102
rect 3154 471978 3774 472046
rect 3154 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 3774 471978
rect 3154 454350 3774 471922
rect 3154 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 3774 454350
rect 3154 454226 3774 454294
rect 3154 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 3774 454226
rect 3154 454102 3774 454170
rect 3154 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 3774 454102
rect 3154 453978 3774 454046
rect 3154 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 3774 453978
rect 3154 436350 3774 453922
rect 3154 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 3774 436350
rect 3154 436226 3774 436294
rect 3154 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 3774 436226
rect 3154 436102 3774 436170
rect 3154 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 3774 436102
rect 3154 435978 3774 436046
rect 3154 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 3774 435978
rect 3154 418350 3774 435922
rect 3154 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 3774 418350
rect 3154 418226 3774 418294
rect 3154 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 3774 418226
rect 3154 418102 3774 418170
rect 3154 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 3774 418102
rect 3154 417978 3774 418046
rect 3154 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 3774 417978
rect 3154 400350 3774 417922
rect 3154 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 3774 400350
rect 3154 400226 3774 400294
rect 3154 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 3774 400226
rect 3154 400102 3774 400170
rect 3154 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 3774 400102
rect 3154 399978 3774 400046
rect 3154 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 3774 399978
rect 3154 382350 3774 399922
rect 3154 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 3774 382350
rect 3154 382226 3774 382294
rect 3154 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 3774 382226
rect 3154 382102 3774 382170
rect 3154 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 3774 382102
rect 3154 381978 3774 382046
rect 3154 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 3774 381978
rect 3154 364350 3774 381922
rect 3154 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 3774 364350
rect 3154 364226 3774 364294
rect 3154 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 3774 364226
rect 3154 364102 3774 364170
rect 3154 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 3774 364102
rect 3154 363978 3774 364046
rect 3154 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 3774 363978
rect 3154 346350 3774 363922
rect 3154 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 3774 346350
rect 3154 346226 3774 346294
rect 3154 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 3774 346226
rect 3154 346102 3774 346170
rect 3154 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 3774 346102
rect 3154 345978 3774 346046
rect 3154 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 3774 345978
rect 3154 328350 3774 345922
rect 3154 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 3774 328350
rect 3154 328226 3774 328294
rect 3154 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 3774 328226
rect 3154 328102 3774 328170
rect 3154 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 3774 328102
rect 3154 327978 3774 328046
rect 3154 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 3774 327978
rect 3154 310350 3774 327922
rect 3154 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 3774 310350
rect 3154 310226 3774 310294
rect 3154 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 3774 310226
rect 3154 310102 3774 310170
rect 3154 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 3774 310102
rect 3154 309978 3774 310046
rect 3154 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 3774 309978
rect 3154 292350 3774 309922
rect 3154 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 3774 292350
rect 3154 292226 3774 292294
rect 3154 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 3774 292226
rect 3154 292102 3774 292170
rect 3154 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 3774 292102
rect 3154 291978 3774 292046
rect 3154 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 3774 291978
rect 3154 274350 3774 291922
rect 3154 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 3774 274350
rect 3154 274226 3774 274294
rect 3154 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 3774 274226
rect 3154 274102 3774 274170
rect 3154 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 3774 274102
rect 3154 273978 3774 274046
rect 3154 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 3774 273978
rect 3154 256350 3774 273922
rect 3154 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 3774 256350
rect 3154 256226 3774 256294
rect 3154 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 3774 256226
rect 3154 256102 3774 256170
rect 3154 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 3774 256102
rect 3154 255978 3774 256046
rect 3154 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 3774 255978
rect 3154 238350 3774 255922
rect 3154 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 3774 238350
rect 3154 238226 3774 238294
rect 3154 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 3774 238226
rect 3154 238102 3774 238170
rect 3154 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 3774 238102
rect 3154 237978 3774 238046
rect 3154 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 3774 237978
rect 3154 220350 3774 237922
rect 3154 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 3774 220350
rect 3154 220226 3774 220294
rect 3154 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 3774 220226
rect 3154 220102 3774 220170
rect 3154 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 3774 220102
rect 3154 219978 3774 220046
rect 3154 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 3774 219978
rect 3154 202350 3774 219922
rect 3154 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 3774 202350
rect 3154 202226 3774 202294
rect 3154 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 3774 202226
rect 3154 202102 3774 202170
rect 3154 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 3774 202102
rect 3154 201978 3774 202046
rect 3154 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 3774 201978
rect 3154 184350 3774 201922
rect 3154 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 3774 184350
rect 3154 184226 3774 184294
rect 3154 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 3774 184226
rect 3154 184102 3774 184170
rect 3154 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 3774 184102
rect 3154 183978 3774 184046
rect 3154 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 3774 183978
rect 3154 166350 3774 183922
rect 3154 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 3774 166350
rect 3154 166226 3774 166294
rect 3154 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 3774 166226
rect 3154 166102 3774 166170
rect 3154 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 3774 166102
rect 3154 165978 3774 166046
rect 3154 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 3774 165978
rect 3154 148350 3774 165922
rect 3154 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 3774 148350
rect 3154 148226 3774 148294
rect 3154 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 3774 148226
rect 3154 148102 3774 148170
rect 3154 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 3774 148102
rect 3154 147978 3774 148046
rect 3154 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 3774 147978
rect 3154 130350 3774 147922
rect 3154 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 3774 130350
rect 3154 130226 3774 130294
rect 3154 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 3774 130226
rect 3154 130102 3774 130170
rect 3154 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 3774 130102
rect 3154 129978 3774 130046
rect 3154 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 3774 129978
rect 3154 112350 3774 129922
rect 3154 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 3774 112350
rect 3154 112226 3774 112294
rect 3154 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 3774 112226
rect 3154 112102 3774 112170
rect 3154 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 3774 112102
rect 3154 111978 3774 112046
rect 3154 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 3774 111978
rect 3154 94350 3774 111922
rect 3154 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 3774 94350
rect 3154 94226 3774 94294
rect 3154 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 3774 94226
rect 3154 94102 3774 94170
rect 3154 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 3774 94102
rect 3154 93978 3774 94046
rect 3154 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 3774 93978
rect 3154 76350 3774 93922
rect 3154 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 3774 76350
rect 3154 76226 3774 76294
rect 3154 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 3774 76226
rect 3154 76102 3774 76170
rect 3154 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 3774 76102
rect 3154 75978 3774 76046
rect 3154 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 3774 75978
rect 3154 58350 3774 75922
rect 3154 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 3774 58350
rect 3154 58226 3774 58294
rect 3154 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 3774 58226
rect 3154 58102 3774 58170
rect 3154 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 3774 58102
rect 3154 57978 3774 58046
rect 3154 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 3774 57978
rect 3154 40350 3774 57922
rect 3154 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 3774 40350
rect 3154 40226 3774 40294
rect 3154 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 3774 40226
rect 3154 40102 3774 40170
rect 3154 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 3774 40102
rect 3154 39978 3774 40046
rect 3154 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 3774 39978
rect 3154 22350 3774 39922
rect 3154 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 3774 22350
rect 3154 22226 3774 22294
rect 3154 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 3774 22226
rect 3154 22102 3774 22170
rect 3154 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 3774 22102
rect 3154 21978 3774 22046
rect 3154 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 3774 21978
rect 3154 4350 3774 21922
rect 3154 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 3774 4350
rect 3154 4226 3774 4294
rect 3154 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 3774 4226
rect 3154 4102 3774 4170
rect 3154 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 3774 4102
rect 3154 3978 3774 4046
rect 3154 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 3774 3978
rect 3154 -160 3774 3922
rect 3154 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 3774 -160
rect 3154 -284 3774 -216
rect 3154 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 3774 -284
rect 3154 -408 3774 -340
rect 3154 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 3774 -408
rect 3154 -532 3774 -464
rect 3154 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 3774 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 3154 -1644 3774 -588
rect 6874 598172 7494 598268
rect 6874 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 7494 598172
rect 6874 598048 7494 598116
rect 6874 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 7494 598048
rect 6874 597924 7494 597992
rect 6874 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 7494 597924
rect 6874 597800 7494 597868
rect 6874 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 7494 597800
rect 6874 586350 7494 597744
rect 6874 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 7494 586350
rect 6874 586226 7494 586294
rect 6874 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 7494 586226
rect 6874 586102 7494 586170
rect 6874 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 7494 586102
rect 6874 585978 7494 586046
rect 6874 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 7494 585978
rect 6874 568350 7494 585922
rect 6874 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 7494 568350
rect 6874 568226 7494 568294
rect 6874 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 7494 568226
rect 6874 568102 7494 568170
rect 6874 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 7494 568102
rect 6874 567978 7494 568046
rect 6874 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 7494 567978
rect 6874 550350 7494 567922
rect 6874 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 7494 550350
rect 6874 550226 7494 550294
rect 6874 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 7494 550226
rect 6874 550102 7494 550170
rect 6874 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 7494 550102
rect 6874 549978 7494 550046
rect 6874 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 7494 549978
rect 6874 532350 7494 549922
rect 6874 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 7494 532350
rect 6874 532226 7494 532294
rect 6874 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 7494 532226
rect 6874 532102 7494 532170
rect 6874 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 7494 532102
rect 6874 531978 7494 532046
rect 6874 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 7494 531978
rect 6874 514350 7494 531922
rect 6874 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 7494 514350
rect 6874 514226 7494 514294
rect 6874 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 7494 514226
rect 6874 514102 7494 514170
rect 6874 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 7494 514102
rect 6874 513978 7494 514046
rect 6874 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 7494 513978
rect 6874 496350 7494 513922
rect 6874 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 7494 496350
rect 6874 496226 7494 496294
rect 6874 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 7494 496226
rect 6874 496102 7494 496170
rect 6874 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 7494 496102
rect 6874 495978 7494 496046
rect 6874 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 7494 495978
rect 6874 478350 7494 495922
rect 6874 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 7494 478350
rect 6874 478226 7494 478294
rect 6874 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 7494 478226
rect 6874 478102 7494 478170
rect 6874 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 7494 478102
rect 6874 477978 7494 478046
rect 6874 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 7494 477978
rect 6874 460350 7494 477922
rect 6874 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 7494 460350
rect 6874 460226 7494 460294
rect 6874 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 7494 460226
rect 6874 460102 7494 460170
rect 6874 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 7494 460102
rect 6874 459978 7494 460046
rect 6874 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 7494 459978
rect 6874 442350 7494 459922
rect 6874 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 7494 442350
rect 6874 442226 7494 442294
rect 6874 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 7494 442226
rect 6874 442102 7494 442170
rect 6874 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 7494 442102
rect 6874 441978 7494 442046
rect 6874 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 7494 441978
rect 6874 424350 7494 441922
rect 6874 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 7494 424350
rect 6874 424226 7494 424294
rect 6874 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 7494 424226
rect 6874 424102 7494 424170
rect 6874 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 7494 424102
rect 6874 423978 7494 424046
rect 6874 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 7494 423978
rect 6874 406350 7494 423922
rect 6874 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 7494 406350
rect 6874 406226 7494 406294
rect 6874 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 7494 406226
rect 6874 406102 7494 406170
rect 6874 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 7494 406102
rect 6874 405978 7494 406046
rect 6874 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 7494 405978
rect 6874 388350 7494 405922
rect 6874 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 7494 388350
rect 6874 388226 7494 388294
rect 6874 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 7494 388226
rect 6874 388102 7494 388170
rect 6874 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 7494 388102
rect 6874 387978 7494 388046
rect 6874 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 7494 387978
rect 6874 370350 7494 387922
rect 6874 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 7494 370350
rect 6874 370226 7494 370294
rect 6874 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 7494 370226
rect 6874 370102 7494 370170
rect 6874 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 7494 370102
rect 6874 369978 7494 370046
rect 6874 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 7494 369978
rect 6874 352350 7494 369922
rect 6874 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 7494 352350
rect 6874 352226 7494 352294
rect 6874 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 7494 352226
rect 6874 352102 7494 352170
rect 6874 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 7494 352102
rect 6874 351978 7494 352046
rect 6874 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 7494 351978
rect 6874 334350 7494 351922
rect 6874 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 7494 334350
rect 6874 334226 7494 334294
rect 6874 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 7494 334226
rect 6874 334102 7494 334170
rect 6874 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 7494 334102
rect 6874 333978 7494 334046
rect 6874 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 7494 333978
rect 6874 316350 7494 333922
rect 6874 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 7494 316350
rect 6874 316226 7494 316294
rect 6874 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 7494 316226
rect 6874 316102 7494 316170
rect 6874 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 7494 316102
rect 6874 315978 7494 316046
rect 6874 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 7494 315978
rect 6874 298350 7494 315922
rect 6874 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 7494 298350
rect 6874 298226 7494 298294
rect 6874 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 7494 298226
rect 6874 298102 7494 298170
rect 6874 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 7494 298102
rect 6874 297978 7494 298046
rect 6874 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 7494 297978
rect 6874 280350 7494 297922
rect 6874 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 7494 280350
rect 6874 280226 7494 280294
rect 6874 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 7494 280226
rect 6874 280102 7494 280170
rect 6874 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 7494 280102
rect 6874 279978 7494 280046
rect 6874 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 7494 279978
rect 6874 262350 7494 279922
rect 6874 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 7494 262350
rect 6874 262226 7494 262294
rect 6874 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 7494 262226
rect 6874 262102 7494 262170
rect 6874 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 7494 262102
rect 6874 261978 7494 262046
rect 6874 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 7494 261978
rect 6874 244350 7494 261922
rect 6874 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 7494 244350
rect 6874 244226 7494 244294
rect 6874 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 7494 244226
rect 6874 244102 7494 244170
rect 6874 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 7494 244102
rect 6874 243978 7494 244046
rect 6874 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 7494 243978
rect 6874 226350 7494 243922
rect 6874 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 7494 226350
rect 6874 226226 7494 226294
rect 6874 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 7494 226226
rect 6874 226102 7494 226170
rect 6874 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 7494 226102
rect 6874 225978 7494 226046
rect 6874 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 7494 225978
rect 6874 208350 7494 225922
rect 6874 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 7494 208350
rect 6874 208226 7494 208294
rect 6874 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 7494 208226
rect 6874 208102 7494 208170
rect 6874 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 7494 208102
rect 6874 207978 7494 208046
rect 6874 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 7494 207978
rect 6874 190350 7494 207922
rect 6874 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 7494 190350
rect 6874 190226 7494 190294
rect 6874 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 7494 190226
rect 6874 190102 7494 190170
rect 6874 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 7494 190102
rect 6874 189978 7494 190046
rect 6874 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 7494 189978
rect 6874 172350 7494 189922
rect 6874 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 7494 172350
rect 6874 172226 7494 172294
rect 6874 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 7494 172226
rect 6874 172102 7494 172170
rect 6874 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 7494 172102
rect 6874 171978 7494 172046
rect 6874 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 7494 171978
rect 6874 154350 7494 171922
rect 6874 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 7494 154350
rect 6874 154226 7494 154294
rect 6874 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 7494 154226
rect 6874 154102 7494 154170
rect 6874 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 7494 154102
rect 6874 153978 7494 154046
rect 6874 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 7494 153978
rect 6874 136350 7494 153922
rect 6874 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 7494 136350
rect 6874 136226 7494 136294
rect 6874 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 7494 136226
rect 6874 136102 7494 136170
rect 6874 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 7494 136102
rect 6874 135978 7494 136046
rect 6874 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 7494 135978
rect 6874 118350 7494 135922
rect 6874 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 7494 118350
rect 6874 118226 7494 118294
rect 6874 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 7494 118226
rect 6874 118102 7494 118170
rect 6874 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 7494 118102
rect 6874 117978 7494 118046
rect 6874 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 7494 117978
rect 6874 100350 7494 117922
rect 6874 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 7494 100350
rect 6874 100226 7494 100294
rect 6874 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 7494 100226
rect 6874 100102 7494 100170
rect 6874 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 7494 100102
rect 6874 99978 7494 100046
rect 6874 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 7494 99978
rect 6874 82350 7494 99922
rect 6874 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 7494 82350
rect 6874 82226 7494 82294
rect 6874 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 7494 82226
rect 6874 82102 7494 82170
rect 6874 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 7494 82102
rect 6874 81978 7494 82046
rect 6874 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 7494 81978
rect 6874 64350 7494 81922
rect 6874 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 7494 64350
rect 6874 64226 7494 64294
rect 6874 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 7494 64226
rect 6874 64102 7494 64170
rect 6874 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 7494 64102
rect 6874 63978 7494 64046
rect 6874 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 7494 63978
rect 6874 46350 7494 63922
rect 6874 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 7494 46350
rect 6874 46226 7494 46294
rect 6874 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 7494 46226
rect 6874 46102 7494 46170
rect 6874 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 7494 46102
rect 6874 45978 7494 46046
rect 6874 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 7494 45978
rect 6874 28350 7494 45922
rect 6874 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 7494 28350
rect 6874 28226 7494 28294
rect 6874 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 7494 28226
rect 6874 28102 7494 28170
rect 6874 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 7494 28102
rect 6874 27978 7494 28046
rect 6874 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 7494 27978
rect 6874 10350 7494 27922
rect 6874 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 7494 10350
rect 6874 10226 7494 10294
rect 6874 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 7494 10226
rect 6874 10102 7494 10170
rect 6874 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 7494 10102
rect 6874 9978 7494 10046
rect 6874 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 7494 9978
rect 6874 -1120 7494 9922
rect 6874 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 7494 -1120
rect 6874 -1244 7494 -1176
rect 6874 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 7494 -1244
rect 6874 -1368 7494 -1300
rect 6874 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 7494 -1368
rect 6874 -1492 7494 -1424
rect 6874 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 7494 -1492
rect 6874 -1644 7494 -1548
rect 21154 597212 21774 598268
rect 21154 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 21774 597212
rect 21154 597088 21774 597156
rect 21154 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 21774 597088
rect 21154 596964 21774 597032
rect 21154 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 21774 596964
rect 21154 596840 21774 596908
rect 21154 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 21774 596840
rect 21154 580350 21774 596784
rect 21154 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 21774 580350
rect 21154 580226 21774 580294
rect 21154 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 21774 580226
rect 21154 580102 21774 580170
rect 21154 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 21774 580102
rect 21154 579978 21774 580046
rect 21154 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 21774 579978
rect 21154 562350 21774 579922
rect 21154 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 21774 562350
rect 21154 562226 21774 562294
rect 21154 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 21774 562226
rect 21154 562102 21774 562170
rect 21154 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 21774 562102
rect 21154 561978 21774 562046
rect 21154 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 21774 561978
rect 21154 544350 21774 561922
rect 21154 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 21774 544350
rect 21154 544226 21774 544294
rect 21154 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 21774 544226
rect 21154 544102 21774 544170
rect 21154 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 21774 544102
rect 21154 543978 21774 544046
rect 21154 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 21774 543978
rect 21154 526350 21774 543922
rect 21154 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 21774 526350
rect 21154 526226 21774 526294
rect 21154 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 21774 526226
rect 21154 526102 21774 526170
rect 21154 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 21774 526102
rect 21154 525978 21774 526046
rect 21154 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 21774 525978
rect 21154 508350 21774 525922
rect 21154 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 21774 508350
rect 21154 508226 21774 508294
rect 21154 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 21774 508226
rect 21154 508102 21774 508170
rect 21154 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 21774 508102
rect 21154 507978 21774 508046
rect 21154 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 21774 507978
rect 21154 490350 21774 507922
rect 21154 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 21774 490350
rect 21154 490226 21774 490294
rect 21154 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 21774 490226
rect 21154 490102 21774 490170
rect 21154 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 21774 490102
rect 21154 489978 21774 490046
rect 21154 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 21774 489978
rect 21154 472350 21774 489922
rect 21154 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 21774 472350
rect 21154 472226 21774 472294
rect 21154 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 21774 472226
rect 21154 472102 21774 472170
rect 21154 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 21774 472102
rect 21154 471978 21774 472046
rect 21154 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 21774 471978
rect 21154 454350 21774 471922
rect 21154 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 21774 454350
rect 21154 454226 21774 454294
rect 21154 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 21774 454226
rect 21154 454102 21774 454170
rect 21154 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 21774 454102
rect 21154 453978 21774 454046
rect 21154 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 21774 453978
rect 21154 436350 21774 453922
rect 21154 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 21774 436350
rect 21154 436226 21774 436294
rect 21154 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 21774 436226
rect 21154 436102 21774 436170
rect 21154 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 21774 436102
rect 21154 435978 21774 436046
rect 21154 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 21774 435978
rect 21154 418350 21774 435922
rect 21154 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 21774 418350
rect 21154 418226 21774 418294
rect 21154 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 21774 418226
rect 21154 418102 21774 418170
rect 21154 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 21774 418102
rect 21154 417978 21774 418046
rect 21154 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 21774 417978
rect 21154 400350 21774 417922
rect 21154 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 21774 400350
rect 21154 400226 21774 400294
rect 21154 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 21774 400226
rect 21154 400102 21774 400170
rect 21154 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 21774 400102
rect 21154 399978 21774 400046
rect 21154 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 21774 399978
rect 21154 382350 21774 399922
rect 21154 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 21774 382350
rect 21154 382226 21774 382294
rect 21154 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 21774 382226
rect 21154 382102 21774 382170
rect 21154 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 21774 382102
rect 21154 381978 21774 382046
rect 21154 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 21774 381978
rect 21154 364350 21774 381922
rect 21154 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 21774 364350
rect 21154 364226 21774 364294
rect 21154 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 21774 364226
rect 21154 364102 21774 364170
rect 21154 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 21774 364102
rect 21154 363978 21774 364046
rect 21154 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 21774 363978
rect 21154 346350 21774 363922
rect 21154 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 21774 346350
rect 21154 346226 21774 346294
rect 21154 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 21774 346226
rect 21154 346102 21774 346170
rect 21154 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 21774 346102
rect 21154 345978 21774 346046
rect 21154 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 21774 345978
rect 21154 328350 21774 345922
rect 21154 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 21774 328350
rect 21154 328226 21774 328294
rect 21154 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 21774 328226
rect 21154 328102 21774 328170
rect 21154 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 21774 328102
rect 21154 327978 21774 328046
rect 21154 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 21774 327978
rect 21154 310350 21774 327922
rect 21154 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 21774 310350
rect 21154 310226 21774 310294
rect 21154 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 21774 310226
rect 21154 310102 21774 310170
rect 21154 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 21774 310102
rect 21154 309978 21774 310046
rect 21154 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 21774 309978
rect 21154 292350 21774 309922
rect 21154 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 21774 292350
rect 21154 292226 21774 292294
rect 21154 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 21774 292226
rect 21154 292102 21774 292170
rect 21154 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 21774 292102
rect 21154 291978 21774 292046
rect 21154 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 21774 291978
rect 21154 274350 21774 291922
rect 21154 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 21774 274350
rect 21154 274226 21774 274294
rect 21154 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 21774 274226
rect 21154 274102 21774 274170
rect 21154 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 21774 274102
rect 21154 273978 21774 274046
rect 21154 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 21774 273978
rect 21154 256350 21774 273922
rect 21154 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 21774 256350
rect 21154 256226 21774 256294
rect 21154 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 21774 256226
rect 21154 256102 21774 256170
rect 21154 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 21774 256102
rect 21154 255978 21774 256046
rect 21154 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 21774 255978
rect 21154 238350 21774 255922
rect 21154 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 21774 238350
rect 21154 238226 21774 238294
rect 21154 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 21774 238226
rect 21154 238102 21774 238170
rect 21154 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 21774 238102
rect 21154 237978 21774 238046
rect 21154 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 21774 237978
rect 21154 220350 21774 237922
rect 21154 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 21774 220350
rect 21154 220226 21774 220294
rect 21154 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 21774 220226
rect 21154 220102 21774 220170
rect 21154 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 21774 220102
rect 21154 219978 21774 220046
rect 21154 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 21774 219978
rect 21154 202350 21774 219922
rect 21154 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 21774 202350
rect 21154 202226 21774 202294
rect 21154 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 21774 202226
rect 21154 202102 21774 202170
rect 21154 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 21774 202102
rect 21154 201978 21774 202046
rect 21154 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 21774 201978
rect 21154 184350 21774 201922
rect 21154 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 21774 184350
rect 21154 184226 21774 184294
rect 21154 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 21774 184226
rect 21154 184102 21774 184170
rect 21154 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 21774 184102
rect 21154 183978 21774 184046
rect 21154 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 21774 183978
rect 21154 166350 21774 183922
rect 21154 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 21774 166350
rect 21154 166226 21774 166294
rect 21154 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 21774 166226
rect 21154 166102 21774 166170
rect 21154 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 21774 166102
rect 21154 165978 21774 166046
rect 21154 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 21774 165978
rect 21154 148350 21774 165922
rect 21154 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 21774 148350
rect 21154 148226 21774 148294
rect 21154 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 21774 148226
rect 21154 148102 21774 148170
rect 21154 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 21774 148102
rect 21154 147978 21774 148046
rect 21154 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 21774 147978
rect 21154 130350 21774 147922
rect 21154 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 21774 130350
rect 21154 130226 21774 130294
rect 21154 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 21774 130226
rect 21154 130102 21774 130170
rect 21154 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 21774 130102
rect 21154 129978 21774 130046
rect 21154 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 21774 129978
rect 21154 112350 21774 129922
rect 21154 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 21774 112350
rect 21154 112226 21774 112294
rect 21154 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 21774 112226
rect 21154 112102 21774 112170
rect 21154 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 21774 112102
rect 21154 111978 21774 112046
rect 21154 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 21774 111978
rect 21154 94350 21774 111922
rect 21154 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 21774 94350
rect 21154 94226 21774 94294
rect 21154 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 21774 94226
rect 21154 94102 21774 94170
rect 21154 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 21774 94102
rect 21154 93978 21774 94046
rect 21154 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 21774 93978
rect 21154 76350 21774 93922
rect 21154 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 21774 76350
rect 21154 76226 21774 76294
rect 21154 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 21774 76226
rect 21154 76102 21774 76170
rect 21154 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 21774 76102
rect 21154 75978 21774 76046
rect 21154 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 21774 75978
rect 21154 58350 21774 75922
rect 21154 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 21774 58350
rect 21154 58226 21774 58294
rect 21154 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 21774 58226
rect 21154 58102 21774 58170
rect 21154 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 21774 58102
rect 21154 57978 21774 58046
rect 21154 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 21774 57978
rect 21154 40350 21774 57922
rect 21154 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 21774 40350
rect 21154 40226 21774 40294
rect 21154 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 21774 40226
rect 21154 40102 21774 40170
rect 21154 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 21774 40102
rect 21154 39978 21774 40046
rect 21154 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 21774 39978
rect 21154 22350 21774 39922
rect 21154 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 21774 22350
rect 21154 22226 21774 22294
rect 21154 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 21774 22226
rect 21154 22102 21774 22170
rect 21154 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 21774 22102
rect 21154 21978 21774 22046
rect 21154 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 21774 21978
rect 21154 4350 21774 21922
rect 21154 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 21774 4350
rect 21154 4226 21774 4294
rect 21154 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 21774 4226
rect 21154 4102 21774 4170
rect 21154 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 21774 4102
rect 21154 3978 21774 4046
rect 21154 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 21774 3978
rect 21154 -160 21774 3922
rect 21154 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 21774 -160
rect 21154 -284 21774 -216
rect 21154 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 21774 -284
rect 21154 -408 21774 -340
rect 21154 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 21774 -408
rect 21154 -532 21774 -464
rect 21154 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 21774 -532
rect 21154 -1644 21774 -588
rect 24874 598172 25494 598268
rect 24874 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 25494 598172
rect 24874 598048 25494 598116
rect 24874 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 25494 598048
rect 24874 597924 25494 597992
rect 24874 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 25494 597924
rect 24874 597800 25494 597868
rect 24874 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 25494 597800
rect 24874 586350 25494 597744
rect 24874 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 25494 586350
rect 24874 586226 25494 586294
rect 24874 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 25494 586226
rect 24874 586102 25494 586170
rect 24874 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 25494 586102
rect 24874 585978 25494 586046
rect 24874 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 25494 585978
rect 24874 568350 25494 585922
rect 24874 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 25494 568350
rect 24874 568226 25494 568294
rect 24874 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 25494 568226
rect 24874 568102 25494 568170
rect 24874 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 25494 568102
rect 24874 567978 25494 568046
rect 24874 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 25494 567978
rect 24874 550350 25494 567922
rect 24874 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 25494 550350
rect 24874 550226 25494 550294
rect 24874 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 25494 550226
rect 24874 550102 25494 550170
rect 24874 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 25494 550102
rect 24874 549978 25494 550046
rect 24874 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 25494 549978
rect 24874 532350 25494 549922
rect 24874 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 25494 532350
rect 24874 532226 25494 532294
rect 24874 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 25494 532226
rect 24874 532102 25494 532170
rect 24874 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 25494 532102
rect 24874 531978 25494 532046
rect 24874 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 25494 531978
rect 24874 514350 25494 531922
rect 24874 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 25494 514350
rect 24874 514226 25494 514294
rect 24874 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 25494 514226
rect 24874 514102 25494 514170
rect 24874 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 25494 514102
rect 24874 513978 25494 514046
rect 24874 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 25494 513978
rect 24874 496350 25494 513922
rect 24874 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 25494 496350
rect 24874 496226 25494 496294
rect 24874 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 25494 496226
rect 24874 496102 25494 496170
rect 24874 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 25494 496102
rect 24874 495978 25494 496046
rect 24874 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 25494 495978
rect 24874 478350 25494 495922
rect 24874 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 25494 478350
rect 24874 478226 25494 478294
rect 24874 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 25494 478226
rect 24874 478102 25494 478170
rect 24874 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 25494 478102
rect 24874 477978 25494 478046
rect 24874 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 25494 477978
rect 24874 460350 25494 477922
rect 24874 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 25494 460350
rect 24874 460226 25494 460294
rect 24874 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 25494 460226
rect 24874 460102 25494 460170
rect 24874 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 25494 460102
rect 24874 459978 25494 460046
rect 24874 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 25494 459978
rect 24874 442350 25494 459922
rect 24874 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 25494 442350
rect 24874 442226 25494 442294
rect 24874 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 25494 442226
rect 24874 442102 25494 442170
rect 24874 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 25494 442102
rect 24874 441978 25494 442046
rect 24874 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 25494 441978
rect 24874 424350 25494 441922
rect 24874 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 25494 424350
rect 24874 424226 25494 424294
rect 24874 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 25494 424226
rect 24874 424102 25494 424170
rect 24874 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 25494 424102
rect 24874 423978 25494 424046
rect 24874 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 25494 423978
rect 24874 406350 25494 423922
rect 24874 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 25494 406350
rect 24874 406226 25494 406294
rect 24874 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 25494 406226
rect 24874 406102 25494 406170
rect 24874 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 25494 406102
rect 24874 405978 25494 406046
rect 24874 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 25494 405978
rect 24874 388350 25494 405922
rect 24874 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 25494 388350
rect 24874 388226 25494 388294
rect 24874 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 25494 388226
rect 24874 388102 25494 388170
rect 24874 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 25494 388102
rect 24874 387978 25494 388046
rect 24874 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 25494 387978
rect 24874 370350 25494 387922
rect 24874 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 25494 370350
rect 24874 370226 25494 370294
rect 24874 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 25494 370226
rect 24874 370102 25494 370170
rect 24874 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 25494 370102
rect 24874 369978 25494 370046
rect 24874 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 25494 369978
rect 24874 352350 25494 369922
rect 24874 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 25494 352350
rect 24874 352226 25494 352294
rect 24874 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 25494 352226
rect 24874 352102 25494 352170
rect 24874 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 25494 352102
rect 24874 351978 25494 352046
rect 24874 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 25494 351978
rect 24874 334350 25494 351922
rect 24874 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 25494 334350
rect 24874 334226 25494 334294
rect 24874 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 25494 334226
rect 24874 334102 25494 334170
rect 24874 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 25494 334102
rect 24874 333978 25494 334046
rect 24874 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 25494 333978
rect 24874 316350 25494 333922
rect 24874 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 25494 316350
rect 24874 316226 25494 316294
rect 24874 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 25494 316226
rect 24874 316102 25494 316170
rect 24874 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 25494 316102
rect 24874 315978 25494 316046
rect 24874 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 25494 315978
rect 24874 298350 25494 315922
rect 24874 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 25494 298350
rect 24874 298226 25494 298294
rect 24874 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 25494 298226
rect 24874 298102 25494 298170
rect 24874 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 25494 298102
rect 24874 297978 25494 298046
rect 24874 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 25494 297978
rect 24874 280350 25494 297922
rect 24874 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 25494 280350
rect 24874 280226 25494 280294
rect 24874 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 25494 280226
rect 24874 280102 25494 280170
rect 24874 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 25494 280102
rect 24874 279978 25494 280046
rect 24874 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 25494 279978
rect 24874 262350 25494 279922
rect 24874 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 25494 262350
rect 24874 262226 25494 262294
rect 24874 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 25494 262226
rect 24874 262102 25494 262170
rect 24874 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 25494 262102
rect 24874 261978 25494 262046
rect 24874 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 25494 261978
rect 24874 244350 25494 261922
rect 24874 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 25494 244350
rect 24874 244226 25494 244294
rect 24874 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 25494 244226
rect 24874 244102 25494 244170
rect 24874 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 25494 244102
rect 24874 243978 25494 244046
rect 24874 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 25494 243978
rect 24874 226350 25494 243922
rect 24874 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 25494 226350
rect 24874 226226 25494 226294
rect 24874 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 25494 226226
rect 24874 226102 25494 226170
rect 24874 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 25494 226102
rect 24874 225978 25494 226046
rect 24874 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 25494 225978
rect 24874 208350 25494 225922
rect 24874 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 25494 208350
rect 24874 208226 25494 208294
rect 24874 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 25494 208226
rect 24874 208102 25494 208170
rect 24874 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 25494 208102
rect 24874 207978 25494 208046
rect 24874 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 25494 207978
rect 24874 190350 25494 207922
rect 24874 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 25494 190350
rect 24874 190226 25494 190294
rect 24874 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 25494 190226
rect 24874 190102 25494 190170
rect 24874 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 25494 190102
rect 24874 189978 25494 190046
rect 24874 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 25494 189978
rect 24874 172350 25494 189922
rect 24874 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 25494 172350
rect 24874 172226 25494 172294
rect 24874 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 25494 172226
rect 24874 172102 25494 172170
rect 24874 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 25494 172102
rect 24874 171978 25494 172046
rect 24874 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 25494 171978
rect 24874 154350 25494 171922
rect 24874 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 25494 154350
rect 24874 154226 25494 154294
rect 24874 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 25494 154226
rect 24874 154102 25494 154170
rect 24874 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 25494 154102
rect 24874 153978 25494 154046
rect 24874 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 25494 153978
rect 24874 136350 25494 153922
rect 24874 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 25494 136350
rect 24874 136226 25494 136294
rect 24874 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 25494 136226
rect 24874 136102 25494 136170
rect 24874 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 25494 136102
rect 24874 135978 25494 136046
rect 24874 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 25494 135978
rect 24874 118350 25494 135922
rect 24874 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 25494 118350
rect 24874 118226 25494 118294
rect 24874 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 25494 118226
rect 24874 118102 25494 118170
rect 24874 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 25494 118102
rect 24874 117978 25494 118046
rect 24874 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 25494 117978
rect 24874 100350 25494 117922
rect 24874 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 25494 100350
rect 24874 100226 25494 100294
rect 24874 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 25494 100226
rect 24874 100102 25494 100170
rect 24874 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 25494 100102
rect 24874 99978 25494 100046
rect 24874 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 25494 99978
rect 24874 82350 25494 99922
rect 24874 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 25494 82350
rect 24874 82226 25494 82294
rect 24874 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 25494 82226
rect 24874 82102 25494 82170
rect 24874 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 25494 82102
rect 24874 81978 25494 82046
rect 24874 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 25494 81978
rect 24874 64350 25494 81922
rect 24874 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 25494 64350
rect 24874 64226 25494 64294
rect 24874 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 25494 64226
rect 24874 64102 25494 64170
rect 24874 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 25494 64102
rect 24874 63978 25494 64046
rect 24874 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 25494 63978
rect 24874 46350 25494 63922
rect 24874 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 25494 46350
rect 24874 46226 25494 46294
rect 24874 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 25494 46226
rect 24874 46102 25494 46170
rect 24874 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 25494 46102
rect 24874 45978 25494 46046
rect 24874 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 25494 45978
rect 24874 28350 25494 45922
rect 24874 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 25494 28350
rect 24874 28226 25494 28294
rect 24874 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 25494 28226
rect 24874 28102 25494 28170
rect 24874 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 25494 28102
rect 24874 27978 25494 28046
rect 24874 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 25494 27978
rect 24874 10350 25494 27922
rect 24874 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 25494 10350
rect 24874 10226 25494 10294
rect 24874 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 25494 10226
rect 24874 10102 25494 10170
rect 24874 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 25494 10102
rect 24874 9978 25494 10046
rect 24874 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 25494 9978
rect 24874 -1120 25494 9922
rect 24874 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 25494 -1120
rect 24874 -1244 25494 -1176
rect 24874 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 25494 -1244
rect 24874 -1368 25494 -1300
rect 24874 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 25494 -1368
rect 24874 -1492 25494 -1424
rect 24874 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 25494 -1492
rect 24874 -1644 25494 -1548
rect 39154 597212 39774 598268
rect 39154 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 39774 597212
rect 39154 597088 39774 597156
rect 39154 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 39774 597088
rect 39154 596964 39774 597032
rect 39154 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 39774 596964
rect 39154 596840 39774 596908
rect 39154 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 39774 596840
rect 39154 580350 39774 596784
rect 39154 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 39774 580350
rect 39154 580226 39774 580294
rect 39154 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 39774 580226
rect 39154 580102 39774 580170
rect 39154 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 39774 580102
rect 39154 579978 39774 580046
rect 39154 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 39774 579978
rect 39154 562350 39774 579922
rect 39154 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 39774 562350
rect 39154 562226 39774 562294
rect 39154 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 39774 562226
rect 39154 562102 39774 562170
rect 39154 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 39774 562102
rect 39154 561978 39774 562046
rect 39154 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 39774 561978
rect 39154 544350 39774 561922
rect 39154 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 39774 544350
rect 39154 544226 39774 544294
rect 39154 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 39774 544226
rect 39154 544102 39774 544170
rect 39154 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 39774 544102
rect 39154 543978 39774 544046
rect 39154 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 39774 543978
rect 39154 526350 39774 543922
rect 39154 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 39774 526350
rect 39154 526226 39774 526294
rect 39154 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 39774 526226
rect 39154 526102 39774 526170
rect 39154 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 39774 526102
rect 39154 525978 39774 526046
rect 39154 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 39774 525978
rect 39154 508350 39774 525922
rect 39154 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 39774 508350
rect 39154 508226 39774 508294
rect 39154 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 39774 508226
rect 39154 508102 39774 508170
rect 39154 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 39774 508102
rect 39154 507978 39774 508046
rect 39154 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 39774 507978
rect 39154 490350 39774 507922
rect 39154 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 39774 490350
rect 39154 490226 39774 490294
rect 39154 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 39774 490226
rect 39154 490102 39774 490170
rect 39154 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 39774 490102
rect 39154 489978 39774 490046
rect 39154 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 39774 489978
rect 39154 472350 39774 489922
rect 39154 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 39774 472350
rect 39154 472226 39774 472294
rect 39154 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 39774 472226
rect 39154 472102 39774 472170
rect 39154 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 39774 472102
rect 39154 471978 39774 472046
rect 39154 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 39774 471978
rect 39154 454350 39774 471922
rect 39154 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 39774 454350
rect 39154 454226 39774 454294
rect 39154 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 39774 454226
rect 39154 454102 39774 454170
rect 39154 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 39774 454102
rect 39154 453978 39774 454046
rect 39154 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 39774 453978
rect 39154 436350 39774 453922
rect 39154 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 39774 436350
rect 39154 436226 39774 436294
rect 39154 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 39774 436226
rect 39154 436102 39774 436170
rect 39154 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 39774 436102
rect 39154 435978 39774 436046
rect 39154 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 39774 435978
rect 39154 418350 39774 435922
rect 39154 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 39774 418350
rect 39154 418226 39774 418294
rect 39154 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 39774 418226
rect 39154 418102 39774 418170
rect 39154 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 39774 418102
rect 39154 417978 39774 418046
rect 39154 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 39774 417978
rect 39154 400350 39774 417922
rect 39154 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 39774 400350
rect 39154 400226 39774 400294
rect 39154 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 39774 400226
rect 39154 400102 39774 400170
rect 39154 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 39774 400102
rect 39154 399978 39774 400046
rect 39154 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 39774 399978
rect 39154 382350 39774 399922
rect 39154 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 39774 382350
rect 39154 382226 39774 382294
rect 39154 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 39774 382226
rect 39154 382102 39774 382170
rect 39154 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 39774 382102
rect 39154 381978 39774 382046
rect 39154 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 39774 381978
rect 39154 364350 39774 381922
rect 39154 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 39774 364350
rect 39154 364226 39774 364294
rect 39154 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 39774 364226
rect 39154 364102 39774 364170
rect 39154 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 39774 364102
rect 39154 363978 39774 364046
rect 39154 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 39774 363978
rect 39154 346350 39774 363922
rect 39154 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 39774 346350
rect 39154 346226 39774 346294
rect 39154 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 39774 346226
rect 39154 346102 39774 346170
rect 39154 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 39774 346102
rect 39154 345978 39774 346046
rect 39154 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 39774 345978
rect 39154 328350 39774 345922
rect 39154 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 39774 328350
rect 39154 328226 39774 328294
rect 39154 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 39774 328226
rect 39154 328102 39774 328170
rect 39154 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 39774 328102
rect 39154 327978 39774 328046
rect 39154 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 39774 327978
rect 39154 310350 39774 327922
rect 39154 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 39774 310350
rect 39154 310226 39774 310294
rect 39154 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 39774 310226
rect 39154 310102 39774 310170
rect 39154 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 39774 310102
rect 39154 309978 39774 310046
rect 39154 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 39774 309978
rect 39154 292350 39774 309922
rect 39154 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 39774 292350
rect 39154 292226 39774 292294
rect 39154 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 39774 292226
rect 39154 292102 39774 292170
rect 39154 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 39774 292102
rect 39154 291978 39774 292046
rect 39154 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 39774 291978
rect 39154 274350 39774 291922
rect 39154 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 39774 274350
rect 39154 274226 39774 274294
rect 39154 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 39774 274226
rect 39154 274102 39774 274170
rect 39154 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 39774 274102
rect 39154 273978 39774 274046
rect 39154 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 39774 273978
rect 39154 256350 39774 273922
rect 39154 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 39774 256350
rect 39154 256226 39774 256294
rect 39154 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 39774 256226
rect 39154 256102 39774 256170
rect 39154 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 39774 256102
rect 39154 255978 39774 256046
rect 39154 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 39774 255978
rect 39154 238350 39774 255922
rect 39154 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 39774 238350
rect 39154 238226 39774 238294
rect 39154 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 39774 238226
rect 39154 238102 39774 238170
rect 39154 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 39774 238102
rect 39154 237978 39774 238046
rect 39154 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 39774 237978
rect 39154 220350 39774 237922
rect 39154 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 39774 220350
rect 39154 220226 39774 220294
rect 39154 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 39774 220226
rect 39154 220102 39774 220170
rect 39154 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 39774 220102
rect 39154 219978 39774 220046
rect 39154 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 39774 219978
rect 39154 202350 39774 219922
rect 39154 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 39774 202350
rect 39154 202226 39774 202294
rect 39154 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 39774 202226
rect 39154 202102 39774 202170
rect 39154 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 39774 202102
rect 39154 201978 39774 202046
rect 39154 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 39774 201978
rect 39154 184350 39774 201922
rect 39154 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 39774 184350
rect 39154 184226 39774 184294
rect 39154 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 39774 184226
rect 39154 184102 39774 184170
rect 39154 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 39774 184102
rect 39154 183978 39774 184046
rect 39154 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 39774 183978
rect 39154 166350 39774 183922
rect 39154 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 39774 166350
rect 39154 166226 39774 166294
rect 39154 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 39774 166226
rect 39154 166102 39774 166170
rect 39154 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 39774 166102
rect 39154 165978 39774 166046
rect 39154 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 39774 165978
rect 39154 148350 39774 165922
rect 39154 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 39774 148350
rect 39154 148226 39774 148294
rect 39154 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 39774 148226
rect 39154 148102 39774 148170
rect 39154 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 39774 148102
rect 39154 147978 39774 148046
rect 39154 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 39774 147978
rect 39154 130350 39774 147922
rect 39154 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 39774 130350
rect 39154 130226 39774 130294
rect 39154 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 39774 130226
rect 39154 130102 39774 130170
rect 39154 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 39774 130102
rect 39154 129978 39774 130046
rect 39154 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 39774 129978
rect 39154 112350 39774 129922
rect 39154 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 39774 112350
rect 39154 112226 39774 112294
rect 39154 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 39774 112226
rect 39154 112102 39774 112170
rect 39154 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 39774 112102
rect 39154 111978 39774 112046
rect 39154 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 39774 111978
rect 39154 94350 39774 111922
rect 39154 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 39774 94350
rect 39154 94226 39774 94294
rect 39154 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 39774 94226
rect 39154 94102 39774 94170
rect 39154 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 39774 94102
rect 39154 93978 39774 94046
rect 39154 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 39774 93978
rect 39154 76350 39774 93922
rect 39154 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 39774 76350
rect 39154 76226 39774 76294
rect 39154 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 39774 76226
rect 39154 76102 39774 76170
rect 39154 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 39774 76102
rect 39154 75978 39774 76046
rect 39154 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 39774 75978
rect 39154 58350 39774 75922
rect 39154 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 39774 58350
rect 39154 58226 39774 58294
rect 39154 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 39774 58226
rect 39154 58102 39774 58170
rect 39154 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 39774 58102
rect 39154 57978 39774 58046
rect 39154 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 39774 57978
rect 39154 40350 39774 57922
rect 39154 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 39774 40350
rect 39154 40226 39774 40294
rect 39154 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 39774 40226
rect 39154 40102 39774 40170
rect 39154 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 39774 40102
rect 39154 39978 39774 40046
rect 39154 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 39774 39978
rect 39154 22350 39774 39922
rect 39154 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 39774 22350
rect 39154 22226 39774 22294
rect 39154 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 39774 22226
rect 39154 22102 39774 22170
rect 39154 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 39774 22102
rect 39154 21978 39774 22046
rect 39154 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 39774 21978
rect 39154 4350 39774 21922
rect 39154 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 39774 4350
rect 39154 4226 39774 4294
rect 39154 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 39774 4226
rect 39154 4102 39774 4170
rect 39154 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 39774 4102
rect 39154 3978 39774 4046
rect 39154 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 39774 3978
rect 39154 -160 39774 3922
rect 39154 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 39774 -160
rect 39154 -284 39774 -216
rect 39154 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 39774 -284
rect 39154 -408 39774 -340
rect 39154 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 39774 -408
rect 39154 -532 39774 -464
rect 39154 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 39774 -532
rect 39154 -1644 39774 -588
rect 42874 598172 43494 598268
rect 42874 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 43494 598172
rect 42874 598048 43494 598116
rect 42874 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 43494 598048
rect 42874 597924 43494 597992
rect 42874 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 43494 597924
rect 42874 597800 43494 597868
rect 42874 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 43494 597800
rect 42874 586350 43494 597744
rect 42874 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 43494 586350
rect 42874 586226 43494 586294
rect 42874 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 43494 586226
rect 42874 586102 43494 586170
rect 42874 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 43494 586102
rect 42874 585978 43494 586046
rect 42874 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 43494 585978
rect 42874 568350 43494 585922
rect 42874 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 43494 568350
rect 42874 568226 43494 568294
rect 42874 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 43494 568226
rect 42874 568102 43494 568170
rect 42874 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 43494 568102
rect 42874 567978 43494 568046
rect 42874 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 43494 567978
rect 42874 550350 43494 567922
rect 42874 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 43494 550350
rect 42874 550226 43494 550294
rect 42874 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 43494 550226
rect 42874 550102 43494 550170
rect 42874 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 43494 550102
rect 42874 549978 43494 550046
rect 42874 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 43494 549978
rect 42874 532350 43494 549922
rect 42874 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 43494 532350
rect 42874 532226 43494 532294
rect 42874 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 43494 532226
rect 42874 532102 43494 532170
rect 42874 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 43494 532102
rect 42874 531978 43494 532046
rect 42874 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 43494 531978
rect 42874 514350 43494 531922
rect 42874 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 43494 514350
rect 42874 514226 43494 514294
rect 42874 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 43494 514226
rect 42874 514102 43494 514170
rect 42874 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 43494 514102
rect 42874 513978 43494 514046
rect 42874 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 43494 513978
rect 42874 496350 43494 513922
rect 42874 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 43494 496350
rect 42874 496226 43494 496294
rect 42874 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 43494 496226
rect 42874 496102 43494 496170
rect 42874 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 43494 496102
rect 42874 495978 43494 496046
rect 42874 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 43494 495978
rect 42874 478350 43494 495922
rect 42874 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 43494 478350
rect 42874 478226 43494 478294
rect 42874 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 43494 478226
rect 42874 478102 43494 478170
rect 42874 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 43494 478102
rect 42874 477978 43494 478046
rect 42874 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 43494 477978
rect 42874 460350 43494 477922
rect 42874 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 43494 460350
rect 42874 460226 43494 460294
rect 42874 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 43494 460226
rect 42874 460102 43494 460170
rect 42874 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 43494 460102
rect 42874 459978 43494 460046
rect 42874 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 43494 459978
rect 42874 442350 43494 459922
rect 42874 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 43494 442350
rect 42874 442226 43494 442294
rect 42874 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 43494 442226
rect 42874 442102 43494 442170
rect 42874 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 43494 442102
rect 42874 441978 43494 442046
rect 42874 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 43494 441978
rect 42874 424350 43494 441922
rect 42874 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 43494 424350
rect 42874 424226 43494 424294
rect 42874 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 43494 424226
rect 42874 424102 43494 424170
rect 42874 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 43494 424102
rect 42874 423978 43494 424046
rect 42874 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 43494 423978
rect 42874 406350 43494 423922
rect 42874 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 43494 406350
rect 42874 406226 43494 406294
rect 42874 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 43494 406226
rect 42874 406102 43494 406170
rect 42874 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 43494 406102
rect 42874 405978 43494 406046
rect 42874 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 43494 405978
rect 42874 388350 43494 405922
rect 42874 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 43494 388350
rect 42874 388226 43494 388294
rect 42874 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 43494 388226
rect 42874 388102 43494 388170
rect 42874 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 43494 388102
rect 42874 387978 43494 388046
rect 42874 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 43494 387978
rect 42874 370350 43494 387922
rect 42874 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 43494 370350
rect 42874 370226 43494 370294
rect 42874 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 43494 370226
rect 42874 370102 43494 370170
rect 42874 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 43494 370102
rect 42874 369978 43494 370046
rect 42874 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 43494 369978
rect 42874 352350 43494 369922
rect 42874 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 43494 352350
rect 42874 352226 43494 352294
rect 42874 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 43494 352226
rect 42874 352102 43494 352170
rect 42874 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 43494 352102
rect 42874 351978 43494 352046
rect 42874 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 43494 351978
rect 42874 334350 43494 351922
rect 42874 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 43494 334350
rect 42874 334226 43494 334294
rect 42874 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 43494 334226
rect 42874 334102 43494 334170
rect 42874 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 43494 334102
rect 42874 333978 43494 334046
rect 42874 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 43494 333978
rect 42874 316350 43494 333922
rect 42874 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 43494 316350
rect 42874 316226 43494 316294
rect 42874 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 43494 316226
rect 42874 316102 43494 316170
rect 42874 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 43494 316102
rect 42874 315978 43494 316046
rect 42874 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 43494 315978
rect 42874 298350 43494 315922
rect 42874 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 43494 298350
rect 42874 298226 43494 298294
rect 42874 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 43494 298226
rect 42874 298102 43494 298170
rect 42874 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 43494 298102
rect 42874 297978 43494 298046
rect 42874 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 43494 297978
rect 42874 280350 43494 297922
rect 42874 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 43494 280350
rect 42874 280226 43494 280294
rect 42874 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 43494 280226
rect 42874 280102 43494 280170
rect 42874 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 43494 280102
rect 42874 279978 43494 280046
rect 42874 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 43494 279978
rect 42874 262350 43494 279922
rect 42874 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 43494 262350
rect 42874 262226 43494 262294
rect 42874 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 43494 262226
rect 42874 262102 43494 262170
rect 42874 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 43494 262102
rect 42874 261978 43494 262046
rect 42874 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 43494 261978
rect 42874 244350 43494 261922
rect 42874 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 43494 244350
rect 42874 244226 43494 244294
rect 42874 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 43494 244226
rect 42874 244102 43494 244170
rect 42874 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 43494 244102
rect 42874 243978 43494 244046
rect 42874 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 43494 243978
rect 42874 226350 43494 243922
rect 42874 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 43494 226350
rect 42874 226226 43494 226294
rect 42874 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 43494 226226
rect 42874 226102 43494 226170
rect 42874 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 43494 226102
rect 42874 225978 43494 226046
rect 42874 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 43494 225978
rect 42874 208350 43494 225922
rect 42874 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 43494 208350
rect 42874 208226 43494 208294
rect 42874 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 43494 208226
rect 42874 208102 43494 208170
rect 42874 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 43494 208102
rect 42874 207978 43494 208046
rect 42874 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 43494 207978
rect 42874 190350 43494 207922
rect 42874 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 43494 190350
rect 42874 190226 43494 190294
rect 42874 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 43494 190226
rect 42874 190102 43494 190170
rect 42874 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 43494 190102
rect 42874 189978 43494 190046
rect 42874 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 43494 189978
rect 42874 172350 43494 189922
rect 42874 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 43494 172350
rect 42874 172226 43494 172294
rect 42874 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 43494 172226
rect 42874 172102 43494 172170
rect 42874 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 43494 172102
rect 42874 171978 43494 172046
rect 42874 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 43494 171978
rect 42874 154350 43494 171922
rect 42874 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 43494 154350
rect 42874 154226 43494 154294
rect 42874 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 43494 154226
rect 42874 154102 43494 154170
rect 42874 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 43494 154102
rect 42874 153978 43494 154046
rect 42874 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 43494 153978
rect 42874 136350 43494 153922
rect 42874 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 43494 136350
rect 42874 136226 43494 136294
rect 42874 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 43494 136226
rect 42874 136102 43494 136170
rect 42874 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 43494 136102
rect 42874 135978 43494 136046
rect 42874 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 43494 135978
rect 42874 118350 43494 135922
rect 42874 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 43494 118350
rect 42874 118226 43494 118294
rect 42874 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 43494 118226
rect 42874 118102 43494 118170
rect 42874 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 43494 118102
rect 42874 117978 43494 118046
rect 42874 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 43494 117978
rect 42874 100350 43494 117922
rect 42874 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 43494 100350
rect 42874 100226 43494 100294
rect 42874 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 43494 100226
rect 42874 100102 43494 100170
rect 42874 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 43494 100102
rect 42874 99978 43494 100046
rect 42874 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 43494 99978
rect 42874 82350 43494 99922
rect 42874 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 43494 82350
rect 42874 82226 43494 82294
rect 42874 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 43494 82226
rect 42874 82102 43494 82170
rect 42874 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 43494 82102
rect 42874 81978 43494 82046
rect 42874 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 43494 81978
rect 42874 64350 43494 81922
rect 42874 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 43494 64350
rect 42874 64226 43494 64294
rect 42874 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 43494 64226
rect 42874 64102 43494 64170
rect 42874 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 43494 64102
rect 42874 63978 43494 64046
rect 42874 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 43494 63978
rect 42874 46350 43494 63922
rect 42874 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 43494 46350
rect 42874 46226 43494 46294
rect 42874 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 43494 46226
rect 42874 46102 43494 46170
rect 42874 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 43494 46102
rect 42874 45978 43494 46046
rect 42874 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 43494 45978
rect 42874 28350 43494 45922
rect 42874 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 43494 28350
rect 42874 28226 43494 28294
rect 42874 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 43494 28226
rect 42874 28102 43494 28170
rect 42874 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 43494 28102
rect 42874 27978 43494 28046
rect 42874 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 43494 27978
rect 42874 10350 43494 27922
rect 42874 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 43494 10350
rect 42874 10226 43494 10294
rect 42874 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 43494 10226
rect 42874 10102 43494 10170
rect 42874 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 43494 10102
rect 42874 9978 43494 10046
rect 42874 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 43494 9978
rect 42874 -1120 43494 9922
rect 42874 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 43494 -1120
rect 42874 -1244 43494 -1176
rect 42874 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 43494 -1244
rect 42874 -1368 43494 -1300
rect 42874 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 43494 -1368
rect 42874 -1492 43494 -1424
rect 42874 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 43494 -1492
rect 42874 -1644 43494 -1548
rect 57154 597212 57774 598268
rect 57154 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 57774 597212
rect 57154 597088 57774 597156
rect 57154 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 57774 597088
rect 57154 596964 57774 597032
rect 57154 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 57774 596964
rect 57154 596840 57774 596908
rect 57154 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 57774 596840
rect 57154 580350 57774 596784
rect 57154 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 57774 580350
rect 57154 580226 57774 580294
rect 57154 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 57774 580226
rect 57154 580102 57774 580170
rect 57154 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 57774 580102
rect 57154 579978 57774 580046
rect 57154 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 57774 579978
rect 57154 562350 57774 579922
rect 57154 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 57774 562350
rect 57154 562226 57774 562294
rect 57154 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 57774 562226
rect 57154 562102 57774 562170
rect 57154 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 57774 562102
rect 57154 561978 57774 562046
rect 57154 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 57774 561978
rect 57154 544350 57774 561922
rect 57154 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 57774 544350
rect 57154 544226 57774 544294
rect 57154 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 57774 544226
rect 57154 544102 57774 544170
rect 57154 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 57774 544102
rect 57154 543978 57774 544046
rect 57154 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 57774 543978
rect 57154 526350 57774 543922
rect 57154 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 57774 526350
rect 57154 526226 57774 526294
rect 57154 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 57774 526226
rect 57154 526102 57774 526170
rect 57154 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 57774 526102
rect 57154 525978 57774 526046
rect 57154 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 57774 525978
rect 57154 508350 57774 525922
rect 57154 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 57774 508350
rect 57154 508226 57774 508294
rect 57154 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 57774 508226
rect 57154 508102 57774 508170
rect 57154 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 57774 508102
rect 57154 507978 57774 508046
rect 57154 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 57774 507978
rect 57154 490350 57774 507922
rect 57154 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 57774 490350
rect 57154 490226 57774 490294
rect 57154 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 57774 490226
rect 57154 490102 57774 490170
rect 57154 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 57774 490102
rect 57154 489978 57774 490046
rect 57154 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 57774 489978
rect 57154 472350 57774 489922
rect 57154 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 57774 472350
rect 57154 472226 57774 472294
rect 57154 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 57774 472226
rect 57154 472102 57774 472170
rect 57154 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 57774 472102
rect 57154 471978 57774 472046
rect 57154 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 57774 471978
rect 57154 454350 57774 471922
rect 57154 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 57774 454350
rect 57154 454226 57774 454294
rect 57154 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 57774 454226
rect 57154 454102 57774 454170
rect 57154 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 57774 454102
rect 57154 453978 57774 454046
rect 57154 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 57774 453978
rect 57154 436350 57774 453922
rect 57154 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436294 57774 436350
rect 57154 436226 57774 436294
rect 57154 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436170 57774 436226
rect 57154 436102 57774 436170
rect 57154 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436046 57774 436102
rect 57154 435978 57774 436046
rect 57154 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435922 57774 435978
rect 57154 418350 57774 435922
rect 57154 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 57774 418350
rect 57154 418226 57774 418294
rect 57154 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 57774 418226
rect 57154 418102 57774 418170
rect 57154 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 57774 418102
rect 57154 417978 57774 418046
rect 57154 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 57774 417978
rect 57154 400350 57774 417922
rect 57154 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 57774 400350
rect 57154 400226 57774 400294
rect 57154 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 57774 400226
rect 57154 400102 57774 400170
rect 57154 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 57774 400102
rect 57154 399978 57774 400046
rect 57154 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 57774 399978
rect 57154 382350 57774 399922
rect 57154 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 57774 382350
rect 57154 382226 57774 382294
rect 57154 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 57774 382226
rect 57154 382102 57774 382170
rect 57154 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 57774 382102
rect 57154 381978 57774 382046
rect 57154 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 57774 381978
rect 57154 364350 57774 381922
rect 57154 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 57774 364350
rect 57154 364226 57774 364294
rect 57154 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 57774 364226
rect 57154 364102 57774 364170
rect 57154 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 57774 364102
rect 57154 363978 57774 364046
rect 57154 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 57774 363978
rect 57154 346350 57774 363922
rect 57154 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 57774 346350
rect 57154 346226 57774 346294
rect 57154 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 57774 346226
rect 57154 346102 57774 346170
rect 57154 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 57774 346102
rect 57154 345978 57774 346046
rect 57154 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 57774 345978
rect 57154 328350 57774 345922
rect 57154 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 57774 328350
rect 57154 328226 57774 328294
rect 57154 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 57774 328226
rect 57154 328102 57774 328170
rect 57154 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 57774 328102
rect 57154 327978 57774 328046
rect 57154 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 57774 327978
rect 57154 310350 57774 327922
rect 57154 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 57774 310350
rect 57154 310226 57774 310294
rect 57154 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 57774 310226
rect 57154 310102 57774 310170
rect 57154 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 57774 310102
rect 57154 309978 57774 310046
rect 57154 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 57774 309978
rect 57154 292350 57774 309922
rect 57154 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 57774 292350
rect 57154 292226 57774 292294
rect 57154 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 57774 292226
rect 57154 292102 57774 292170
rect 57154 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 57774 292102
rect 57154 291978 57774 292046
rect 57154 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 57774 291978
rect 57154 274350 57774 291922
rect 57154 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 57774 274350
rect 57154 274226 57774 274294
rect 57154 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 57774 274226
rect 57154 274102 57774 274170
rect 57154 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 57774 274102
rect 57154 273978 57774 274046
rect 57154 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 57774 273978
rect 57154 256350 57774 273922
rect 57154 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 57774 256350
rect 57154 256226 57774 256294
rect 57154 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 57774 256226
rect 57154 256102 57774 256170
rect 57154 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 57774 256102
rect 57154 255978 57774 256046
rect 57154 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 57774 255978
rect 57154 238350 57774 255922
rect 57154 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 57774 238350
rect 57154 238226 57774 238294
rect 57154 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 57774 238226
rect 57154 238102 57774 238170
rect 57154 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 57774 238102
rect 57154 237978 57774 238046
rect 57154 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 57774 237978
rect 57154 220350 57774 237922
rect 57154 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 57774 220350
rect 57154 220226 57774 220294
rect 57154 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 57774 220226
rect 57154 220102 57774 220170
rect 57154 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 57774 220102
rect 57154 219978 57774 220046
rect 57154 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 57774 219978
rect 57154 202350 57774 219922
rect 57154 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 57774 202350
rect 57154 202226 57774 202294
rect 57154 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 57774 202226
rect 57154 202102 57774 202170
rect 57154 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 57774 202102
rect 57154 201978 57774 202046
rect 57154 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 57774 201978
rect 57154 184350 57774 201922
rect 57154 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 57774 184350
rect 57154 184226 57774 184294
rect 57154 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 57774 184226
rect 57154 184102 57774 184170
rect 57154 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 57774 184102
rect 57154 183978 57774 184046
rect 57154 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 57774 183978
rect 57154 166350 57774 183922
rect 57154 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 57774 166350
rect 57154 166226 57774 166294
rect 57154 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 57774 166226
rect 57154 166102 57774 166170
rect 57154 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 57774 166102
rect 57154 165978 57774 166046
rect 57154 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 57774 165978
rect 57154 148350 57774 165922
rect 57154 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 57774 148350
rect 57154 148226 57774 148294
rect 57154 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 57774 148226
rect 57154 148102 57774 148170
rect 57154 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 57774 148102
rect 57154 147978 57774 148046
rect 57154 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 57774 147978
rect 57154 130350 57774 147922
rect 57154 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 57774 130350
rect 57154 130226 57774 130294
rect 57154 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 57774 130226
rect 57154 130102 57774 130170
rect 57154 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 57774 130102
rect 57154 129978 57774 130046
rect 57154 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 57774 129978
rect 57154 112350 57774 129922
rect 57154 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 57774 112350
rect 57154 112226 57774 112294
rect 57154 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 57774 112226
rect 57154 112102 57774 112170
rect 57154 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 57774 112102
rect 57154 111978 57774 112046
rect 57154 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 57774 111978
rect 57154 94350 57774 111922
rect 57154 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 57774 94350
rect 57154 94226 57774 94294
rect 57154 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 57774 94226
rect 57154 94102 57774 94170
rect 57154 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 57774 94102
rect 57154 93978 57774 94046
rect 57154 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 57774 93978
rect 57154 76350 57774 93922
rect 57154 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 57774 76350
rect 57154 76226 57774 76294
rect 57154 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 57774 76226
rect 57154 76102 57774 76170
rect 57154 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 57774 76102
rect 57154 75978 57774 76046
rect 57154 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 57774 75978
rect 57154 58350 57774 75922
rect 57154 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 57774 58350
rect 57154 58226 57774 58294
rect 57154 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 57774 58226
rect 57154 58102 57774 58170
rect 57154 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 57774 58102
rect 57154 57978 57774 58046
rect 57154 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 57774 57978
rect 57154 40350 57774 57922
rect 57154 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 57774 40350
rect 57154 40226 57774 40294
rect 57154 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 57774 40226
rect 57154 40102 57774 40170
rect 57154 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 57774 40102
rect 57154 39978 57774 40046
rect 57154 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 57774 39978
rect 57154 22350 57774 39922
rect 57154 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 57774 22350
rect 57154 22226 57774 22294
rect 57154 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 57774 22226
rect 57154 22102 57774 22170
rect 57154 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 57774 22102
rect 57154 21978 57774 22046
rect 57154 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 57774 21978
rect 57154 4350 57774 21922
rect 57154 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 57774 4350
rect 57154 4226 57774 4294
rect 57154 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 57774 4226
rect 57154 4102 57774 4170
rect 57154 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 57774 4102
rect 57154 3978 57774 4046
rect 57154 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 57774 3978
rect 57154 -160 57774 3922
rect 57154 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 57774 -160
rect 57154 -284 57774 -216
rect 57154 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 57774 -284
rect 57154 -408 57774 -340
rect 57154 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 57774 -408
rect 57154 -532 57774 -464
rect 57154 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 57774 -532
rect 57154 -1644 57774 -588
rect 60874 598172 61494 598268
rect 60874 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 61494 598172
rect 60874 598048 61494 598116
rect 60874 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 61494 598048
rect 60874 597924 61494 597992
rect 60874 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 61494 597924
rect 60874 597800 61494 597868
rect 60874 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 61494 597800
rect 60874 586350 61494 597744
rect 60874 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 61494 586350
rect 60874 586226 61494 586294
rect 60874 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 61494 586226
rect 60874 586102 61494 586170
rect 60874 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 61494 586102
rect 60874 585978 61494 586046
rect 60874 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 61494 585978
rect 60874 568350 61494 585922
rect 60874 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 61494 568350
rect 60874 568226 61494 568294
rect 60874 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 61494 568226
rect 60874 568102 61494 568170
rect 60874 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 61494 568102
rect 60874 567978 61494 568046
rect 60874 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 61494 567978
rect 60874 550350 61494 567922
rect 60874 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 61494 550350
rect 60874 550226 61494 550294
rect 60874 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 61494 550226
rect 60874 550102 61494 550170
rect 60874 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 61494 550102
rect 60874 549978 61494 550046
rect 60874 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 61494 549978
rect 60874 532350 61494 549922
rect 60874 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 61494 532350
rect 60874 532226 61494 532294
rect 60874 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 61494 532226
rect 60874 532102 61494 532170
rect 60874 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 61494 532102
rect 60874 531978 61494 532046
rect 60874 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 61494 531978
rect 60874 514350 61494 531922
rect 60874 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 61494 514350
rect 60874 514226 61494 514294
rect 60874 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 61494 514226
rect 60874 514102 61494 514170
rect 60874 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 61494 514102
rect 60874 513978 61494 514046
rect 60874 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 61494 513978
rect 60874 496350 61494 513922
rect 60874 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 61494 496350
rect 60874 496226 61494 496294
rect 60874 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 61494 496226
rect 60874 496102 61494 496170
rect 60874 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 61494 496102
rect 60874 495978 61494 496046
rect 60874 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 61494 495978
rect 60874 478350 61494 495922
rect 60874 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 61494 478350
rect 60874 478226 61494 478294
rect 60874 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 61494 478226
rect 60874 478102 61494 478170
rect 60874 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 61494 478102
rect 60874 477978 61494 478046
rect 60874 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 61494 477978
rect 60874 460350 61494 477922
rect 60874 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 61494 460350
rect 60874 460226 61494 460294
rect 60874 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 61494 460226
rect 60874 460102 61494 460170
rect 60874 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 61494 460102
rect 60874 459978 61494 460046
rect 60874 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 61494 459978
rect 60874 442350 61494 459922
rect 60874 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 61494 442350
rect 60874 442226 61494 442294
rect 60874 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 61494 442226
rect 60874 442102 61494 442170
rect 60874 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 61494 442102
rect 60874 441978 61494 442046
rect 60874 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 61494 441978
rect 60874 424350 61494 441922
rect 60874 424294 60970 424350
rect 61026 424294 61094 424350
rect 61150 424294 61218 424350
rect 61274 424294 61342 424350
rect 61398 424294 61494 424350
rect 60874 424226 61494 424294
rect 60874 424170 60970 424226
rect 61026 424170 61094 424226
rect 61150 424170 61218 424226
rect 61274 424170 61342 424226
rect 61398 424170 61494 424226
rect 60874 424102 61494 424170
rect 60874 424046 60970 424102
rect 61026 424046 61094 424102
rect 61150 424046 61218 424102
rect 61274 424046 61342 424102
rect 61398 424046 61494 424102
rect 60874 423978 61494 424046
rect 60874 423922 60970 423978
rect 61026 423922 61094 423978
rect 61150 423922 61218 423978
rect 61274 423922 61342 423978
rect 61398 423922 61494 423978
rect 60874 406350 61494 423922
rect 60874 406294 60970 406350
rect 61026 406294 61094 406350
rect 61150 406294 61218 406350
rect 61274 406294 61342 406350
rect 61398 406294 61494 406350
rect 60874 406226 61494 406294
rect 60874 406170 60970 406226
rect 61026 406170 61094 406226
rect 61150 406170 61218 406226
rect 61274 406170 61342 406226
rect 61398 406170 61494 406226
rect 60874 406102 61494 406170
rect 60874 406046 60970 406102
rect 61026 406046 61094 406102
rect 61150 406046 61218 406102
rect 61274 406046 61342 406102
rect 61398 406046 61494 406102
rect 60874 405978 61494 406046
rect 60874 405922 60970 405978
rect 61026 405922 61094 405978
rect 61150 405922 61218 405978
rect 61274 405922 61342 405978
rect 61398 405922 61494 405978
rect 60874 388350 61494 405922
rect 60874 388294 60970 388350
rect 61026 388294 61094 388350
rect 61150 388294 61218 388350
rect 61274 388294 61342 388350
rect 61398 388294 61494 388350
rect 60874 388226 61494 388294
rect 60874 388170 60970 388226
rect 61026 388170 61094 388226
rect 61150 388170 61218 388226
rect 61274 388170 61342 388226
rect 61398 388170 61494 388226
rect 60874 388102 61494 388170
rect 60874 388046 60970 388102
rect 61026 388046 61094 388102
rect 61150 388046 61218 388102
rect 61274 388046 61342 388102
rect 61398 388046 61494 388102
rect 60874 387978 61494 388046
rect 60874 387922 60970 387978
rect 61026 387922 61094 387978
rect 61150 387922 61218 387978
rect 61274 387922 61342 387978
rect 61398 387922 61494 387978
rect 60874 370350 61494 387922
rect 60874 370294 60970 370350
rect 61026 370294 61094 370350
rect 61150 370294 61218 370350
rect 61274 370294 61342 370350
rect 61398 370294 61494 370350
rect 60874 370226 61494 370294
rect 60874 370170 60970 370226
rect 61026 370170 61094 370226
rect 61150 370170 61218 370226
rect 61274 370170 61342 370226
rect 61398 370170 61494 370226
rect 60874 370102 61494 370170
rect 60874 370046 60970 370102
rect 61026 370046 61094 370102
rect 61150 370046 61218 370102
rect 61274 370046 61342 370102
rect 61398 370046 61494 370102
rect 60874 369978 61494 370046
rect 60874 369922 60970 369978
rect 61026 369922 61094 369978
rect 61150 369922 61218 369978
rect 61274 369922 61342 369978
rect 61398 369922 61494 369978
rect 60874 352350 61494 369922
rect 60874 352294 60970 352350
rect 61026 352294 61094 352350
rect 61150 352294 61218 352350
rect 61274 352294 61342 352350
rect 61398 352294 61494 352350
rect 60874 352226 61494 352294
rect 60874 352170 60970 352226
rect 61026 352170 61094 352226
rect 61150 352170 61218 352226
rect 61274 352170 61342 352226
rect 61398 352170 61494 352226
rect 60874 352102 61494 352170
rect 60874 352046 60970 352102
rect 61026 352046 61094 352102
rect 61150 352046 61218 352102
rect 61274 352046 61342 352102
rect 61398 352046 61494 352102
rect 60874 351978 61494 352046
rect 60874 351922 60970 351978
rect 61026 351922 61094 351978
rect 61150 351922 61218 351978
rect 61274 351922 61342 351978
rect 61398 351922 61494 351978
rect 60874 334350 61494 351922
rect 60874 334294 60970 334350
rect 61026 334294 61094 334350
rect 61150 334294 61218 334350
rect 61274 334294 61342 334350
rect 61398 334294 61494 334350
rect 60874 334226 61494 334294
rect 60874 334170 60970 334226
rect 61026 334170 61094 334226
rect 61150 334170 61218 334226
rect 61274 334170 61342 334226
rect 61398 334170 61494 334226
rect 60874 334102 61494 334170
rect 60874 334046 60970 334102
rect 61026 334046 61094 334102
rect 61150 334046 61218 334102
rect 61274 334046 61342 334102
rect 61398 334046 61494 334102
rect 60874 333978 61494 334046
rect 60874 333922 60970 333978
rect 61026 333922 61094 333978
rect 61150 333922 61218 333978
rect 61274 333922 61342 333978
rect 61398 333922 61494 333978
rect 60874 316350 61494 333922
rect 60874 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 61494 316350
rect 60874 316226 61494 316294
rect 60874 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 61494 316226
rect 60874 316102 61494 316170
rect 60874 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 61494 316102
rect 60874 315978 61494 316046
rect 60874 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 61494 315978
rect 60874 298350 61494 315922
rect 60874 298294 60970 298350
rect 61026 298294 61094 298350
rect 61150 298294 61218 298350
rect 61274 298294 61342 298350
rect 61398 298294 61494 298350
rect 60874 298226 61494 298294
rect 60874 298170 60970 298226
rect 61026 298170 61094 298226
rect 61150 298170 61218 298226
rect 61274 298170 61342 298226
rect 61398 298170 61494 298226
rect 60874 298102 61494 298170
rect 60874 298046 60970 298102
rect 61026 298046 61094 298102
rect 61150 298046 61218 298102
rect 61274 298046 61342 298102
rect 61398 298046 61494 298102
rect 60874 297978 61494 298046
rect 60874 297922 60970 297978
rect 61026 297922 61094 297978
rect 61150 297922 61218 297978
rect 61274 297922 61342 297978
rect 61398 297922 61494 297978
rect 60874 280350 61494 297922
rect 60874 280294 60970 280350
rect 61026 280294 61094 280350
rect 61150 280294 61218 280350
rect 61274 280294 61342 280350
rect 61398 280294 61494 280350
rect 60874 280226 61494 280294
rect 60874 280170 60970 280226
rect 61026 280170 61094 280226
rect 61150 280170 61218 280226
rect 61274 280170 61342 280226
rect 61398 280170 61494 280226
rect 60874 280102 61494 280170
rect 60874 280046 60970 280102
rect 61026 280046 61094 280102
rect 61150 280046 61218 280102
rect 61274 280046 61342 280102
rect 61398 280046 61494 280102
rect 60874 279978 61494 280046
rect 60874 279922 60970 279978
rect 61026 279922 61094 279978
rect 61150 279922 61218 279978
rect 61274 279922 61342 279978
rect 61398 279922 61494 279978
rect 60874 262350 61494 279922
rect 60874 262294 60970 262350
rect 61026 262294 61094 262350
rect 61150 262294 61218 262350
rect 61274 262294 61342 262350
rect 61398 262294 61494 262350
rect 60874 262226 61494 262294
rect 60874 262170 60970 262226
rect 61026 262170 61094 262226
rect 61150 262170 61218 262226
rect 61274 262170 61342 262226
rect 61398 262170 61494 262226
rect 60874 262102 61494 262170
rect 60874 262046 60970 262102
rect 61026 262046 61094 262102
rect 61150 262046 61218 262102
rect 61274 262046 61342 262102
rect 61398 262046 61494 262102
rect 60874 261978 61494 262046
rect 60874 261922 60970 261978
rect 61026 261922 61094 261978
rect 61150 261922 61218 261978
rect 61274 261922 61342 261978
rect 61398 261922 61494 261978
rect 60874 244350 61494 261922
rect 60874 244294 60970 244350
rect 61026 244294 61094 244350
rect 61150 244294 61218 244350
rect 61274 244294 61342 244350
rect 61398 244294 61494 244350
rect 60874 244226 61494 244294
rect 60874 244170 60970 244226
rect 61026 244170 61094 244226
rect 61150 244170 61218 244226
rect 61274 244170 61342 244226
rect 61398 244170 61494 244226
rect 60874 244102 61494 244170
rect 60874 244046 60970 244102
rect 61026 244046 61094 244102
rect 61150 244046 61218 244102
rect 61274 244046 61342 244102
rect 61398 244046 61494 244102
rect 60874 243978 61494 244046
rect 60874 243922 60970 243978
rect 61026 243922 61094 243978
rect 61150 243922 61218 243978
rect 61274 243922 61342 243978
rect 61398 243922 61494 243978
rect 60874 226350 61494 243922
rect 60874 226294 60970 226350
rect 61026 226294 61094 226350
rect 61150 226294 61218 226350
rect 61274 226294 61342 226350
rect 61398 226294 61494 226350
rect 60874 226226 61494 226294
rect 60874 226170 60970 226226
rect 61026 226170 61094 226226
rect 61150 226170 61218 226226
rect 61274 226170 61342 226226
rect 61398 226170 61494 226226
rect 60874 226102 61494 226170
rect 60874 226046 60970 226102
rect 61026 226046 61094 226102
rect 61150 226046 61218 226102
rect 61274 226046 61342 226102
rect 61398 226046 61494 226102
rect 60874 225978 61494 226046
rect 60874 225922 60970 225978
rect 61026 225922 61094 225978
rect 61150 225922 61218 225978
rect 61274 225922 61342 225978
rect 61398 225922 61494 225978
rect 60874 208350 61494 225922
rect 60874 208294 60970 208350
rect 61026 208294 61094 208350
rect 61150 208294 61218 208350
rect 61274 208294 61342 208350
rect 61398 208294 61494 208350
rect 60874 208226 61494 208294
rect 60874 208170 60970 208226
rect 61026 208170 61094 208226
rect 61150 208170 61218 208226
rect 61274 208170 61342 208226
rect 61398 208170 61494 208226
rect 60874 208102 61494 208170
rect 60874 208046 60970 208102
rect 61026 208046 61094 208102
rect 61150 208046 61218 208102
rect 61274 208046 61342 208102
rect 61398 208046 61494 208102
rect 60874 207978 61494 208046
rect 60874 207922 60970 207978
rect 61026 207922 61094 207978
rect 61150 207922 61218 207978
rect 61274 207922 61342 207978
rect 61398 207922 61494 207978
rect 60874 190350 61494 207922
rect 60874 190294 60970 190350
rect 61026 190294 61094 190350
rect 61150 190294 61218 190350
rect 61274 190294 61342 190350
rect 61398 190294 61494 190350
rect 60874 190226 61494 190294
rect 60874 190170 60970 190226
rect 61026 190170 61094 190226
rect 61150 190170 61218 190226
rect 61274 190170 61342 190226
rect 61398 190170 61494 190226
rect 60874 190102 61494 190170
rect 60874 190046 60970 190102
rect 61026 190046 61094 190102
rect 61150 190046 61218 190102
rect 61274 190046 61342 190102
rect 61398 190046 61494 190102
rect 60874 189978 61494 190046
rect 60874 189922 60970 189978
rect 61026 189922 61094 189978
rect 61150 189922 61218 189978
rect 61274 189922 61342 189978
rect 61398 189922 61494 189978
rect 60874 172350 61494 189922
rect 60874 172294 60970 172350
rect 61026 172294 61094 172350
rect 61150 172294 61218 172350
rect 61274 172294 61342 172350
rect 61398 172294 61494 172350
rect 60874 172226 61494 172294
rect 60874 172170 60970 172226
rect 61026 172170 61094 172226
rect 61150 172170 61218 172226
rect 61274 172170 61342 172226
rect 61398 172170 61494 172226
rect 60874 172102 61494 172170
rect 60874 172046 60970 172102
rect 61026 172046 61094 172102
rect 61150 172046 61218 172102
rect 61274 172046 61342 172102
rect 61398 172046 61494 172102
rect 60874 171978 61494 172046
rect 60874 171922 60970 171978
rect 61026 171922 61094 171978
rect 61150 171922 61218 171978
rect 61274 171922 61342 171978
rect 61398 171922 61494 171978
rect 60874 154350 61494 171922
rect 60874 154294 60970 154350
rect 61026 154294 61094 154350
rect 61150 154294 61218 154350
rect 61274 154294 61342 154350
rect 61398 154294 61494 154350
rect 60874 154226 61494 154294
rect 60874 154170 60970 154226
rect 61026 154170 61094 154226
rect 61150 154170 61218 154226
rect 61274 154170 61342 154226
rect 61398 154170 61494 154226
rect 60874 154102 61494 154170
rect 60874 154046 60970 154102
rect 61026 154046 61094 154102
rect 61150 154046 61218 154102
rect 61274 154046 61342 154102
rect 61398 154046 61494 154102
rect 60874 153978 61494 154046
rect 60874 153922 60970 153978
rect 61026 153922 61094 153978
rect 61150 153922 61218 153978
rect 61274 153922 61342 153978
rect 61398 153922 61494 153978
rect 60874 136350 61494 153922
rect 60874 136294 60970 136350
rect 61026 136294 61094 136350
rect 61150 136294 61218 136350
rect 61274 136294 61342 136350
rect 61398 136294 61494 136350
rect 60874 136226 61494 136294
rect 60874 136170 60970 136226
rect 61026 136170 61094 136226
rect 61150 136170 61218 136226
rect 61274 136170 61342 136226
rect 61398 136170 61494 136226
rect 60874 136102 61494 136170
rect 60874 136046 60970 136102
rect 61026 136046 61094 136102
rect 61150 136046 61218 136102
rect 61274 136046 61342 136102
rect 61398 136046 61494 136102
rect 60874 135978 61494 136046
rect 60874 135922 60970 135978
rect 61026 135922 61094 135978
rect 61150 135922 61218 135978
rect 61274 135922 61342 135978
rect 61398 135922 61494 135978
rect 60874 118350 61494 135922
rect 60874 118294 60970 118350
rect 61026 118294 61094 118350
rect 61150 118294 61218 118350
rect 61274 118294 61342 118350
rect 61398 118294 61494 118350
rect 60874 118226 61494 118294
rect 60874 118170 60970 118226
rect 61026 118170 61094 118226
rect 61150 118170 61218 118226
rect 61274 118170 61342 118226
rect 61398 118170 61494 118226
rect 60874 118102 61494 118170
rect 60874 118046 60970 118102
rect 61026 118046 61094 118102
rect 61150 118046 61218 118102
rect 61274 118046 61342 118102
rect 61398 118046 61494 118102
rect 60874 117978 61494 118046
rect 60874 117922 60970 117978
rect 61026 117922 61094 117978
rect 61150 117922 61218 117978
rect 61274 117922 61342 117978
rect 61398 117922 61494 117978
rect 60874 100350 61494 117922
rect 60874 100294 60970 100350
rect 61026 100294 61094 100350
rect 61150 100294 61218 100350
rect 61274 100294 61342 100350
rect 61398 100294 61494 100350
rect 60874 100226 61494 100294
rect 60874 100170 60970 100226
rect 61026 100170 61094 100226
rect 61150 100170 61218 100226
rect 61274 100170 61342 100226
rect 61398 100170 61494 100226
rect 60874 100102 61494 100170
rect 60874 100046 60970 100102
rect 61026 100046 61094 100102
rect 61150 100046 61218 100102
rect 61274 100046 61342 100102
rect 61398 100046 61494 100102
rect 60874 99978 61494 100046
rect 60874 99922 60970 99978
rect 61026 99922 61094 99978
rect 61150 99922 61218 99978
rect 61274 99922 61342 99978
rect 61398 99922 61494 99978
rect 60874 82350 61494 99922
rect 60874 82294 60970 82350
rect 61026 82294 61094 82350
rect 61150 82294 61218 82350
rect 61274 82294 61342 82350
rect 61398 82294 61494 82350
rect 60874 82226 61494 82294
rect 60874 82170 60970 82226
rect 61026 82170 61094 82226
rect 61150 82170 61218 82226
rect 61274 82170 61342 82226
rect 61398 82170 61494 82226
rect 60874 82102 61494 82170
rect 60874 82046 60970 82102
rect 61026 82046 61094 82102
rect 61150 82046 61218 82102
rect 61274 82046 61342 82102
rect 61398 82046 61494 82102
rect 60874 81978 61494 82046
rect 60874 81922 60970 81978
rect 61026 81922 61094 81978
rect 61150 81922 61218 81978
rect 61274 81922 61342 81978
rect 61398 81922 61494 81978
rect 60874 64350 61494 81922
rect 60874 64294 60970 64350
rect 61026 64294 61094 64350
rect 61150 64294 61218 64350
rect 61274 64294 61342 64350
rect 61398 64294 61494 64350
rect 60874 64226 61494 64294
rect 60874 64170 60970 64226
rect 61026 64170 61094 64226
rect 61150 64170 61218 64226
rect 61274 64170 61342 64226
rect 61398 64170 61494 64226
rect 60874 64102 61494 64170
rect 60874 64046 60970 64102
rect 61026 64046 61094 64102
rect 61150 64046 61218 64102
rect 61274 64046 61342 64102
rect 61398 64046 61494 64102
rect 60874 63978 61494 64046
rect 60874 63922 60970 63978
rect 61026 63922 61094 63978
rect 61150 63922 61218 63978
rect 61274 63922 61342 63978
rect 61398 63922 61494 63978
rect 60874 46350 61494 63922
rect 60874 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 61494 46350
rect 60874 46226 61494 46294
rect 60874 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 61494 46226
rect 60874 46102 61494 46170
rect 60874 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 61494 46102
rect 60874 45978 61494 46046
rect 60874 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 61494 45978
rect 60874 28350 61494 45922
rect 60874 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 61494 28350
rect 60874 28226 61494 28294
rect 60874 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 61494 28226
rect 60874 28102 61494 28170
rect 60874 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 61494 28102
rect 60874 27978 61494 28046
rect 60874 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 61494 27978
rect 60874 10350 61494 27922
rect 60874 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 61494 10350
rect 60874 10226 61494 10294
rect 60874 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 61494 10226
rect 60874 10102 61494 10170
rect 60874 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 61494 10102
rect 60874 9978 61494 10046
rect 60874 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 61494 9978
rect 60874 -1120 61494 9922
rect 60874 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 61494 -1120
rect 60874 -1244 61494 -1176
rect 60874 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 61494 -1244
rect 60874 -1368 61494 -1300
rect 60874 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 61494 -1368
rect 60874 -1492 61494 -1424
rect 60874 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 61494 -1492
rect 60874 -1644 61494 -1548
rect 75154 597212 75774 598268
rect 75154 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 75774 597212
rect 75154 597088 75774 597156
rect 75154 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 75774 597088
rect 75154 596964 75774 597032
rect 75154 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 75774 596964
rect 75154 596840 75774 596908
rect 75154 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 75774 596840
rect 75154 580350 75774 596784
rect 75154 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 75774 580350
rect 75154 580226 75774 580294
rect 75154 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 75774 580226
rect 75154 580102 75774 580170
rect 75154 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 75774 580102
rect 75154 579978 75774 580046
rect 75154 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 75774 579978
rect 75154 562350 75774 579922
rect 75154 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 75774 562350
rect 75154 562226 75774 562294
rect 75154 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 75774 562226
rect 75154 562102 75774 562170
rect 75154 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 75774 562102
rect 75154 561978 75774 562046
rect 75154 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 75774 561978
rect 75154 544350 75774 561922
rect 75154 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 75774 544350
rect 75154 544226 75774 544294
rect 75154 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 75774 544226
rect 75154 544102 75774 544170
rect 75154 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 75774 544102
rect 75154 543978 75774 544046
rect 75154 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 75774 543978
rect 75154 526350 75774 543922
rect 75154 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 75774 526350
rect 75154 526226 75774 526294
rect 75154 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 75774 526226
rect 75154 526102 75774 526170
rect 75154 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 75774 526102
rect 75154 525978 75774 526046
rect 75154 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 75774 525978
rect 75154 508350 75774 525922
rect 75154 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 75774 508350
rect 75154 508226 75774 508294
rect 75154 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 75774 508226
rect 75154 508102 75774 508170
rect 75154 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 75774 508102
rect 75154 507978 75774 508046
rect 75154 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 75774 507978
rect 75154 490350 75774 507922
rect 75154 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 75774 490350
rect 75154 490226 75774 490294
rect 75154 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 75774 490226
rect 75154 490102 75774 490170
rect 75154 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 75774 490102
rect 75154 489978 75774 490046
rect 75154 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 75774 489978
rect 75154 472350 75774 489922
rect 75154 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 75774 472350
rect 75154 472226 75774 472294
rect 75154 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 75774 472226
rect 75154 472102 75774 472170
rect 75154 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 75774 472102
rect 75154 471978 75774 472046
rect 75154 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 75774 471978
rect 75154 454350 75774 471922
rect 75154 454294 75250 454350
rect 75306 454294 75374 454350
rect 75430 454294 75498 454350
rect 75554 454294 75622 454350
rect 75678 454294 75774 454350
rect 75154 454226 75774 454294
rect 75154 454170 75250 454226
rect 75306 454170 75374 454226
rect 75430 454170 75498 454226
rect 75554 454170 75622 454226
rect 75678 454170 75774 454226
rect 75154 454102 75774 454170
rect 75154 454046 75250 454102
rect 75306 454046 75374 454102
rect 75430 454046 75498 454102
rect 75554 454046 75622 454102
rect 75678 454046 75774 454102
rect 75154 453978 75774 454046
rect 75154 453922 75250 453978
rect 75306 453922 75374 453978
rect 75430 453922 75498 453978
rect 75554 453922 75622 453978
rect 75678 453922 75774 453978
rect 75154 436350 75774 453922
rect 75154 436294 75250 436350
rect 75306 436294 75374 436350
rect 75430 436294 75498 436350
rect 75554 436294 75622 436350
rect 75678 436294 75774 436350
rect 75154 436226 75774 436294
rect 75154 436170 75250 436226
rect 75306 436170 75374 436226
rect 75430 436170 75498 436226
rect 75554 436170 75622 436226
rect 75678 436170 75774 436226
rect 75154 436102 75774 436170
rect 75154 436046 75250 436102
rect 75306 436046 75374 436102
rect 75430 436046 75498 436102
rect 75554 436046 75622 436102
rect 75678 436046 75774 436102
rect 75154 435978 75774 436046
rect 75154 435922 75250 435978
rect 75306 435922 75374 435978
rect 75430 435922 75498 435978
rect 75554 435922 75622 435978
rect 75678 435922 75774 435978
rect 75154 418350 75774 435922
rect 75154 418294 75250 418350
rect 75306 418294 75374 418350
rect 75430 418294 75498 418350
rect 75554 418294 75622 418350
rect 75678 418294 75774 418350
rect 75154 418226 75774 418294
rect 75154 418170 75250 418226
rect 75306 418170 75374 418226
rect 75430 418170 75498 418226
rect 75554 418170 75622 418226
rect 75678 418170 75774 418226
rect 75154 418102 75774 418170
rect 75154 418046 75250 418102
rect 75306 418046 75374 418102
rect 75430 418046 75498 418102
rect 75554 418046 75622 418102
rect 75678 418046 75774 418102
rect 75154 417978 75774 418046
rect 75154 417922 75250 417978
rect 75306 417922 75374 417978
rect 75430 417922 75498 417978
rect 75554 417922 75622 417978
rect 75678 417922 75774 417978
rect 75154 400350 75774 417922
rect 75154 400294 75250 400350
rect 75306 400294 75374 400350
rect 75430 400294 75498 400350
rect 75554 400294 75622 400350
rect 75678 400294 75774 400350
rect 75154 400226 75774 400294
rect 75154 400170 75250 400226
rect 75306 400170 75374 400226
rect 75430 400170 75498 400226
rect 75554 400170 75622 400226
rect 75678 400170 75774 400226
rect 75154 400102 75774 400170
rect 75154 400046 75250 400102
rect 75306 400046 75374 400102
rect 75430 400046 75498 400102
rect 75554 400046 75622 400102
rect 75678 400046 75774 400102
rect 75154 399978 75774 400046
rect 75154 399922 75250 399978
rect 75306 399922 75374 399978
rect 75430 399922 75498 399978
rect 75554 399922 75622 399978
rect 75678 399922 75774 399978
rect 75154 382350 75774 399922
rect 75154 382294 75250 382350
rect 75306 382294 75374 382350
rect 75430 382294 75498 382350
rect 75554 382294 75622 382350
rect 75678 382294 75774 382350
rect 75154 382226 75774 382294
rect 75154 382170 75250 382226
rect 75306 382170 75374 382226
rect 75430 382170 75498 382226
rect 75554 382170 75622 382226
rect 75678 382170 75774 382226
rect 75154 382102 75774 382170
rect 75154 382046 75250 382102
rect 75306 382046 75374 382102
rect 75430 382046 75498 382102
rect 75554 382046 75622 382102
rect 75678 382046 75774 382102
rect 75154 381978 75774 382046
rect 75154 381922 75250 381978
rect 75306 381922 75374 381978
rect 75430 381922 75498 381978
rect 75554 381922 75622 381978
rect 75678 381922 75774 381978
rect 75154 364350 75774 381922
rect 75154 364294 75250 364350
rect 75306 364294 75374 364350
rect 75430 364294 75498 364350
rect 75554 364294 75622 364350
rect 75678 364294 75774 364350
rect 75154 364226 75774 364294
rect 75154 364170 75250 364226
rect 75306 364170 75374 364226
rect 75430 364170 75498 364226
rect 75554 364170 75622 364226
rect 75678 364170 75774 364226
rect 75154 364102 75774 364170
rect 75154 364046 75250 364102
rect 75306 364046 75374 364102
rect 75430 364046 75498 364102
rect 75554 364046 75622 364102
rect 75678 364046 75774 364102
rect 75154 363978 75774 364046
rect 75154 363922 75250 363978
rect 75306 363922 75374 363978
rect 75430 363922 75498 363978
rect 75554 363922 75622 363978
rect 75678 363922 75774 363978
rect 75154 346350 75774 363922
rect 75154 346294 75250 346350
rect 75306 346294 75374 346350
rect 75430 346294 75498 346350
rect 75554 346294 75622 346350
rect 75678 346294 75774 346350
rect 75154 346226 75774 346294
rect 75154 346170 75250 346226
rect 75306 346170 75374 346226
rect 75430 346170 75498 346226
rect 75554 346170 75622 346226
rect 75678 346170 75774 346226
rect 75154 346102 75774 346170
rect 75154 346046 75250 346102
rect 75306 346046 75374 346102
rect 75430 346046 75498 346102
rect 75554 346046 75622 346102
rect 75678 346046 75774 346102
rect 75154 345978 75774 346046
rect 75154 345922 75250 345978
rect 75306 345922 75374 345978
rect 75430 345922 75498 345978
rect 75554 345922 75622 345978
rect 75678 345922 75774 345978
rect 75154 328350 75774 345922
rect 75154 328294 75250 328350
rect 75306 328294 75374 328350
rect 75430 328294 75498 328350
rect 75554 328294 75622 328350
rect 75678 328294 75774 328350
rect 75154 328226 75774 328294
rect 75154 328170 75250 328226
rect 75306 328170 75374 328226
rect 75430 328170 75498 328226
rect 75554 328170 75622 328226
rect 75678 328170 75774 328226
rect 75154 328102 75774 328170
rect 75154 328046 75250 328102
rect 75306 328046 75374 328102
rect 75430 328046 75498 328102
rect 75554 328046 75622 328102
rect 75678 328046 75774 328102
rect 75154 327978 75774 328046
rect 75154 327922 75250 327978
rect 75306 327922 75374 327978
rect 75430 327922 75498 327978
rect 75554 327922 75622 327978
rect 75678 327922 75774 327978
rect 75154 310350 75774 327922
rect 75154 310294 75250 310350
rect 75306 310294 75374 310350
rect 75430 310294 75498 310350
rect 75554 310294 75622 310350
rect 75678 310294 75774 310350
rect 75154 310226 75774 310294
rect 75154 310170 75250 310226
rect 75306 310170 75374 310226
rect 75430 310170 75498 310226
rect 75554 310170 75622 310226
rect 75678 310170 75774 310226
rect 75154 310102 75774 310170
rect 75154 310046 75250 310102
rect 75306 310046 75374 310102
rect 75430 310046 75498 310102
rect 75554 310046 75622 310102
rect 75678 310046 75774 310102
rect 75154 309978 75774 310046
rect 75154 309922 75250 309978
rect 75306 309922 75374 309978
rect 75430 309922 75498 309978
rect 75554 309922 75622 309978
rect 75678 309922 75774 309978
rect 75154 292350 75774 309922
rect 75154 292294 75250 292350
rect 75306 292294 75374 292350
rect 75430 292294 75498 292350
rect 75554 292294 75622 292350
rect 75678 292294 75774 292350
rect 75154 292226 75774 292294
rect 75154 292170 75250 292226
rect 75306 292170 75374 292226
rect 75430 292170 75498 292226
rect 75554 292170 75622 292226
rect 75678 292170 75774 292226
rect 75154 292102 75774 292170
rect 75154 292046 75250 292102
rect 75306 292046 75374 292102
rect 75430 292046 75498 292102
rect 75554 292046 75622 292102
rect 75678 292046 75774 292102
rect 75154 291978 75774 292046
rect 75154 291922 75250 291978
rect 75306 291922 75374 291978
rect 75430 291922 75498 291978
rect 75554 291922 75622 291978
rect 75678 291922 75774 291978
rect 75154 274350 75774 291922
rect 75154 274294 75250 274350
rect 75306 274294 75374 274350
rect 75430 274294 75498 274350
rect 75554 274294 75622 274350
rect 75678 274294 75774 274350
rect 75154 274226 75774 274294
rect 75154 274170 75250 274226
rect 75306 274170 75374 274226
rect 75430 274170 75498 274226
rect 75554 274170 75622 274226
rect 75678 274170 75774 274226
rect 75154 274102 75774 274170
rect 75154 274046 75250 274102
rect 75306 274046 75374 274102
rect 75430 274046 75498 274102
rect 75554 274046 75622 274102
rect 75678 274046 75774 274102
rect 75154 273978 75774 274046
rect 75154 273922 75250 273978
rect 75306 273922 75374 273978
rect 75430 273922 75498 273978
rect 75554 273922 75622 273978
rect 75678 273922 75774 273978
rect 75154 256350 75774 273922
rect 75154 256294 75250 256350
rect 75306 256294 75374 256350
rect 75430 256294 75498 256350
rect 75554 256294 75622 256350
rect 75678 256294 75774 256350
rect 75154 256226 75774 256294
rect 75154 256170 75250 256226
rect 75306 256170 75374 256226
rect 75430 256170 75498 256226
rect 75554 256170 75622 256226
rect 75678 256170 75774 256226
rect 75154 256102 75774 256170
rect 75154 256046 75250 256102
rect 75306 256046 75374 256102
rect 75430 256046 75498 256102
rect 75554 256046 75622 256102
rect 75678 256046 75774 256102
rect 75154 255978 75774 256046
rect 75154 255922 75250 255978
rect 75306 255922 75374 255978
rect 75430 255922 75498 255978
rect 75554 255922 75622 255978
rect 75678 255922 75774 255978
rect 75154 238350 75774 255922
rect 75154 238294 75250 238350
rect 75306 238294 75374 238350
rect 75430 238294 75498 238350
rect 75554 238294 75622 238350
rect 75678 238294 75774 238350
rect 75154 238226 75774 238294
rect 75154 238170 75250 238226
rect 75306 238170 75374 238226
rect 75430 238170 75498 238226
rect 75554 238170 75622 238226
rect 75678 238170 75774 238226
rect 75154 238102 75774 238170
rect 75154 238046 75250 238102
rect 75306 238046 75374 238102
rect 75430 238046 75498 238102
rect 75554 238046 75622 238102
rect 75678 238046 75774 238102
rect 75154 237978 75774 238046
rect 75154 237922 75250 237978
rect 75306 237922 75374 237978
rect 75430 237922 75498 237978
rect 75554 237922 75622 237978
rect 75678 237922 75774 237978
rect 75154 220350 75774 237922
rect 75154 220294 75250 220350
rect 75306 220294 75374 220350
rect 75430 220294 75498 220350
rect 75554 220294 75622 220350
rect 75678 220294 75774 220350
rect 75154 220226 75774 220294
rect 75154 220170 75250 220226
rect 75306 220170 75374 220226
rect 75430 220170 75498 220226
rect 75554 220170 75622 220226
rect 75678 220170 75774 220226
rect 75154 220102 75774 220170
rect 75154 220046 75250 220102
rect 75306 220046 75374 220102
rect 75430 220046 75498 220102
rect 75554 220046 75622 220102
rect 75678 220046 75774 220102
rect 75154 219978 75774 220046
rect 75154 219922 75250 219978
rect 75306 219922 75374 219978
rect 75430 219922 75498 219978
rect 75554 219922 75622 219978
rect 75678 219922 75774 219978
rect 75154 202350 75774 219922
rect 75154 202294 75250 202350
rect 75306 202294 75374 202350
rect 75430 202294 75498 202350
rect 75554 202294 75622 202350
rect 75678 202294 75774 202350
rect 75154 202226 75774 202294
rect 75154 202170 75250 202226
rect 75306 202170 75374 202226
rect 75430 202170 75498 202226
rect 75554 202170 75622 202226
rect 75678 202170 75774 202226
rect 75154 202102 75774 202170
rect 75154 202046 75250 202102
rect 75306 202046 75374 202102
rect 75430 202046 75498 202102
rect 75554 202046 75622 202102
rect 75678 202046 75774 202102
rect 75154 201978 75774 202046
rect 75154 201922 75250 201978
rect 75306 201922 75374 201978
rect 75430 201922 75498 201978
rect 75554 201922 75622 201978
rect 75678 201922 75774 201978
rect 75154 184350 75774 201922
rect 75154 184294 75250 184350
rect 75306 184294 75374 184350
rect 75430 184294 75498 184350
rect 75554 184294 75622 184350
rect 75678 184294 75774 184350
rect 75154 184226 75774 184294
rect 75154 184170 75250 184226
rect 75306 184170 75374 184226
rect 75430 184170 75498 184226
rect 75554 184170 75622 184226
rect 75678 184170 75774 184226
rect 75154 184102 75774 184170
rect 75154 184046 75250 184102
rect 75306 184046 75374 184102
rect 75430 184046 75498 184102
rect 75554 184046 75622 184102
rect 75678 184046 75774 184102
rect 75154 183978 75774 184046
rect 75154 183922 75250 183978
rect 75306 183922 75374 183978
rect 75430 183922 75498 183978
rect 75554 183922 75622 183978
rect 75678 183922 75774 183978
rect 75154 166350 75774 183922
rect 75154 166294 75250 166350
rect 75306 166294 75374 166350
rect 75430 166294 75498 166350
rect 75554 166294 75622 166350
rect 75678 166294 75774 166350
rect 75154 166226 75774 166294
rect 75154 166170 75250 166226
rect 75306 166170 75374 166226
rect 75430 166170 75498 166226
rect 75554 166170 75622 166226
rect 75678 166170 75774 166226
rect 75154 166102 75774 166170
rect 75154 166046 75250 166102
rect 75306 166046 75374 166102
rect 75430 166046 75498 166102
rect 75554 166046 75622 166102
rect 75678 166046 75774 166102
rect 75154 165978 75774 166046
rect 75154 165922 75250 165978
rect 75306 165922 75374 165978
rect 75430 165922 75498 165978
rect 75554 165922 75622 165978
rect 75678 165922 75774 165978
rect 75154 148350 75774 165922
rect 75154 148294 75250 148350
rect 75306 148294 75374 148350
rect 75430 148294 75498 148350
rect 75554 148294 75622 148350
rect 75678 148294 75774 148350
rect 75154 148226 75774 148294
rect 75154 148170 75250 148226
rect 75306 148170 75374 148226
rect 75430 148170 75498 148226
rect 75554 148170 75622 148226
rect 75678 148170 75774 148226
rect 75154 148102 75774 148170
rect 75154 148046 75250 148102
rect 75306 148046 75374 148102
rect 75430 148046 75498 148102
rect 75554 148046 75622 148102
rect 75678 148046 75774 148102
rect 75154 147978 75774 148046
rect 75154 147922 75250 147978
rect 75306 147922 75374 147978
rect 75430 147922 75498 147978
rect 75554 147922 75622 147978
rect 75678 147922 75774 147978
rect 75154 130350 75774 147922
rect 75154 130294 75250 130350
rect 75306 130294 75374 130350
rect 75430 130294 75498 130350
rect 75554 130294 75622 130350
rect 75678 130294 75774 130350
rect 75154 130226 75774 130294
rect 75154 130170 75250 130226
rect 75306 130170 75374 130226
rect 75430 130170 75498 130226
rect 75554 130170 75622 130226
rect 75678 130170 75774 130226
rect 75154 130102 75774 130170
rect 75154 130046 75250 130102
rect 75306 130046 75374 130102
rect 75430 130046 75498 130102
rect 75554 130046 75622 130102
rect 75678 130046 75774 130102
rect 75154 129978 75774 130046
rect 75154 129922 75250 129978
rect 75306 129922 75374 129978
rect 75430 129922 75498 129978
rect 75554 129922 75622 129978
rect 75678 129922 75774 129978
rect 75154 112350 75774 129922
rect 75154 112294 75250 112350
rect 75306 112294 75374 112350
rect 75430 112294 75498 112350
rect 75554 112294 75622 112350
rect 75678 112294 75774 112350
rect 75154 112226 75774 112294
rect 75154 112170 75250 112226
rect 75306 112170 75374 112226
rect 75430 112170 75498 112226
rect 75554 112170 75622 112226
rect 75678 112170 75774 112226
rect 75154 112102 75774 112170
rect 75154 112046 75250 112102
rect 75306 112046 75374 112102
rect 75430 112046 75498 112102
rect 75554 112046 75622 112102
rect 75678 112046 75774 112102
rect 75154 111978 75774 112046
rect 75154 111922 75250 111978
rect 75306 111922 75374 111978
rect 75430 111922 75498 111978
rect 75554 111922 75622 111978
rect 75678 111922 75774 111978
rect 75154 94350 75774 111922
rect 75154 94294 75250 94350
rect 75306 94294 75374 94350
rect 75430 94294 75498 94350
rect 75554 94294 75622 94350
rect 75678 94294 75774 94350
rect 75154 94226 75774 94294
rect 75154 94170 75250 94226
rect 75306 94170 75374 94226
rect 75430 94170 75498 94226
rect 75554 94170 75622 94226
rect 75678 94170 75774 94226
rect 75154 94102 75774 94170
rect 75154 94046 75250 94102
rect 75306 94046 75374 94102
rect 75430 94046 75498 94102
rect 75554 94046 75622 94102
rect 75678 94046 75774 94102
rect 75154 93978 75774 94046
rect 75154 93922 75250 93978
rect 75306 93922 75374 93978
rect 75430 93922 75498 93978
rect 75554 93922 75622 93978
rect 75678 93922 75774 93978
rect 75154 76350 75774 93922
rect 75154 76294 75250 76350
rect 75306 76294 75374 76350
rect 75430 76294 75498 76350
rect 75554 76294 75622 76350
rect 75678 76294 75774 76350
rect 75154 76226 75774 76294
rect 75154 76170 75250 76226
rect 75306 76170 75374 76226
rect 75430 76170 75498 76226
rect 75554 76170 75622 76226
rect 75678 76170 75774 76226
rect 75154 76102 75774 76170
rect 75154 76046 75250 76102
rect 75306 76046 75374 76102
rect 75430 76046 75498 76102
rect 75554 76046 75622 76102
rect 75678 76046 75774 76102
rect 75154 75978 75774 76046
rect 75154 75922 75250 75978
rect 75306 75922 75374 75978
rect 75430 75922 75498 75978
rect 75554 75922 75622 75978
rect 75678 75922 75774 75978
rect 75154 58350 75774 75922
rect 75154 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 75774 58350
rect 75154 58226 75774 58294
rect 75154 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 75774 58226
rect 75154 58102 75774 58170
rect 75154 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 75774 58102
rect 75154 57978 75774 58046
rect 75154 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 75774 57978
rect 75154 40350 75774 57922
rect 75154 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 75774 40350
rect 75154 40226 75774 40294
rect 75154 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 75774 40226
rect 75154 40102 75774 40170
rect 75154 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 75774 40102
rect 75154 39978 75774 40046
rect 75154 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 75774 39978
rect 75154 22350 75774 39922
rect 75154 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 75774 22350
rect 75154 22226 75774 22294
rect 75154 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 75774 22226
rect 75154 22102 75774 22170
rect 75154 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 75774 22102
rect 75154 21978 75774 22046
rect 75154 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 75774 21978
rect 75154 4350 75774 21922
rect 75154 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 75774 4350
rect 75154 4226 75774 4294
rect 75154 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 75774 4226
rect 75154 4102 75774 4170
rect 75154 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 75774 4102
rect 75154 3978 75774 4046
rect 75154 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 75774 3978
rect 75154 -160 75774 3922
rect 75154 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 75774 -160
rect 75154 -284 75774 -216
rect 75154 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 75774 -284
rect 75154 -408 75774 -340
rect 75154 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 75774 -408
rect 75154 -532 75774 -464
rect 75154 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 75774 -532
rect 75154 -1644 75774 -588
rect 78874 598172 79494 598268
rect 78874 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 79494 598172
rect 78874 598048 79494 598116
rect 78874 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 79494 598048
rect 78874 597924 79494 597992
rect 78874 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 79494 597924
rect 78874 597800 79494 597868
rect 78874 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 79494 597800
rect 78874 586350 79494 597744
rect 78874 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 79494 586350
rect 78874 586226 79494 586294
rect 78874 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 79494 586226
rect 78874 586102 79494 586170
rect 78874 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 79494 586102
rect 78874 585978 79494 586046
rect 78874 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 79494 585978
rect 78874 568350 79494 585922
rect 78874 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 79494 568350
rect 78874 568226 79494 568294
rect 78874 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 79494 568226
rect 78874 568102 79494 568170
rect 78874 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 79494 568102
rect 78874 567978 79494 568046
rect 78874 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 79494 567978
rect 78874 550350 79494 567922
rect 78874 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 79494 550350
rect 78874 550226 79494 550294
rect 78874 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 79494 550226
rect 78874 550102 79494 550170
rect 78874 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 79494 550102
rect 78874 549978 79494 550046
rect 78874 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 79494 549978
rect 78874 532350 79494 549922
rect 78874 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 79494 532350
rect 78874 532226 79494 532294
rect 78874 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 79494 532226
rect 78874 532102 79494 532170
rect 78874 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 79494 532102
rect 78874 531978 79494 532046
rect 78874 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 79494 531978
rect 78874 514350 79494 531922
rect 78874 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 79494 514350
rect 78874 514226 79494 514294
rect 78874 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 79494 514226
rect 78874 514102 79494 514170
rect 78874 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 79494 514102
rect 78874 513978 79494 514046
rect 78874 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 79494 513978
rect 78874 496350 79494 513922
rect 78874 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 79494 496350
rect 78874 496226 79494 496294
rect 78874 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 79494 496226
rect 78874 496102 79494 496170
rect 78874 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 79494 496102
rect 78874 495978 79494 496046
rect 78874 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 79494 495978
rect 78874 478350 79494 495922
rect 78874 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 79494 478350
rect 78874 478226 79494 478294
rect 78874 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 79494 478226
rect 78874 478102 79494 478170
rect 78874 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 79494 478102
rect 78874 477978 79494 478046
rect 78874 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 79494 477978
rect 78874 460350 79494 477922
rect 78874 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 79494 460350
rect 78874 460226 79494 460294
rect 78874 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 79494 460226
rect 78874 460102 79494 460170
rect 78874 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 79494 460102
rect 78874 459978 79494 460046
rect 78874 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 79494 459978
rect 78874 442350 79494 459922
rect 78874 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 79494 442350
rect 78874 442226 79494 442294
rect 78874 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 79494 442226
rect 78874 442102 79494 442170
rect 78874 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 79494 442102
rect 78874 441978 79494 442046
rect 78874 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 79494 441978
rect 78874 424350 79494 441922
rect 78874 424294 78970 424350
rect 79026 424294 79094 424350
rect 79150 424294 79218 424350
rect 79274 424294 79342 424350
rect 79398 424294 79494 424350
rect 78874 424226 79494 424294
rect 78874 424170 78970 424226
rect 79026 424170 79094 424226
rect 79150 424170 79218 424226
rect 79274 424170 79342 424226
rect 79398 424170 79494 424226
rect 78874 424102 79494 424170
rect 78874 424046 78970 424102
rect 79026 424046 79094 424102
rect 79150 424046 79218 424102
rect 79274 424046 79342 424102
rect 79398 424046 79494 424102
rect 78874 423978 79494 424046
rect 78874 423922 78970 423978
rect 79026 423922 79094 423978
rect 79150 423922 79218 423978
rect 79274 423922 79342 423978
rect 79398 423922 79494 423978
rect 78874 406350 79494 423922
rect 78874 406294 78970 406350
rect 79026 406294 79094 406350
rect 79150 406294 79218 406350
rect 79274 406294 79342 406350
rect 79398 406294 79494 406350
rect 78874 406226 79494 406294
rect 78874 406170 78970 406226
rect 79026 406170 79094 406226
rect 79150 406170 79218 406226
rect 79274 406170 79342 406226
rect 79398 406170 79494 406226
rect 78874 406102 79494 406170
rect 78874 406046 78970 406102
rect 79026 406046 79094 406102
rect 79150 406046 79218 406102
rect 79274 406046 79342 406102
rect 79398 406046 79494 406102
rect 78874 405978 79494 406046
rect 78874 405922 78970 405978
rect 79026 405922 79094 405978
rect 79150 405922 79218 405978
rect 79274 405922 79342 405978
rect 79398 405922 79494 405978
rect 78874 388350 79494 405922
rect 78874 388294 78970 388350
rect 79026 388294 79094 388350
rect 79150 388294 79218 388350
rect 79274 388294 79342 388350
rect 79398 388294 79494 388350
rect 78874 388226 79494 388294
rect 78874 388170 78970 388226
rect 79026 388170 79094 388226
rect 79150 388170 79218 388226
rect 79274 388170 79342 388226
rect 79398 388170 79494 388226
rect 78874 388102 79494 388170
rect 78874 388046 78970 388102
rect 79026 388046 79094 388102
rect 79150 388046 79218 388102
rect 79274 388046 79342 388102
rect 79398 388046 79494 388102
rect 78874 387978 79494 388046
rect 78874 387922 78970 387978
rect 79026 387922 79094 387978
rect 79150 387922 79218 387978
rect 79274 387922 79342 387978
rect 79398 387922 79494 387978
rect 78874 370350 79494 387922
rect 78874 370294 78970 370350
rect 79026 370294 79094 370350
rect 79150 370294 79218 370350
rect 79274 370294 79342 370350
rect 79398 370294 79494 370350
rect 78874 370226 79494 370294
rect 78874 370170 78970 370226
rect 79026 370170 79094 370226
rect 79150 370170 79218 370226
rect 79274 370170 79342 370226
rect 79398 370170 79494 370226
rect 78874 370102 79494 370170
rect 78874 370046 78970 370102
rect 79026 370046 79094 370102
rect 79150 370046 79218 370102
rect 79274 370046 79342 370102
rect 79398 370046 79494 370102
rect 78874 369978 79494 370046
rect 78874 369922 78970 369978
rect 79026 369922 79094 369978
rect 79150 369922 79218 369978
rect 79274 369922 79342 369978
rect 79398 369922 79494 369978
rect 78874 352350 79494 369922
rect 78874 352294 78970 352350
rect 79026 352294 79094 352350
rect 79150 352294 79218 352350
rect 79274 352294 79342 352350
rect 79398 352294 79494 352350
rect 78874 352226 79494 352294
rect 78874 352170 78970 352226
rect 79026 352170 79094 352226
rect 79150 352170 79218 352226
rect 79274 352170 79342 352226
rect 79398 352170 79494 352226
rect 78874 352102 79494 352170
rect 78874 352046 78970 352102
rect 79026 352046 79094 352102
rect 79150 352046 79218 352102
rect 79274 352046 79342 352102
rect 79398 352046 79494 352102
rect 78874 351978 79494 352046
rect 78874 351922 78970 351978
rect 79026 351922 79094 351978
rect 79150 351922 79218 351978
rect 79274 351922 79342 351978
rect 79398 351922 79494 351978
rect 78874 334350 79494 351922
rect 78874 334294 78970 334350
rect 79026 334294 79094 334350
rect 79150 334294 79218 334350
rect 79274 334294 79342 334350
rect 79398 334294 79494 334350
rect 78874 334226 79494 334294
rect 78874 334170 78970 334226
rect 79026 334170 79094 334226
rect 79150 334170 79218 334226
rect 79274 334170 79342 334226
rect 79398 334170 79494 334226
rect 78874 334102 79494 334170
rect 78874 334046 78970 334102
rect 79026 334046 79094 334102
rect 79150 334046 79218 334102
rect 79274 334046 79342 334102
rect 79398 334046 79494 334102
rect 78874 333978 79494 334046
rect 78874 333922 78970 333978
rect 79026 333922 79094 333978
rect 79150 333922 79218 333978
rect 79274 333922 79342 333978
rect 79398 333922 79494 333978
rect 78874 316350 79494 333922
rect 78874 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 79494 316350
rect 78874 316226 79494 316294
rect 78874 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 79494 316226
rect 78874 316102 79494 316170
rect 78874 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 79494 316102
rect 78874 315978 79494 316046
rect 78874 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 79494 315978
rect 78874 298350 79494 315922
rect 78874 298294 78970 298350
rect 79026 298294 79094 298350
rect 79150 298294 79218 298350
rect 79274 298294 79342 298350
rect 79398 298294 79494 298350
rect 78874 298226 79494 298294
rect 78874 298170 78970 298226
rect 79026 298170 79094 298226
rect 79150 298170 79218 298226
rect 79274 298170 79342 298226
rect 79398 298170 79494 298226
rect 78874 298102 79494 298170
rect 78874 298046 78970 298102
rect 79026 298046 79094 298102
rect 79150 298046 79218 298102
rect 79274 298046 79342 298102
rect 79398 298046 79494 298102
rect 78874 297978 79494 298046
rect 78874 297922 78970 297978
rect 79026 297922 79094 297978
rect 79150 297922 79218 297978
rect 79274 297922 79342 297978
rect 79398 297922 79494 297978
rect 78874 280350 79494 297922
rect 78874 280294 78970 280350
rect 79026 280294 79094 280350
rect 79150 280294 79218 280350
rect 79274 280294 79342 280350
rect 79398 280294 79494 280350
rect 78874 280226 79494 280294
rect 78874 280170 78970 280226
rect 79026 280170 79094 280226
rect 79150 280170 79218 280226
rect 79274 280170 79342 280226
rect 79398 280170 79494 280226
rect 78874 280102 79494 280170
rect 78874 280046 78970 280102
rect 79026 280046 79094 280102
rect 79150 280046 79218 280102
rect 79274 280046 79342 280102
rect 79398 280046 79494 280102
rect 78874 279978 79494 280046
rect 78874 279922 78970 279978
rect 79026 279922 79094 279978
rect 79150 279922 79218 279978
rect 79274 279922 79342 279978
rect 79398 279922 79494 279978
rect 78874 262350 79494 279922
rect 78874 262294 78970 262350
rect 79026 262294 79094 262350
rect 79150 262294 79218 262350
rect 79274 262294 79342 262350
rect 79398 262294 79494 262350
rect 78874 262226 79494 262294
rect 78874 262170 78970 262226
rect 79026 262170 79094 262226
rect 79150 262170 79218 262226
rect 79274 262170 79342 262226
rect 79398 262170 79494 262226
rect 78874 262102 79494 262170
rect 78874 262046 78970 262102
rect 79026 262046 79094 262102
rect 79150 262046 79218 262102
rect 79274 262046 79342 262102
rect 79398 262046 79494 262102
rect 78874 261978 79494 262046
rect 78874 261922 78970 261978
rect 79026 261922 79094 261978
rect 79150 261922 79218 261978
rect 79274 261922 79342 261978
rect 79398 261922 79494 261978
rect 78874 244350 79494 261922
rect 78874 244294 78970 244350
rect 79026 244294 79094 244350
rect 79150 244294 79218 244350
rect 79274 244294 79342 244350
rect 79398 244294 79494 244350
rect 78874 244226 79494 244294
rect 78874 244170 78970 244226
rect 79026 244170 79094 244226
rect 79150 244170 79218 244226
rect 79274 244170 79342 244226
rect 79398 244170 79494 244226
rect 78874 244102 79494 244170
rect 78874 244046 78970 244102
rect 79026 244046 79094 244102
rect 79150 244046 79218 244102
rect 79274 244046 79342 244102
rect 79398 244046 79494 244102
rect 78874 243978 79494 244046
rect 78874 243922 78970 243978
rect 79026 243922 79094 243978
rect 79150 243922 79218 243978
rect 79274 243922 79342 243978
rect 79398 243922 79494 243978
rect 78874 226350 79494 243922
rect 78874 226294 78970 226350
rect 79026 226294 79094 226350
rect 79150 226294 79218 226350
rect 79274 226294 79342 226350
rect 79398 226294 79494 226350
rect 78874 226226 79494 226294
rect 78874 226170 78970 226226
rect 79026 226170 79094 226226
rect 79150 226170 79218 226226
rect 79274 226170 79342 226226
rect 79398 226170 79494 226226
rect 78874 226102 79494 226170
rect 78874 226046 78970 226102
rect 79026 226046 79094 226102
rect 79150 226046 79218 226102
rect 79274 226046 79342 226102
rect 79398 226046 79494 226102
rect 78874 225978 79494 226046
rect 78874 225922 78970 225978
rect 79026 225922 79094 225978
rect 79150 225922 79218 225978
rect 79274 225922 79342 225978
rect 79398 225922 79494 225978
rect 78874 208350 79494 225922
rect 78874 208294 78970 208350
rect 79026 208294 79094 208350
rect 79150 208294 79218 208350
rect 79274 208294 79342 208350
rect 79398 208294 79494 208350
rect 78874 208226 79494 208294
rect 78874 208170 78970 208226
rect 79026 208170 79094 208226
rect 79150 208170 79218 208226
rect 79274 208170 79342 208226
rect 79398 208170 79494 208226
rect 78874 208102 79494 208170
rect 78874 208046 78970 208102
rect 79026 208046 79094 208102
rect 79150 208046 79218 208102
rect 79274 208046 79342 208102
rect 79398 208046 79494 208102
rect 78874 207978 79494 208046
rect 78874 207922 78970 207978
rect 79026 207922 79094 207978
rect 79150 207922 79218 207978
rect 79274 207922 79342 207978
rect 79398 207922 79494 207978
rect 78874 190350 79494 207922
rect 78874 190294 78970 190350
rect 79026 190294 79094 190350
rect 79150 190294 79218 190350
rect 79274 190294 79342 190350
rect 79398 190294 79494 190350
rect 78874 190226 79494 190294
rect 78874 190170 78970 190226
rect 79026 190170 79094 190226
rect 79150 190170 79218 190226
rect 79274 190170 79342 190226
rect 79398 190170 79494 190226
rect 78874 190102 79494 190170
rect 78874 190046 78970 190102
rect 79026 190046 79094 190102
rect 79150 190046 79218 190102
rect 79274 190046 79342 190102
rect 79398 190046 79494 190102
rect 78874 189978 79494 190046
rect 78874 189922 78970 189978
rect 79026 189922 79094 189978
rect 79150 189922 79218 189978
rect 79274 189922 79342 189978
rect 79398 189922 79494 189978
rect 78874 172350 79494 189922
rect 78874 172294 78970 172350
rect 79026 172294 79094 172350
rect 79150 172294 79218 172350
rect 79274 172294 79342 172350
rect 79398 172294 79494 172350
rect 78874 172226 79494 172294
rect 78874 172170 78970 172226
rect 79026 172170 79094 172226
rect 79150 172170 79218 172226
rect 79274 172170 79342 172226
rect 79398 172170 79494 172226
rect 78874 172102 79494 172170
rect 78874 172046 78970 172102
rect 79026 172046 79094 172102
rect 79150 172046 79218 172102
rect 79274 172046 79342 172102
rect 79398 172046 79494 172102
rect 78874 171978 79494 172046
rect 78874 171922 78970 171978
rect 79026 171922 79094 171978
rect 79150 171922 79218 171978
rect 79274 171922 79342 171978
rect 79398 171922 79494 171978
rect 78874 154350 79494 171922
rect 78874 154294 78970 154350
rect 79026 154294 79094 154350
rect 79150 154294 79218 154350
rect 79274 154294 79342 154350
rect 79398 154294 79494 154350
rect 78874 154226 79494 154294
rect 78874 154170 78970 154226
rect 79026 154170 79094 154226
rect 79150 154170 79218 154226
rect 79274 154170 79342 154226
rect 79398 154170 79494 154226
rect 78874 154102 79494 154170
rect 78874 154046 78970 154102
rect 79026 154046 79094 154102
rect 79150 154046 79218 154102
rect 79274 154046 79342 154102
rect 79398 154046 79494 154102
rect 78874 153978 79494 154046
rect 78874 153922 78970 153978
rect 79026 153922 79094 153978
rect 79150 153922 79218 153978
rect 79274 153922 79342 153978
rect 79398 153922 79494 153978
rect 78874 136350 79494 153922
rect 78874 136294 78970 136350
rect 79026 136294 79094 136350
rect 79150 136294 79218 136350
rect 79274 136294 79342 136350
rect 79398 136294 79494 136350
rect 78874 136226 79494 136294
rect 78874 136170 78970 136226
rect 79026 136170 79094 136226
rect 79150 136170 79218 136226
rect 79274 136170 79342 136226
rect 79398 136170 79494 136226
rect 78874 136102 79494 136170
rect 78874 136046 78970 136102
rect 79026 136046 79094 136102
rect 79150 136046 79218 136102
rect 79274 136046 79342 136102
rect 79398 136046 79494 136102
rect 78874 135978 79494 136046
rect 78874 135922 78970 135978
rect 79026 135922 79094 135978
rect 79150 135922 79218 135978
rect 79274 135922 79342 135978
rect 79398 135922 79494 135978
rect 78874 118350 79494 135922
rect 78874 118294 78970 118350
rect 79026 118294 79094 118350
rect 79150 118294 79218 118350
rect 79274 118294 79342 118350
rect 79398 118294 79494 118350
rect 78874 118226 79494 118294
rect 78874 118170 78970 118226
rect 79026 118170 79094 118226
rect 79150 118170 79218 118226
rect 79274 118170 79342 118226
rect 79398 118170 79494 118226
rect 78874 118102 79494 118170
rect 78874 118046 78970 118102
rect 79026 118046 79094 118102
rect 79150 118046 79218 118102
rect 79274 118046 79342 118102
rect 79398 118046 79494 118102
rect 78874 117978 79494 118046
rect 78874 117922 78970 117978
rect 79026 117922 79094 117978
rect 79150 117922 79218 117978
rect 79274 117922 79342 117978
rect 79398 117922 79494 117978
rect 78874 100350 79494 117922
rect 78874 100294 78970 100350
rect 79026 100294 79094 100350
rect 79150 100294 79218 100350
rect 79274 100294 79342 100350
rect 79398 100294 79494 100350
rect 78874 100226 79494 100294
rect 78874 100170 78970 100226
rect 79026 100170 79094 100226
rect 79150 100170 79218 100226
rect 79274 100170 79342 100226
rect 79398 100170 79494 100226
rect 78874 100102 79494 100170
rect 78874 100046 78970 100102
rect 79026 100046 79094 100102
rect 79150 100046 79218 100102
rect 79274 100046 79342 100102
rect 79398 100046 79494 100102
rect 78874 99978 79494 100046
rect 78874 99922 78970 99978
rect 79026 99922 79094 99978
rect 79150 99922 79218 99978
rect 79274 99922 79342 99978
rect 79398 99922 79494 99978
rect 78874 82350 79494 99922
rect 78874 82294 78970 82350
rect 79026 82294 79094 82350
rect 79150 82294 79218 82350
rect 79274 82294 79342 82350
rect 79398 82294 79494 82350
rect 78874 82226 79494 82294
rect 78874 82170 78970 82226
rect 79026 82170 79094 82226
rect 79150 82170 79218 82226
rect 79274 82170 79342 82226
rect 79398 82170 79494 82226
rect 78874 82102 79494 82170
rect 78874 82046 78970 82102
rect 79026 82046 79094 82102
rect 79150 82046 79218 82102
rect 79274 82046 79342 82102
rect 79398 82046 79494 82102
rect 78874 81978 79494 82046
rect 78874 81922 78970 81978
rect 79026 81922 79094 81978
rect 79150 81922 79218 81978
rect 79274 81922 79342 81978
rect 79398 81922 79494 81978
rect 78874 64350 79494 81922
rect 78874 64294 78970 64350
rect 79026 64294 79094 64350
rect 79150 64294 79218 64350
rect 79274 64294 79342 64350
rect 79398 64294 79494 64350
rect 78874 64226 79494 64294
rect 78874 64170 78970 64226
rect 79026 64170 79094 64226
rect 79150 64170 79218 64226
rect 79274 64170 79342 64226
rect 79398 64170 79494 64226
rect 78874 64102 79494 64170
rect 78874 64046 78970 64102
rect 79026 64046 79094 64102
rect 79150 64046 79218 64102
rect 79274 64046 79342 64102
rect 79398 64046 79494 64102
rect 78874 63978 79494 64046
rect 78874 63922 78970 63978
rect 79026 63922 79094 63978
rect 79150 63922 79218 63978
rect 79274 63922 79342 63978
rect 79398 63922 79494 63978
rect 78874 46350 79494 63922
rect 78874 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 79494 46350
rect 78874 46226 79494 46294
rect 78874 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 79494 46226
rect 78874 46102 79494 46170
rect 78874 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 79494 46102
rect 78874 45978 79494 46046
rect 78874 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 79494 45978
rect 78874 28350 79494 45922
rect 78874 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 79494 28350
rect 78874 28226 79494 28294
rect 78874 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 79494 28226
rect 78874 28102 79494 28170
rect 78874 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 79494 28102
rect 78874 27978 79494 28046
rect 78874 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 79494 27978
rect 78874 10350 79494 27922
rect 78874 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 79494 10350
rect 78874 10226 79494 10294
rect 78874 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 79494 10226
rect 78874 10102 79494 10170
rect 78874 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 79494 10102
rect 78874 9978 79494 10046
rect 78874 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 79494 9978
rect 78874 -1120 79494 9922
rect 78874 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 79494 -1120
rect 78874 -1244 79494 -1176
rect 78874 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 79494 -1244
rect 78874 -1368 79494 -1300
rect 78874 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 79494 -1368
rect 78874 -1492 79494 -1424
rect 78874 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 79494 -1492
rect 78874 -1644 79494 -1548
rect 93154 597212 93774 598268
rect 93154 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 93774 597212
rect 93154 597088 93774 597156
rect 93154 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 93774 597088
rect 93154 596964 93774 597032
rect 93154 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 93774 596964
rect 93154 596840 93774 596908
rect 93154 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 93774 596840
rect 93154 580350 93774 596784
rect 93154 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 93774 580350
rect 93154 580226 93774 580294
rect 93154 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 93774 580226
rect 93154 580102 93774 580170
rect 93154 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 93774 580102
rect 93154 579978 93774 580046
rect 93154 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 93774 579978
rect 93154 562350 93774 579922
rect 93154 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 93774 562350
rect 93154 562226 93774 562294
rect 93154 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 93774 562226
rect 93154 562102 93774 562170
rect 93154 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 93774 562102
rect 93154 561978 93774 562046
rect 93154 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 93774 561978
rect 93154 544350 93774 561922
rect 93154 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 93774 544350
rect 93154 544226 93774 544294
rect 93154 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 93774 544226
rect 93154 544102 93774 544170
rect 93154 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 93774 544102
rect 93154 543978 93774 544046
rect 93154 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 93774 543978
rect 93154 526350 93774 543922
rect 93154 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 93774 526350
rect 93154 526226 93774 526294
rect 93154 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 93774 526226
rect 93154 526102 93774 526170
rect 93154 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 93774 526102
rect 93154 525978 93774 526046
rect 93154 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 93774 525978
rect 93154 508350 93774 525922
rect 93154 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 93774 508350
rect 93154 508226 93774 508294
rect 93154 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 93774 508226
rect 93154 508102 93774 508170
rect 93154 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 93774 508102
rect 93154 507978 93774 508046
rect 93154 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 93774 507978
rect 93154 490350 93774 507922
rect 93154 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 93774 490350
rect 93154 490226 93774 490294
rect 93154 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 93774 490226
rect 93154 490102 93774 490170
rect 93154 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 93774 490102
rect 93154 489978 93774 490046
rect 93154 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 93774 489978
rect 93154 472350 93774 489922
rect 93154 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 93774 472350
rect 93154 472226 93774 472294
rect 93154 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 93774 472226
rect 93154 472102 93774 472170
rect 93154 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 93774 472102
rect 93154 471978 93774 472046
rect 93154 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 93774 471978
rect 93154 454350 93774 471922
rect 93154 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 93774 454350
rect 93154 454226 93774 454294
rect 93154 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 93774 454226
rect 93154 454102 93774 454170
rect 93154 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 93774 454102
rect 93154 453978 93774 454046
rect 93154 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 93774 453978
rect 93154 436350 93774 453922
rect 93154 436294 93250 436350
rect 93306 436294 93374 436350
rect 93430 436294 93498 436350
rect 93554 436294 93622 436350
rect 93678 436294 93774 436350
rect 93154 436226 93774 436294
rect 93154 436170 93250 436226
rect 93306 436170 93374 436226
rect 93430 436170 93498 436226
rect 93554 436170 93622 436226
rect 93678 436170 93774 436226
rect 93154 436102 93774 436170
rect 93154 436046 93250 436102
rect 93306 436046 93374 436102
rect 93430 436046 93498 436102
rect 93554 436046 93622 436102
rect 93678 436046 93774 436102
rect 93154 435978 93774 436046
rect 93154 435922 93250 435978
rect 93306 435922 93374 435978
rect 93430 435922 93498 435978
rect 93554 435922 93622 435978
rect 93678 435922 93774 435978
rect 93154 418350 93774 435922
rect 93154 418294 93250 418350
rect 93306 418294 93374 418350
rect 93430 418294 93498 418350
rect 93554 418294 93622 418350
rect 93678 418294 93774 418350
rect 93154 418226 93774 418294
rect 93154 418170 93250 418226
rect 93306 418170 93374 418226
rect 93430 418170 93498 418226
rect 93554 418170 93622 418226
rect 93678 418170 93774 418226
rect 93154 418102 93774 418170
rect 93154 418046 93250 418102
rect 93306 418046 93374 418102
rect 93430 418046 93498 418102
rect 93554 418046 93622 418102
rect 93678 418046 93774 418102
rect 93154 417978 93774 418046
rect 93154 417922 93250 417978
rect 93306 417922 93374 417978
rect 93430 417922 93498 417978
rect 93554 417922 93622 417978
rect 93678 417922 93774 417978
rect 93154 400350 93774 417922
rect 93154 400294 93250 400350
rect 93306 400294 93374 400350
rect 93430 400294 93498 400350
rect 93554 400294 93622 400350
rect 93678 400294 93774 400350
rect 93154 400226 93774 400294
rect 93154 400170 93250 400226
rect 93306 400170 93374 400226
rect 93430 400170 93498 400226
rect 93554 400170 93622 400226
rect 93678 400170 93774 400226
rect 93154 400102 93774 400170
rect 93154 400046 93250 400102
rect 93306 400046 93374 400102
rect 93430 400046 93498 400102
rect 93554 400046 93622 400102
rect 93678 400046 93774 400102
rect 93154 399978 93774 400046
rect 93154 399922 93250 399978
rect 93306 399922 93374 399978
rect 93430 399922 93498 399978
rect 93554 399922 93622 399978
rect 93678 399922 93774 399978
rect 93154 382350 93774 399922
rect 93154 382294 93250 382350
rect 93306 382294 93374 382350
rect 93430 382294 93498 382350
rect 93554 382294 93622 382350
rect 93678 382294 93774 382350
rect 93154 382226 93774 382294
rect 93154 382170 93250 382226
rect 93306 382170 93374 382226
rect 93430 382170 93498 382226
rect 93554 382170 93622 382226
rect 93678 382170 93774 382226
rect 93154 382102 93774 382170
rect 93154 382046 93250 382102
rect 93306 382046 93374 382102
rect 93430 382046 93498 382102
rect 93554 382046 93622 382102
rect 93678 382046 93774 382102
rect 93154 381978 93774 382046
rect 93154 381922 93250 381978
rect 93306 381922 93374 381978
rect 93430 381922 93498 381978
rect 93554 381922 93622 381978
rect 93678 381922 93774 381978
rect 93154 364350 93774 381922
rect 93154 364294 93250 364350
rect 93306 364294 93374 364350
rect 93430 364294 93498 364350
rect 93554 364294 93622 364350
rect 93678 364294 93774 364350
rect 93154 364226 93774 364294
rect 93154 364170 93250 364226
rect 93306 364170 93374 364226
rect 93430 364170 93498 364226
rect 93554 364170 93622 364226
rect 93678 364170 93774 364226
rect 93154 364102 93774 364170
rect 93154 364046 93250 364102
rect 93306 364046 93374 364102
rect 93430 364046 93498 364102
rect 93554 364046 93622 364102
rect 93678 364046 93774 364102
rect 93154 363978 93774 364046
rect 93154 363922 93250 363978
rect 93306 363922 93374 363978
rect 93430 363922 93498 363978
rect 93554 363922 93622 363978
rect 93678 363922 93774 363978
rect 93154 346350 93774 363922
rect 93154 346294 93250 346350
rect 93306 346294 93374 346350
rect 93430 346294 93498 346350
rect 93554 346294 93622 346350
rect 93678 346294 93774 346350
rect 93154 346226 93774 346294
rect 93154 346170 93250 346226
rect 93306 346170 93374 346226
rect 93430 346170 93498 346226
rect 93554 346170 93622 346226
rect 93678 346170 93774 346226
rect 93154 346102 93774 346170
rect 93154 346046 93250 346102
rect 93306 346046 93374 346102
rect 93430 346046 93498 346102
rect 93554 346046 93622 346102
rect 93678 346046 93774 346102
rect 93154 345978 93774 346046
rect 93154 345922 93250 345978
rect 93306 345922 93374 345978
rect 93430 345922 93498 345978
rect 93554 345922 93622 345978
rect 93678 345922 93774 345978
rect 93154 328350 93774 345922
rect 93154 328294 93250 328350
rect 93306 328294 93374 328350
rect 93430 328294 93498 328350
rect 93554 328294 93622 328350
rect 93678 328294 93774 328350
rect 93154 328226 93774 328294
rect 93154 328170 93250 328226
rect 93306 328170 93374 328226
rect 93430 328170 93498 328226
rect 93554 328170 93622 328226
rect 93678 328170 93774 328226
rect 93154 328102 93774 328170
rect 93154 328046 93250 328102
rect 93306 328046 93374 328102
rect 93430 328046 93498 328102
rect 93554 328046 93622 328102
rect 93678 328046 93774 328102
rect 93154 327978 93774 328046
rect 93154 327922 93250 327978
rect 93306 327922 93374 327978
rect 93430 327922 93498 327978
rect 93554 327922 93622 327978
rect 93678 327922 93774 327978
rect 93154 310350 93774 327922
rect 93154 310294 93250 310350
rect 93306 310294 93374 310350
rect 93430 310294 93498 310350
rect 93554 310294 93622 310350
rect 93678 310294 93774 310350
rect 93154 310226 93774 310294
rect 93154 310170 93250 310226
rect 93306 310170 93374 310226
rect 93430 310170 93498 310226
rect 93554 310170 93622 310226
rect 93678 310170 93774 310226
rect 93154 310102 93774 310170
rect 93154 310046 93250 310102
rect 93306 310046 93374 310102
rect 93430 310046 93498 310102
rect 93554 310046 93622 310102
rect 93678 310046 93774 310102
rect 93154 309978 93774 310046
rect 93154 309922 93250 309978
rect 93306 309922 93374 309978
rect 93430 309922 93498 309978
rect 93554 309922 93622 309978
rect 93678 309922 93774 309978
rect 93154 292350 93774 309922
rect 93154 292294 93250 292350
rect 93306 292294 93374 292350
rect 93430 292294 93498 292350
rect 93554 292294 93622 292350
rect 93678 292294 93774 292350
rect 93154 292226 93774 292294
rect 93154 292170 93250 292226
rect 93306 292170 93374 292226
rect 93430 292170 93498 292226
rect 93554 292170 93622 292226
rect 93678 292170 93774 292226
rect 93154 292102 93774 292170
rect 93154 292046 93250 292102
rect 93306 292046 93374 292102
rect 93430 292046 93498 292102
rect 93554 292046 93622 292102
rect 93678 292046 93774 292102
rect 93154 291978 93774 292046
rect 93154 291922 93250 291978
rect 93306 291922 93374 291978
rect 93430 291922 93498 291978
rect 93554 291922 93622 291978
rect 93678 291922 93774 291978
rect 93154 274350 93774 291922
rect 93154 274294 93250 274350
rect 93306 274294 93374 274350
rect 93430 274294 93498 274350
rect 93554 274294 93622 274350
rect 93678 274294 93774 274350
rect 93154 274226 93774 274294
rect 93154 274170 93250 274226
rect 93306 274170 93374 274226
rect 93430 274170 93498 274226
rect 93554 274170 93622 274226
rect 93678 274170 93774 274226
rect 93154 274102 93774 274170
rect 93154 274046 93250 274102
rect 93306 274046 93374 274102
rect 93430 274046 93498 274102
rect 93554 274046 93622 274102
rect 93678 274046 93774 274102
rect 93154 273978 93774 274046
rect 93154 273922 93250 273978
rect 93306 273922 93374 273978
rect 93430 273922 93498 273978
rect 93554 273922 93622 273978
rect 93678 273922 93774 273978
rect 93154 256350 93774 273922
rect 93154 256294 93250 256350
rect 93306 256294 93374 256350
rect 93430 256294 93498 256350
rect 93554 256294 93622 256350
rect 93678 256294 93774 256350
rect 93154 256226 93774 256294
rect 93154 256170 93250 256226
rect 93306 256170 93374 256226
rect 93430 256170 93498 256226
rect 93554 256170 93622 256226
rect 93678 256170 93774 256226
rect 93154 256102 93774 256170
rect 93154 256046 93250 256102
rect 93306 256046 93374 256102
rect 93430 256046 93498 256102
rect 93554 256046 93622 256102
rect 93678 256046 93774 256102
rect 93154 255978 93774 256046
rect 93154 255922 93250 255978
rect 93306 255922 93374 255978
rect 93430 255922 93498 255978
rect 93554 255922 93622 255978
rect 93678 255922 93774 255978
rect 93154 238350 93774 255922
rect 93154 238294 93250 238350
rect 93306 238294 93374 238350
rect 93430 238294 93498 238350
rect 93554 238294 93622 238350
rect 93678 238294 93774 238350
rect 93154 238226 93774 238294
rect 93154 238170 93250 238226
rect 93306 238170 93374 238226
rect 93430 238170 93498 238226
rect 93554 238170 93622 238226
rect 93678 238170 93774 238226
rect 93154 238102 93774 238170
rect 93154 238046 93250 238102
rect 93306 238046 93374 238102
rect 93430 238046 93498 238102
rect 93554 238046 93622 238102
rect 93678 238046 93774 238102
rect 93154 237978 93774 238046
rect 93154 237922 93250 237978
rect 93306 237922 93374 237978
rect 93430 237922 93498 237978
rect 93554 237922 93622 237978
rect 93678 237922 93774 237978
rect 93154 220350 93774 237922
rect 93154 220294 93250 220350
rect 93306 220294 93374 220350
rect 93430 220294 93498 220350
rect 93554 220294 93622 220350
rect 93678 220294 93774 220350
rect 93154 220226 93774 220294
rect 93154 220170 93250 220226
rect 93306 220170 93374 220226
rect 93430 220170 93498 220226
rect 93554 220170 93622 220226
rect 93678 220170 93774 220226
rect 93154 220102 93774 220170
rect 93154 220046 93250 220102
rect 93306 220046 93374 220102
rect 93430 220046 93498 220102
rect 93554 220046 93622 220102
rect 93678 220046 93774 220102
rect 93154 219978 93774 220046
rect 93154 219922 93250 219978
rect 93306 219922 93374 219978
rect 93430 219922 93498 219978
rect 93554 219922 93622 219978
rect 93678 219922 93774 219978
rect 93154 202350 93774 219922
rect 93154 202294 93250 202350
rect 93306 202294 93374 202350
rect 93430 202294 93498 202350
rect 93554 202294 93622 202350
rect 93678 202294 93774 202350
rect 93154 202226 93774 202294
rect 93154 202170 93250 202226
rect 93306 202170 93374 202226
rect 93430 202170 93498 202226
rect 93554 202170 93622 202226
rect 93678 202170 93774 202226
rect 93154 202102 93774 202170
rect 93154 202046 93250 202102
rect 93306 202046 93374 202102
rect 93430 202046 93498 202102
rect 93554 202046 93622 202102
rect 93678 202046 93774 202102
rect 93154 201978 93774 202046
rect 93154 201922 93250 201978
rect 93306 201922 93374 201978
rect 93430 201922 93498 201978
rect 93554 201922 93622 201978
rect 93678 201922 93774 201978
rect 93154 184350 93774 201922
rect 93154 184294 93250 184350
rect 93306 184294 93374 184350
rect 93430 184294 93498 184350
rect 93554 184294 93622 184350
rect 93678 184294 93774 184350
rect 93154 184226 93774 184294
rect 93154 184170 93250 184226
rect 93306 184170 93374 184226
rect 93430 184170 93498 184226
rect 93554 184170 93622 184226
rect 93678 184170 93774 184226
rect 93154 184102 93774 184170
rect 93154 184046 93250 184102
rect 93306 184046 93374 184102
rect 93430 184046 93498 184102
rect 93554 184046 93622 184102
rect 93678 184046 93774 184102
rect 93154 183978 93774 184046
rect 93154 183922 93250 183978
rect 93306 183922 93374 183978
rect 93430 183922 93498 183978
rect 93554 183922 93622 183978
rect 93678 183922 93774 183978
rect 93154 166350 93774 183922
rect 93154 166294 93250 166350
rect 93306 166294 93374 166350
rect 93430 166294 93498 166350
rect 93554 166294 93622 166350
rect 93678 166294 93774 166350
rect 93154 166226 93774 166294
rect 93154 166170 93250 166226
rect 93306 166170 93374 166226
rect 93430 166170 93498 166226
rect 93554 166170 93622 166226
rect 93678 166170 93774 166226
rect 93154 166102 93774 166170
rect 93154 166046 93250 166102
rect 93306 166046 93374 166102
rect 93430 166046 93498 166102
rect 93554 166046 93622 166102
rect 93678 166046 93774 166102
rect 93154 165978 93774 166046
rect 93154 165922 93250 165978
rect 93306 165922 93374 165978
rect 93430 165922 93498 165978
rect 93554 165922 93622 165978
rect 93678 165922 93774 165978
rect 93154 148350 93774 165922
rect 93154 148294 93250 148350
rect 93306 148294 93374 148350
rect 93430 148294 93498 148350
rect 93554 148294 93622 148350
rect 93678 148294 93774 148350
rect 93154 148226 93774 148294
rect 93154 148170 93250 148226
rect 93306 148170 93374 148226
rect 93430 148170 93498 148226
rect 93554 148170 93622 148226
rect 93678 148170 93774 148226
rect 93154 148102 93774 148170
rect 93154 148046 93250 148102
rect 93306 148046 93374 148102
rect 93430 148046 93498 148102
rect 93554 148046 93622 148102
rect 93678 148046 93774 148102
rect 93154 147978 93774 148046
rect 93154 147922 93250 147978
rect 93306 147922 93374 147978
rect 93430 147922 93498 147978
rect 93554 147922 93622 147978
rect 93678 147922 93774 147978
rect 93154 130350 93774 147922
rect 93154 130294 93250 130350
rect 93306 130294 93374 130350
rect 93430 130294 93498 130350
rect 93554 130294 93622 130350
rect 93678 130294 93774 130350
rect 93154 130226 93774 130294
rect 93154 130170 93250 130226
rect 93306 130170 93374 130226
rect 93430 130170 93498 130226
rect 93554 130170 93622 130226
rect 93678 130170 93774 130226
rect 93154 130102 93774 130170
rect 93154 130046 93250 130102
rect 93306 130046 93374 130102
rect 93430 130046 93498 130102
rect 93554 130046 93622 130102
rect 93678 130046 93774 130102
rect 93154 129978 93774 130046
rect 93154 129922 93250 129978
rect 93306 129922 93374 129978
rect 93430 129922 93498 129978
rect 93554 129922 93622 129978
rect 93678 129922 93774 129978
rect 93154 112350 93774 129922
rect 93154 112294 93250 112350
rect 93306 112294 93374 112350
rect 93430 112294 93498 112350
rect 93554 112294 93622 112350
rect 93678 112294 93774 112350
rect 93154 112226 93774 112294
rect 93154 112170 93250 112226
rect 93306 112170 93374 112226
rect 93430 112170 93498 112226
rect 93554 112170 93622 112226
rect 93678 112170 93774 112226
rect 93154 112102 93774 112170
rect 93154 112046 93250 112102
rect 93306 112046 93374 112102
rect 93430 112046 93498 112102
rect 93554 112046 93622 112102
rect 93678 112046 93774 112102
rect 93154 111978 93774 112046
rect 93154 111922 93250 111978
rect 93306 111922 93374 111978
rect 93430 111922 93498 111978
rect 93554 111922 93622 111978
rect 93678 111922 93774 111978
rect 93154 94350 93774 111922
rect 93154 94294 93250 94350
rect 93306 94294 93374 94350
rect 93430 94294 93498 94350
rect 93554 94294 93622 94350
rect 93678 94294 93774 94350
rect 93154 94226 93774 94294
rect 93154 94170 93250 94226
rect 93306 94170 93374 94226
rect 93430 94170 93498 94226
rect 93554 94170 93622 94226
rect 93678 94170 93774 94226
rect 93154 94102 93774 94170
rect 93154 94046 93250 94102
rect 93306 94046 93374 94102
rect 93430 94046 93498 94102
rect 93554 94046 93622 94102
rect 93678 94046 93774 94102
rect 93154 93978 93774 94046
rect 93154 93922 93250 93978
rect 93306 93922 93374 93978
rect 93430 93922 93498 93978
rect 93554 93922 93622 93978
rect 93678 93922 93774 93978
rect 93154 76350 93774 93922
rect 93154 76294 93250 76350
rect 93306 76294 93374 76350
rect 93430 76294 93498 76350
rect 93554 76294 93622 76350
rect 93678 76294 93774 76350
rect 93154 76226 93774 76294
rect 93154 76170 93250 76226
rect 93306 76170 93374 76226
rect 93430 76170 93498 76226
rect 93554 76170 93622 76226
rect 93678 76170 93774 76226
rect 93154 76102 93774 76170
rect 93154 76046 93250 76102
rect 93306 76046 93374 76102
rect 93430 76046 93498 76102
rect 93554 76046 93622 76102
rect 93678 76046 93774 76102
rect 93154 75978 93774 76046
rect 93154 75922 93250 75978
rect 93306 75922 93374 75978
rect 93430 75922 93498 75978
rect 93554 75922 93622 75978
rect 93678 75922 93774 75978
rect 93154 58350 93774 75922
rect 93154 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 93774 58350
rect 93154 58226 93774 58294
rect 93154 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 93774 58226
rect 93154 58102 93774 58170
rect 93154 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 93774 58102
rect 93154 57978 93774 58046
rect 93154 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 93774 57978
rect 93154 40350 93774 57922
rect 93154 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 93774 40350
rect 93154 40226 93774 40294
rect 93154 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 93774 40226
rect 93154 40102 93774 40170
rect 93154 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 93774 40102
rect 93154 39978 93774 40046
rect 93154 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 93774 39978
rect 93154 22350 93774 39922
rect 93154 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 93774 22350
rect 93154 22226 93774 22294
rect 93154 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 93774 22226
rect 93154 22102 93774 22170
rect 93154 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 93774 22102
rect 93154 21978 93774 22046
rect 93154 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 93774 21978
rect 93154 4350 93774 21922
rect 93154 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 93774 4350
rect 93154 4226 93774 4294
rect 93154 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 93774 4226
rect 93154 4102 93774 4170
rect 93154 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 93774 4102
rect 93154 3978 93774 4046
rect 93154 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 93774 3978
rect 93154 -160 93774 3922
rect 93154 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 93774 -160
rect 93154 -284 93774 -216
rect 93154 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 93774 -284
rect 93154 -408 93774 -340
rect 93154 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 93774 -408
rect 93154 -532 93774 -464
rect 93154 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 93774 -532
rect 93154 -1644 93774 -588
rect 96874 598172 97494 598268
rect 96874 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 97494 598172
rect 96874 598048 97494 598116
rect 96874 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 97494 598048
rect 96874 597924 97494 597992
rect 96874 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 97494 597924
rect 96874 597800 97494 597868
rect 96874 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 97494 597800
rect 96874 586350 97494 597744
rect 96874 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 97494 586350
rect 96874 586226 97494 586294
rect 96874 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 97494 586226
rect 96874 586102 97494 586170
rect 96874 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 97494 586102
rect 96874 585978 97494 586046
rect 96874 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 97494 585978
rect 96874 568350 97494 585922
rect 96874 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 97494 568350
rect 96874 568226 97494 568294
rect 96874 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 97494 568226
rect 96874 568102 97494 568170
rect 96874 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 97494 568102
rect 96874 567978 97494 568046
rect 96874 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 97494 567978
rect 96874 550350 97494 567922
rect 96874 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 97494 550350
rect 96874 550226 97494 550294
rect 96874 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 97494 550226
rect 96874 550102 97494 550170
rect 96874 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 97494 550102
rect 96874 549978 97494 550046
rect 96874 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 97494 549978
rect 96874 532350 97494 549922
rect 96874 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 97494 532350
rect 96874 532226 97494 532294
rect 96874 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 97494 532226
rect 96874 532102 97494 532170
rect 96874 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 97494 532102
rect 96874 531978 97494 532046
rect 96874 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 97494 531978
rect 96874 514350 97494 531922
rect 96874 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 97494 514350
rect 96874 514226 97494 514294
rect 96874 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 97494 514226
rect 96874 514102 97494 514170
rect 96874 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 97494 514102
rect 96874 513978 97494 514046
rect 96874 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 97494 513978
rect 96874 496350 97494 513922
rect 96874 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 97494 496350
rect 96874 496226 97494 496294
rect 96874 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 97494 496226
rect 96874 496102 97494 496170
rect 96874 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 97494 496102
rect 96874 495978 97494 496046
rect 96874 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 97494 495978
rect 96874 478350 97494 495922
rect 96874 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 97494 478350
rect 96874 478226 97494 478294
rect 96874 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 97494 478226
rect 96874 478102 97494 478170
rect 96874 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 97494 478102
rect 96874 477978 97494 478046
rect 96874 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 97494 477978
rect 96874 460350 97494 477922
rect 96874 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 97494 460350
rect 96874 460226 97494 460294
rect 96874 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 97494 460226
rect 96874 460102 97494 460170
rect 96874 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 97494 460102
rect 96874 459978 97494 460046
rect 96874 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 97494 459978
rect 96874 442350 97494 459922
rect 96874 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 97494 442350
rect 96874 442226 97494 442294
rect 96874 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 97494 442226
rect 96874 442102 97494 442170
rect 96874 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 97494 442102
rect 96874 441978 97494 442046
rect 96874 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 97494 441978
rect 96874 424350 97494 441922
rect 96874 424294 96970 424350
rect 97026 424294 97094 424350
rect 97150 424294 97218 424350
rect 97274 424294 97342 424350
rect 97398 424294 97494 424350
rect 96874 424226 97494 424294
rect 96874 424170 96970 424226
rect 97026 424170 97094 424226
rect 97150 424170 97218 424226
rect 97274 424170 97342 424226
rect 97398 424170 97494 424226
rect 96874 424102 97494 424170
rect 96874 424046 96970 424102
rect 97026 424046 97094 424102
rect 97150 424046 97218 424102
rect 97274 424046 97342 424102
rect 97398 424046 97494 424102
rect 96874 423978 97494 424046
rect 96874 423922 96970 423978
rect 97026 423922 97094 423978
rect 97150 423922 97218 423978
rect 97274 423922 97342 423978
rect 97398 423922 97494 423978
rect 96874 406350 97494 423922
rect 96874 406294 96970 406350
rect 97026 406294 97094 406350
rect 97150 406294 97218 406350
rect 97274 406294 97342 406350
rect 97398 406294 97494 406350
rect 96874 406226 97494 406294
rect 96874 406170 96970 406226
rect 97026 406170 97094 406226
rect 97150 406170 97218 406226
rect 97274 406170 97342 406226
rect 97398 406170 97494 406226
rect 96874 406102 97494 406170
rect 96874 406046 96970 406102
rect 97026 406046 97094 406102
rect 97150 406046 97218 406102
rect 97274 406046 97342 406102
rect 97398 406046 97494 406102
rect 96874 405978 97494 406046
rect 96874 405922 96970 405978
rect 97026 405922 97094 405978
rect 97150 405922 97218 405978
rect 97274 405922 97342 405978
rect 97398 405922 97494 405978
rect 96874 388350 97494 405922
rect 96874 388294 96970 388350
rect 97026 388294 97094 388350
rect 97150 388294 97218 388350
rect 97274 388294 97342 388350
rect 97398 388294 97494 388350
rect 96874 388226 97494 388294
rect 96874 388170 96970 388226
rect 97026 388170 97094 388226
rect 97150 388170 97218 388226
rect 97274 388170 97342 388226
rect 97398 388170 97494 388226
rect 96874 388102 97494 388170
rect 96874 388046 96970 388102
rect 97026 388046 97094 388102
rect 97150 388046 97218 388102
rect 97274 388046 97342 388102
rect 97398 388046 97494 388102
rect 96874 387978 97494 388046
rect 96874 387922 96970 387978
rect 97026 387922 97094 387978
rect 97150 387922 97218 387978
rect 97274 387922 97342 387978
rect 97398 387922 97494 387978
rect 96874 370350 97494 387922
rect 96874 370294 96970 370350
rect 97026 370294 97094 370350
rect 97150 370294 97218 370350
rect 97274 370294 97342 370350
rect 97398 370294 97494 370350
rect 96874 370226 97494 370294
rect 96874 370170 96970 370226
rect 97026 370170 97094 370226
rect 97150 370170 97218 370226
rect 97274 370170 97342 370226
rect 97398 370170 97494 370226
rect 96874 370102 97494 370170
rect 96874 370046 96970 370102
rect 97026 370046 97094 370102
rect 97150 370046 97218 370102
rect 97274 370046 97342 370102
rect 97398 370046 97494 370102
rect 96874 369978 97494 370046
rect 96874 369922 96970 369978
rect 97026 369922 97094 369978
rect 97150 369922 97218 369978
rect 97274 369922 97342 369978
rect 97398 369922 97494 369978
rect 96874 352350 97494 369922
rect 96874 352294 96970 352350
rect 97026 352294 97094 352350
rect 97150 352294 97218 352350
rect 97274 352294 97342 352350
rect 97398 352294 97494 352350
rect 96874 352226 97494 352294
rect 96874 352170 96970 352226
rect 97026 352170 97094 352226
rect 97150 352170 97218 352226
rect 97274 352170 97342 352226
rect 97398 352170 97494 352226
rect 96874 352102 97494 352170
rect 96874 352046 96970 352102
rect 97026 352046 97094 352102
rect 97150 352046 97218 352102
rect 97274 352046 97342 352102
rect 97398 352046 97494 352102
rect 96874 351978 97494 352046
rect 96874 351922 96970 351978
rect 97026 351922 97094 351978
rect 97150 351922 97218 351978
rect 97274 351922 97342 351978
rect 97398 351922 97494 351978
rect 96874 334350 97494 351922
rect 96874 334294 96970 334350
rect 97026 334294 97094 334350
rect 97150 334294 97218 334350
rect 97274 334294 97342 334350
rect 97398 334294 97494 334350
rect 96874 334226 97494 334294
rect 96874 334170 96970 334226
rect 97026 334170 97094 334226
rect 97150 334170 97218 334226
rect 97274 334170 97342 334226
rect 97398 334170 97494 334226
rect 96874 334102 97494 334170
rect 96874 334046 96970 334102
rect 97026 334046 97094 334102
rect 97150 334046 97218 334102
rect 97274 334046 97342 334102
rect 97398 334046 97494 334102
rect 96874 333978 97494 334046
rect 96874 333922 96970 333978
rect 97026 333922 97094 333978
rect 97150 333922 97218 333978
rect 97274 333922 97342 333978
rect 97398 333922 97494 333978
rect 96874 316350 97494 333922
rect 96874 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 97494 316350
rect 96874 316226 97494 316294
rect 96874 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 97494 316226
rect 96874 316102 97494 316170
rect 96874 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 97494 316102
rect 96874 315978 97494 316046
rect 96874 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 97494 315978
rect 96874 298350 97494 315922
rect 96874 298294 96970 298350
rect 97026 298294 97094 298350
rect 97150 298294 97218 298350
rect 97274 298294 97342 298350
rect 97398 298294 97494 298350
rect 96874 298226 97494 298294
rect 96874 298170 96970 298226
rect 97026 298170 97094 298226
rect 97150 298170 97218 298226
rect 97274 298170 97342 298226
rect 97398 298170 97494 298226
rect 96874 298102 97494 298170
rect 96874 298046 96970 298102
rect 97026 298046 97094 298102
rect 97150 298046 97218 298102
rect 97274 298046 97342 298102
rect 97398 298046 97494 298102
rect 96874 297978 97494 298046
rect 96874 297922 96970 297978
rect 97026 297922 97094 297978
rect 97150 297922 97218 297978
rect 97274 297922 97342 297978
rect 97398 297922 97494 297978
rect 96874 280350 97494 297922
rect 96874 280294 96970 280350
rect 97026 280294 97094 280350
rect 97150 280294 97218 280350
rect 97274 280294 97342 280350
rect 97398 280294 97494 280350
rect 96874 280226 97494 280294
rect 96874 280170 96970 280226
rect 97026 280170 97094 280226
rect 97150 280170 97218 280226
rect 97274 280170 97342 280226
rect 97398 280170 97494 280226
rect 96874 280102 97494 280170
rect 96874 280046 96970 280102
rect 97026 280046 97094 280102
rect 97150 280046 97218 280102
rect 97274 280046 97342 280102
rect 97398 280046 97494 280102
rect 96874 279978 97494 280046
rect 96874 279922 96970 279978
rect 97026 279922 97094 279978
rect 97150 279922 97218 279978
rect 97274 279922 97342 279978
rect 97398 279922 97494 279978
rect 96874 262350 97494 279922
rect 96874 262294 96970 262350
rect 97026 262294 97094 262350
rect 97150 262294 97218 262350
rect 97274 262294 97342 262350
rect 97398 262294 97494 262350
rect 96874 262226 97494 262294
rect 96874 262170 96970 262226
rect 97026 262170 97094 262226
rect 97150 262170 97218 262226
rect 97274 262170 97342 262226
rect 97398 262170 97494 262226
rect 96874 262102 97494 262170
rect 96874 262046 96970 262102
rect 97026 262046 97094 262102
rect 97150 262046 97218 262102
rect 97274 262046 97342 262102
rect 97398 262046 97494 262102
rect 96874 261978 97494 262046
rect 96874 261922 96970 261978
rect 97026 261922 97094 261978
rect 97150 261922 97218 261978
rect 97274 261922 97342 261978
rect 97398 261922 97494 261978
rect 96874 244350 97494 261922
rect 96874 244294 96970 244350
rect 97026 244294 97094 244350
rect 97150 244294 97218 244350
rect 97274 244294 97342 244350
rect 97398 244294 97494 244350
rect 96874 244226 97494 244294
rect 96874 244170 96970 244226
rect 97026 244170 97094 244226
rect 97150 244170 97218 244226
rect 97274 244170 97342 244226
rect 97398 244170 97494 244226
rect 96874 244102 97494 244170
rect 96874 244046 96970 244102
rect 97026 244046 97094 244102
rect 97150 244046 97218 244102
rect 97274 244046 97342 244102
rect 97398 244046 97494 244102
rect 96874 243978 97494 244046
rect 96874 243922 96970 243978
rect 97026 243922 97094 243978
rect 97150 243922 97218 243978
rect 97274 243922 97342 243978
rect 97398 243922 97494 243978
rect 96874 226350 97494 243922
rect 96874 226294 96970 226350
rect 97026 226294 97094 226350
rect 97150 226294 97218 226350
rect 97274 226294 97342 226350
rect 97398 226294 97494 226350
rect 96874 226226 97494 226294
rect 96874 226170 96970 226226
rect 97026 226170 97094 226226
rect 97150 226170 97218 226226
rect 97274 226170 97342 226226
rect 97398 226170 97494 226226
rect 96874 226102 97494 226170
rect 96874 226046 96970 226102
rect 97026 226046 97094 226102
rect 97150 226046 97218 226102
rect 97274 226046 97342 226102
rect 97398 226046 97494 226102
rect 96874 225978 97494 226046
rect 96874 225922 96970 225978
rect 97026 225922 97094 225978
rect 97150 225922 97218 225978
rect 97274 225922 97342 225978
rect 97398 225922 97494 225978
rect 96874 208350 97494 225922
rect 96874 208294 96970 208350
rect 97026 208294 97094 208350
rect 97150 208294 97218 208350
rect 97274 208294 97342 208350
rect 97398 208294 97494 208350
rect 96874 208226 97494 208294
rect 96874 208170 96970 208226
rect 97026 208170 97094 208226
rect 97150 208170 97218 208226
rect 97274 208170 97342 208226
rect 97398 208170 97494 208226
rect 96874 208102 97494 208170
rect 96874 208046 96970 208102
rect 97026 208046 97094 208102
rect 97150 208046 97218 208102
rect 97274 208046 97342 208102
rect 97398 208046 97494 208102
rect 96874 207978 97494 208046
rect 96874 207922 96970 207978
rect 97026 207922 97094 207978
rect 97150 207922 97218 207978
rect 97274 207922 97342 207978
rect 97398 207922 97494 207978
rect 96874 190350 97494 207922
rect 96874 190294 96970 190350
rect 97026 190294 97094 190350
rect 97150 190294 97218 190350
rect 97274 190294 97342 190350
rect 97398 190294 97494 190350
rect 96874 190226 97494 190294
rect 96874 190170 96970 190226
rect 97026 190170 97094 190226
rect 97150 190170 97218 190226
rect 97274 190170 97342 190226
rect 97398 190170 97494 190226
rect 96874 190102 97494 190170
rect 96874 190046 96970 190102
rect 97026 190046 97094 190102
rect 97150 190046 97218 190102
rect 97274 190046 97342 190102
rect 97398 190046 97494 190102
rect 96874 189978 97494 190046
rect 96874 189922 96970 189978
rect 97026 189922 97094 189978
rect 97150 189922 97218 189978
rect 97274 189922 97342 189978
rect 97398 189922 97494 189978
rect 96874 172350 97494 189922
rect 96874 172294 96970 172350
rect 97026 172294 97094 172350
rect 97150 172294 97218 172350
rect 97274 172294 97342 172350
rect 97398 172294 97494 172350
rect 96874 172226 97494 172294
rect 96874 172170 96970 172226
rect 97026 172170 97094 172226
rect 97150 172170 97218 172226
rect 97274 172170 97342 172226
rect 97398 172170 97494 172226
rect 96874 172102 97494 172170
rect 96874 172046 96970 172102
rect 97026 172046 97094 172102
rect 97150 172046 97218 172102
rect 97274 172046 97342 172102
rect 97398 172046 97494 172102
rect 96874 171978 97494 172046
rect 96874 171922 96970 171978
rect 97026 171922 97094 171978
rect 97150 171922 97218 171978
rect 97274 171922 97342 171978
rect 97398 171922 97494 171978
rect 96874 154350 97494 171922
rect 96874 154294 96970 154350
rect 97026 154294 97094 154350
rect 97150 154294 97218 154350
rect 97274 154294 97342 154350
rect 97398 154294 97494 154350
rect 96874 154226 97494 154294
rect 96874 154170 96970 154226
rect 97026 154170 97094 154226
rect 97150 154170 97218 154226
rect 97274 154170 97342 154226
rect 97398 154170 97494 154226
rect 96874 154102 97494 154170
rect 96874 154046 96970 154102
rect 97026 154046 97094 154102
rect 97150 154046 97218 154102
rect 97274 154046 97342 154102
rect 97398 154046 97494 154102
rect 96874 153978 97494 154046
rect 96874 153922 96970 153978
rect 97026 153922 97094 153978
rect 97150 153922 97218 153978
rect 97274 153922 97342 153978
rect 97398 153922 97494 153978
rect 96874 136350 97494 153922
rect 96874 136294 96970 136350
rect 97026 136294 97094 136350
rect 97150 136294 97218 136350
rect 97274 136294 97342 136350
rect 97398 136294 97494 136350
rect 96874 136226 97494 136294
rect 96874 136170 96970 136226
rect 97026 136170 97094 136226
rect 97150 136170 97218 136226
rect 97274 136170 97342 136226
rect 97398 136170 97494 136226
rect 96874 136102 97494 136170
rect 96874 136046 96970 136102
rect 97026 136046 97094 136102
rect 97150 136046 97218 136102
rect 97274 136046 97342 136102
rect 97398 136046 97494 136102
rect 96874 135978 97494 136046
rect 96874 135922 96970 135978
rect 97026 135922 97094 135978
rect 97150 135922 97218 135978
rect 97274 135922 97342 135978
rect 97398 135922 97494 135978
rect 96874 118350 97494 135922
rect 96874 118294 96970 118350
rect 97026 118294 97094 118350
rect 97150 118294 97218 118350
rect 97274 118294 97342 118350
rect 97398 118294 97494 118350
rect 96874 118226 97494 118294
rect 96874 118170 96970 118226
rect 97026 118170 97094 118226
rect 97150 118170 97218 118226
rect 97274 118170 97342 118226
rect 97398 118170 97494 118226
rect 96874 118102 97494 118170
rect 96874 118046 96970 118102
rect 97026 118046 97094 118102
rect 97150 118046 97218 118102
rect 97274 118046 97342 118102
rect 97398 118046 97494 118102
rect 96874 117978 97494 118046
rect 96874 117922 96970 117978
rect 97026 117922 97094 117978
rect 97150 117922 97218 117978
rect 97274 117922 97342 117978
rect 97398 117922 97494 117978
rect 96874 100350 97494 117922
rect 96874 100294 96970 100350
rect 97026 100294 97094 100350
rect 97150 100294 97218 100350
rect 97274 100294 97342 100350
rect 97398 100294 97494 100350
rect 96874 100226 97494 100294
rect 96874 100170 96970 100226
rect 97026 100170 97094 100226
rect 97150 100170 97218 100226
rect 97274 100170 97342 100226
rect 97398 100170 97494 100226
rect 96874 100102 97494 100170
rect 96874 100046 96970 100102
rect 97026 100046 97094 100102
rect 97150 100046 97218 100102
rect 97274 100046 97342 100102
rect 97398 100046 97494 100102
rect 96874 99978 97494 100046
rect 96874 99922 96970 99978
rect 97026 99922 97094 99978
rect 97150 99922 97218 99978
rect 97274 99922 97342 99978
rect 97398 99922 97494 99978
rect 96874 82350 97494 99922
rect 96874 82294 96970 82350
rect 97026 82294 97094 82350
rect 97150 82294 97218 82350
rect 97274 82294 97342 82350
rect 97398 82294 97494 82350
rect 96874 82226 97494 82294
rect 96874 82170 96970 82226
rect 97026 82170 97094 82226
rect 97150 82170 97218 82226
rect 97274 82170 97342 82226
rect 97398 82170 97494 82226
rect 96874 82102 97494 82170
rect 96874 82046 96970 82102
rect 97026 82046 97094 82102
rect 97150 82046 97218 82102
rect 97274 82046 97342 82102
rect 97398 82046 97494 82102
rect 96874 81978 97494 82046
rect 96874 81922 96970 81978
rect 97026 81922 97094 81978
rect 97150 81922 97218 81978
rect 97274 81922 97342 81978
rect 97398 81922 97494 81978
rect 96874 64350 97494 81922
rect 96874 64294 96970 64350
rect 97026 64294 97094 64350
rect 97150 64294 97218 64350
rect 97274 64294 97342 64350
rect 97398 64294 97494 64350
rect 96874 64226 97494 64294
rect 96874 64170 96970 64226
rect 97026 64170 97094 64226
rect 97150 64170 97218 64226
rect 97274 64170 97342 64226
rect 97398 64170 97494 64226
rect 96874 64102 97494 64170
rect 96874 64046 96970 64102
rect 97026 64046 97094 64102
rect 97150 64046 97218 64102
rect 97274 64046 97342 64102
rect 97398 64046 97494 64102
rect 96874 63978 97494 64046
rect 96874 63922 96970 63978
rect 97026 63922 97094 63978
rect 97150 63922 97218 63978
rect 97274 63922 97342 63978
rect 97398 63922 97494 63978
rect 96874 46350 97494 63922
rect 96874 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 97494 46350
rect 96874 46226 97494 46294
rect 96874 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 97494 46226
rect 96874 46102 97494 46170
rect 96874 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 97494 46102
rect 96874 45978 97494 46046
rect 96874 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 97494 45978
rect 96874 28350 97494 45922
rect 96874 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 97494 28350
rect 96874 28226 97494 28294
rect 96874 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 97494 28226
rect 96874 28102 97494 28170
rect 96874 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 97494 28102
rect 96874 27978 97494 28046
rect 96874 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 97494 27978
rect 96874 10350 97494 27922
rect 96874 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 97494 10350
rect 96874 10226 97494 10294
rect 96874 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 97494 10226
rect 96874 10102 97494 10170
rect 96874 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 97494 10102
rect 96874 9978 97494 10046
rect 96874 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 97494 9978
rect 96874 -1120 97494 9922
rect 96874 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 97494 -1120
rect 96874 -1244 97494 -1176
rect 96874 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 97494 -1244
rect 96874 -1368 97494 -1300
rect 96874 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 97494 -1368
rect 96874 -1492 97494 -1424
rect 96874 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 97494 -1492
rect 96874 -1644 97494 -1548
rect 111154 597212 111774 598268
rect 111154 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 111774 597212
rect 111154 597088 111774 597156
rect 111154 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 111774 597088
rect 111154 596964 111774 597032
rect 111154 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 111774 596964
rect 111154 596840 111774 596908
rect 111154 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 111774 596840
rect 111154 580350 111774 596784
rect 111154 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 111774 580350
rect 111154 580226 111774 580294
rect 111154 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 111774 580226
rect 111154 580102 111774 580170
rect 111154 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 111774 580102
rect 111154 579978 111774 580046
rect 111154 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 111774 579978
rect 111154 562350 111774 579922
rect 111154 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 111774 562350
rect 111154 562226 111774 562294
rect 111154 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 111774 562226
rect 111154 562102 111774 562170
rect 111154 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 111774 562102
rect 111154 561978 111774 562046
rect 111154 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 111774 561978
rect 111154 544350 111774 561922
rect 111154 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 111774 544350
rect 111154 544226 111774 544294
rect 111154 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 111774 544226
rect 111154 544102 111774 544170
rect 111154 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 111774 544102
rect 111154 543978 111774 544046
rect 111154 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 111774 543978
rect 111154 526350 111774 543922
rect 111154 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 111774 526350
rect 111154 526226 111774 526294
rect 111154 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 111774 526226
rect 111154 526102 111774 526170
rect 111154 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 111774 526102
rect 111154 525978 111774 526046
rect 111154 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 111774 525978
rect 111154 508350 111774 525922
rect 111154 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 111774 508350
rect 111154 508226 111774 508294
rect 111154 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 111774 508226
rect 111154 508102 111774 508170
rect 111154 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 111774 508102
rect 111154 507978 111774 508046
rect 111154 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 111774 507978
rect 111154 490350 111774 507922
rect 111154 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 111774 490350
rect 111154 490226 111774 490294
rect 111154 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 111774 490226
rect 111154 490102 111774 490170
rect 111154 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 111774 490102
rect 111154 489978 111774 490046
rect 111154 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 111774 489978
rect 111154 472350 111774 489922
rect 111154 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 111774 472350
rect 111154 472226 111774 472294
rect 111154 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 111774 472226
rect 111154 472102 111774 472170
rect 111154 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 111774 472102
rect 111154 471978 111774 472046
rect 111154 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 111774 471978
rect 111154 454350 111774 471922
rect 111154 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 111774 454350
rect 111154 454226 111774 454294
rect 111154 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 111774 454226
rect 111154 454102 111774 454170
rect 111154 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 111774 454102
rect 111154 453978 111774 454046
rect 111154 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 111774 453978
rect 111154 436350 111774 453922
rect 111154 436294 111250 436350
rect 111306 436294 111374 436350
rect 111430 436294 111498 436350
rect 111554 436294 111622 436350
rect 111678 436294 111774 436350
rect 111154 436226 111774 436294
rect 111154 436170 111250 436226
rect 111306 436170 111374 436226
rect 111430 436170 111498 436226
rect 111554 436170 111622 436226
rect 111678 436170 111774 436226
rect 111154 436102 111774 436170
rect 111154 436046 111250 436102
rect 111306 436046 111374 436102
rect 111430 436046 111498 436102
rect 111554 436046 111622 436102
rect 111678 436046 111774 436102
rect 111154 435978 111774 436046
rect 111154 435922 111250 435978
rect 111306 435922 111374 435978
rect 111430 435922 111498 435978
rect 111554 435922 111622 435978
rect 111678 435922 111774 435978
rect 111154 418350 111774 435922
rect 111154 418294 111250 418350
rect 111306 418294 111374 418350
rect 111430 418294 111498 418350
rect 111554 418294 111622 418350
rect 111678 418294 111774 418350
rect 111154 418226 111774 418294
rect 111154 418170 111250 418226
rect 111306 418170 111374 418226
rect 111430 418170 111498 418226
rect 111554 418170 111622 418226
rect 111678 418170 111774 418226
rect 111154 418102 111774 418170
rect 111154 418046 111250 418102
rect 111306 418046 111374 418102
rect 111430 418046 111498 418102
rect 111554 418046 111622 418102
rect 111678 418046 111774 418102
rect 111154 417978 111774 418046
rect 111154 417922 111250 417978
rect 111306 417922 111374 417978
rect 111430 417922 111498 417978
rect 111554 417922 111622 417978
rect 111678 417922 111774 417978
rect 111154 400350 111774 417922
rect 111154 400294 111250 400350
rect 111306 400294 111374 400350
rect 111430 400294 111498 400350
rect 111554 400294 111622 400350
rect 111678 400294 111774 400350
rect 111154 400226 111774 400294
rect 111154 400170 111250 400226
rect 111306 400170 111374 400226
rect 111430 400170 111498 400226
rect 111554 400170 111622 400226
rect 111678 400170 111774 400226
rect 111154 400102 111774 400170
rect 111154 400046 111250 400102
rect 111306 400046 111374 400102
rect 111430 400046 111498 400102
rect 111554 400046 111622 400102
rect 111678 400046 111774 400102
rect 111154 399978 111774 400046
rect 111154 399922 111250 399978
rect 111306 399922 111374 399978
rect 111430 399922 111498 399978
rect 111554 399922 111622 399978
rect 111678 399922 111774 399978
rect 111154 382350 111774 399922
rect 111154 382294 111250 382350
rect 111306 382294 111374 382350
rect 111430 382294 111498 382350
rect 111554 382294 111622 382350
rect 111678 382294 111774 382350
rect 111154 382226 111774 382294
rect 111154 382170 111250 382226
rect 111306 382170 111374 382226
rect 111430 382170 111498 382226
rect 111554 382170 111622 382226
rect 111678 382170 111774 382226
rect 111154 382102 111774 382170
rect 111154 382046 111250 382102
rect 111306 382046 111374 382102
rect 111430 382046 111498 382102
rect 111554 382046 111622 382102
rect 111678 382046 111774 382102
rect 111154 381978 111774 382046
rect 111154 381922 111250 381978
rect 111306 381922 111374 381978
rect 111430 381922 111498 381978
rect 111554 381922 111622 381978
rect 111678 381922 111774 381978
rect 111154 364350 111774 381922
rect 111154 364294 111250 364350
rect 111306 364294 111374 364350
rect 111430 364294 111498 364350
rect 111554 364294 111622 364350
rect 111678 364294 111774 364350
rect 111154 364226 111774 364294
rect 111154 364170 111250 364226
rect 111306 364170 111374 364226
rect 111430 364170 111498 364226
rect 111554 364170 111622 364226
rect 111678 364170 111774 364226
rect 111154 364102 111774 364170
rect 111154 364046 111250 364102
rect 111306 364046 111374 364102
rect 111430 364046 111498 364102
rect 111554 364046 111622 364102
rect 111678 364046 111774 364102
rect 111154 363978 111774 364046
rect 111154 363922 111250 363978
rect 111306 363922 111374 363978
rect 111430 363922 111498 363978
rect 111554 363922 111622 363978
rect 111678 363922 111774 363978
rect 111154 346350 111774 363922
rect 111154 346294 111250 346350
rect 111306 346294 111374 346350
rect 111430 346294 111498 346350
rect 111554 346294 111622 346350
rect 111678 346294 111774 346350
rect 111154 346226 111774 346294
rect 111154 346170 111250 346226
rect 111306 346170 111374 346226
rect 111430 346170 111498 346226
rect 111554 346170 111622 346226
rect 111678 346170 111774 346226
rect 111154 346102 111774 346170
rect 111154 346046 111250 346102
rect 111306 346046 111374 346102
rect 111430 346046 111498 346102
rect 111554 346046 111622 346102
rect 111678 346046 111774 346102
rect 111154 345978 111774 346046
rect 111154 345922 111250 345978
rect 111306 345922 111374 345978
rect 111430 345922 111498 345978
rect 111554 345922 111622 345978
rect 111678 345922 111774 345978
rect 111154 328350 111774 345922
rect 111154 328294 111250 328350
rect 111306 328294 111374 328350
rect 111430 328294 111498 328350
rect 111554 328294 111622 328350
rect 111678 328294 111774 328350
rect 111154 328226 111774 328294
rect 111154 328170 111250 328226
rect 111306 328170 111374 328226
rect 111430 328170 111498 328226
rect 111554 328170 111622 328226
rect 111678 328170 111774 328226
rect 111154 328102 111774 328170
rect 111154 328046 111250 328102
rect 111306 328046 111374 328102
rect 111430 328046 111498 328102
rect 111554 328046 111622 328102
rect 111678 328046 111774 328102
rect 111154 327978 111774 328046
rect 111154 327922 111250 327978
rect 111306 327922 111374 327978
rect 111430 327922 111498 327978
rect 111554 327922 111622 327978
rect 111678 327922 111774 327978
rect 111154 310350 111774 327922
rect 111154 310294 111250 310350
rect 111306 310294 111374 310350
rect 111430 310294 111498 310350
rect 111554 310294 111622 310350
rect 111678 310294 111774 310350
rect 111154 310226 111774 310294
rect 111154 310170 111250 310226
rect 111306 310170 111374 310226
rect 111430 310170 111498 310226
rect 111554 310170 111622 310226
rect 111678 310170 111774 310226
rect 111154 310102 111774 310170
rect 111154 310046 111250 310102
rect 111306 310046 111374 310102
rect 111430 310046 111498 310102
rect 111554 310046 111622 310102
rect 111678 310046 111774 310102
rect 111154 309978 111774 310046
rect 111154 309922 111250 309978
rect 111306 309922 111374 309978
rect 111430 309922 111498 309978
rect 111554 309922 111622 309978
rect 111678 309922 111774 309978
rect 111154 292350 111774 309922
rect 111154 292294 111250 292350
rect 111306 292294 111374 292350
rect 111430 292294 111498 292350
rect 111554 292294 111622 292350
rect 111678 292294 111774 292350
rect 111154 292226 111774 292294
rect 111154 292170 111250 292226
rect 111306 292170 111374 292226
rect 111430 292170 111498 292226
rect 111554 292170 111622 292226
rect 111678 292170 111774 292226
rect 111154 292102 111774 292170
rect 111154 292046 111250 292102
rect 111306 292046 111374 292102
rect 111430 292046 111498 292102
rect 111554 292046 111622 292102
rect 111678 292046 111774 292102
rect 111154 291978 111774 292046
rect 111154 291922 111250 291978
rect 111306 291922 111374 291978
rect 111430 291922 111498 291978
rect 111554 291922 111622 291978
rect 111678 291922 111774 291978
rect 111154 274350 111774 291922
rect 111154 274294 111250 274350
rect 111306 274294 111374 274350
rect 111430 274294 111498 274350
rect 111554 274294 111622 274350
rect 111678 274294 111774 274350
rect 111154 274226 111774 274294
rect 111154 274170 111250 274226
rect 111306 274170 111374 274226
rect 111430 274170 111498 274226
rect 111554 274170 111622 274226
rect 111678 274170 111774 274226
rect 111154 274102 111774 274170
rect 111154 274046 111250 274102
rect 111306 274046 111374 274102
rect 111430 274046 111498 274102
rect 111554 274046 111622 274102
rect 111678 274046 111774 274102
rect 111154 273978 111774 274046
rect 111154 273922 111250 273978
rect 111306 273922 111374 273978
rect 111430 273922 111498 273978
rect 111554 273922 111622 273978
rect 111678 273922 111774 273978
rect 111154 256350 111774 273922
rect 111154 256294 111250 256350
rect 111306 256294 111374 256350
rect 111430 256294 111498 256350
rect 111554 256294 111622 256350
rect 111678 256294 111774 256350
rect 111154 256226 111774 256294
rect 111154 256170 111250 256226
rect 111306 256170 111374 256226
rect 111430 256170 111498 256226
rect 111554 256170 111622 256226
rect 111678 256170 111774 256226
rect 111154 256102 111774 256170
rect 111154 256046 111250 256102
rect 111306 256046 111374 256102
rect 111430 256046 111498 256102
rect 111554 256046 111622 256102
rect 111678 256046 111774 256102
rect 111154 255978 111774 256046
rect 111154 255922 111250 255978
rect 111306 255922 111374 255978
rect 111430 255922 111498 255978
rect 111554 255922 111622 255978
rect 111678 255922 111774 255978
rect 111154 238350 111774 255922
rect 111154 238294 111250 238350
rect 111306 238294 111374 238350
rect 111430 238294 111498 238350
rect 111554 238294 111622 238350
rect 111678 238294 111774 238350
rect 111154 238226 111774 238294
rect 111154 238170 111250 238226
rect 111306 238170 111374 238226
rect 111430 238170 111498 238226
rect 111554 238170 111622 238226
rect 111678 238170 111774 238226
rect 111154 238102 111774 238170
rect 111154 238046 111250 238102
rect 111306 238046 111374 238102
rect 111430 238046 111498 238102
rect 111554 238046 111622 238102
rect 111678 238046 111774 238102
rect 111154 237978 111774 238046
rect 111154 237922 111250 237978
rect 111306 237922 111374 237978
rect 111430 237922 111498 237978
rect 111554 237922 111622 237978
rect 111678 237922 111774 237978
rect 111154 220350 111774 237922
rect 111154 220294 111250 220350
rect 111306 220294 111374 220350
rect 111430 220294 111498 220350
rect 111554 220294 111622 220350
rect 111678 220294 111774 220350
rect 111154 220226 111774 220294
rect 111154 220170 111250 220226
rect 111306 220170 111374 220226
rect 111430 220170 111498 220226
rect 111554 220170 111622 220226
rect 111678 220170 111774 220226
rect 111154 220102 111774 220170
rect 111154 220046 111250 220102
rect 111306 220046 111374 220102
rect 111430 220046 111498 220102
rect 111554 220046 111622 220102
rect 111678 220046 111774 220102
rect 111154 219978 111774 220046
rect 111154 219922 111250 219978
rect 111306 219922 111374 219978
rect 111430 219922 111498 219978
rect 111554 219922 111622 219978
rect 111678 219922 111774 219978
rect 111154 202350 111774 219922
rect 111154 202294 111250 202350
rect 111306 202294 111374 202350
rect 111430 202294 111498 202350
rect 111554 202294 111622 202350
rect 111678 202294 111774 202350
rect 111154 202226 111774 202294
rect 111154 202170 111250 202226
rect 111306 202170 111374 202226
rect 111430 202170 111498 202226
rect 111554 202170 111622 202226
rect 111678 202170 111774 202226
rect 111154 202102 111774 202170
rect 111154 202046 111250 202102
rect 111306 202046 111374 202102
rect 111430 202046 111498 202102
rect 111554 202046 111622 202102
rect 111678 202046 111774 202102
rect 111154 201978 111774 202046
rect 111154 201922 111250 201978
rect 111306 201922 111374 201978
rect 111430 201922 111498 201978
rect 111554 201922 111622 201978
rect 111678 201922 111774 201978
rect 111154 184350 111774 201922
rect 111154 184294 111250 184350
rect 111306 184294 111374 184350
rect 111430 184294 111498 184350
rect 111554 184294 111622 184350
rect 111678 184294 111774 184350
rect 111154 184226 111774 184294
rect 111154 184170 111250 184226
rect 111306 184170 111374 184226
rect 111430 184170 111498 184226
rect 111554 184170 111622 184226
rect 111678 184170 111774 184226
rect 111154 184102 111774 184170
rect 111154 184046 111250 184102
rect 111306 184046 111374 184102
rect 111430 184046 111498 184102
rect 111554 184046 111622 184102
rect 111678 184046 111774 184102
rect 111154 183978 111774 184046
rect 111154 183922 111250 183978
rect 111306 183922 111374 183978
rect 111430 183922 111498 183978
rect 111554 183922 111622 183978
rect 111678 183922 111774 183978
rect 111154 166350 111774 183922
rect 111154 166294 111250 166350
rect 111306 166294 111374 166350
rect 111430 166294 111498 166350
rect 111554 166294 111622 166350
rect 111678 166294 111774 166350
rect 111154 166226 111774 166294
rect 111154 166170 111250 166226
rect 111306 166170 111374 166226
rect 111430 166170 111498 166226
rect 111554 166170 111622 166226
rect 111678 166170 111774 166226
rect 111154 166102 111774 166170
rect 111154 166046 111250 166102
rect 111306 166046 111374 166102
rect 111430 166046 111498 166102
rect 111554 166046 111622 166102
rect 111678 166046 111774 166102
rect 111154 165978 111774 166046
rect 111154 165922 111250 165978
rect 111306 165922 111374 165978
rect 111430 165922 111498 165978
rect 111554 165922 111622 165978
rect 111678 165922 111774 165978
rect 111154 148350 111774 165922
rect 111154 148294 111250 148350
rect 111306 148294 111374 148350
rect 111430 148294 111498 148350
rect 111554 148294 111622 148350
rect 111678 148294 111774 148350
rect 111154 148226 111774 148294
rect 111154 148170 111250 148226
rect 111306 148170 111374 148226
rect 111430 148170 111498 148226
rect 111554 148170 111622 148226
rect 111678 148170 111774 148226
rect 111154 148102 111774 148170
rect 111154 148046 111250 148102
rect 111306 148046 111374 148102
rect 111430 148046 111498 148102
rect 111554 148046 111622 148102
rect 111678 148046 111774 148102
rect 111154 147978 111774 148046
rect 111154 147922 111250 147978
rect 111306 147922 111374 147978
rect 111430 147922 111498 147978
rect 111554 147922 111622 147978
rect 111678 147922 111774 147978
rect 111154 130350 111774 147922
rect 111154 130294 111250 130350
rect 111306 130294 111374 130350
rect 111430 130294 111498 130350
rect 111554 130294 111622 130350
rect 111678 130294 111774 130350
rect 111154 130226 111774 130294
rect 111154 130170 111250 130226
rect 111306 130170 111374 130226
rect 111430 130170 111498 130226
rect 111554 130170 111622 130226
rect 111678 130170 111774 130226
rect 111154 130102 111774 130170
rect 111154 130046 111250 130102
rect 111306 130046 111374 130102
rect 111430 130046 111498 130102
rect 111554 130046 111622 130102
rect 111678 130046 111774 130102
rect 111154 129978 111774 130046
rect 111154 129922 111250 129978
rect 111306 129922 111374 129978
rect 111430 129922 111498 129978
rect 111554 129922 111622 129978
rect 111678 129922 111774 129978
rect 111154 112350 111774 129922
rect 111154 112294 111250 112350
rect 111306 112294 111374 112350
rect 111430 112294 111498 112350
rect 111554 112294 111622 112350
rect 111678 112294 111774 112350
rect 111154 112226 111774 112294
rect 111154 112170 111250 112226
rect 111306 112170 111374 112226
rect 111430 112170 111498 112226
rect 111554 112170 111622 112226
rect 111678 112170 111774 112226
rect 111154 112102 111774 112170
rect 111154 112046 111250 112102
rect 111306 112046 111374 112102
rect 111430 112046 111498 112102
rect 111554 112046 111622 112102
rect 111678 112046 111774 112102
rect 111154 111978 111774 112046
rect 111154 111922 111250 111978
rect 111306 111922 111374 111978
rect 111430 111922 111498 111978
rect 111554 111922 111622 111978
rect 111678 111922 111774 111978
rect 111154 94350 111774 111922
rect 111154 94294 111250 94350
rect 111306 94294 111374 94350
rect 111430 94294 111498 94350
rect 111554 94294 111622 94350
rect 111678 94294 111774 94350
rect 111154 94226 111774 94294
rect 111154 94170 111250 94226
rect 111306 94170 111374 94226
rect 111430 94170 111498 94226
rect 111554 94170 111622 94226
rect 111678 94170 111774 94226
rect 111154 94102 111774 94170
rect 111154 94046 111250 94102
rect 111306 94046 111374 94102
rect 111430 94046 111498 94102
rect 111554 94046 111622 94102
rect 111678 94046 111774 94102
rect 111154 93978 111774 94046
rect 111154 93922 111250 93978
rect 111306 93922 111374 93978
rect 111430 93922 111498 93978
rect 111554 93922 111622 93978
rect 111678 93922 111774 93978
rect 111154 76350 111774 93922
rect 111154 76294 111250 76350
rect 111306 76294 111374 76350
rect 111430 76294 111498 76350
rect 111554 76294 111622 76350
rect 111678 76294 111774 76350
rect 111154 76226 111774 76294
rect 111154 76170 111250 76226
rect 111306 76170 111374 76226
rect 111430 76170 111498 76226
rect 111554 76170 111622 76226
rect 111678 76170 111774 76226
rect 111154 76102 111774 76170
rect 111154 76046 111250 76102
rect 111306 76046 111374 76102
rect 111430 76046 111498 76102
rect 111554 76046 111622 76102
rect 111678 76046 111774 76102
rect 111154 75978 111774 76046
rect 111154 75922 111250 75978
rect 111306 75922 111374 75978
rect 111430 75922 111498 75978
rect 111554 75922 111622 75978
rect 111678 75922 111774 75978
rect 111154 58350 111774 75922
rect 111154 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 111774 58350
rect 111154 58226 111774 58294
rect 111154 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 111774 58226
rect 111154 58102 111774 58170
rect 111154 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 111774 58102
rect 111154 57978 111774 58046
rect 111154 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 111774 57978
rect 111154 40350 111774 57922
rect 111154 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 111774 40350
rect 111154 40226 111774 40294
rect 111154 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 111774 40226
rect 111154 40102 111774 40170
rect 111154 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 111774 40102
rect 111154 39978 111774 40046
rect 111154 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 111774 39978
rect 111154 22350 111774 39922
rect 111154 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 111774 22350
rect 111154 22226 111774 22294
rect 111154 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 111774 22226
rect 111154 22102 111774 22170
rect 111154 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 111774 22102
rect 111154 21978 111774 22046
rect 111154 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 111774 21978
rect 111154 4350 111774 21922
rect 111154 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 111774 4350
rect 111154 4226 111774 4294
rect 111154 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 111774 4226
rect 111154 4102 111774 4170
rect 111154 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 111774 4102
rect 111154 3978 111774 4046
rect 111154 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 111774 3978
rect 111154 -160 111774 3922
rect 111154 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 111774 -160
rect 111154 -284 111774 -216
rect 111154 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 111774 -284
rect 111154 -408 111774 -340
rect 111154 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 111774 -408
rect 111154 -532 111774 -464
rect 111154 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 111774 -532
rect 111154 -1644 111774 -588
rect 114874 598172 115494 598268
rect 114874 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 115494 598172
rect 114874 598048 115494 598116
rect 114874 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 115494 598048
rect 114874 597924 115494 597992
rect 114874 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 115494 597924
rect 114874 597800 115494 597868
rect 114874 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 115494 597800
rect 114874 586350 115494 597744
rect 114874 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 115494 586350
rect 114874 586226 115494 586294
rect 114874 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 115494 586226
rect 114874 586102 115494 586170
rect 114874 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 115494 586102
rect 114874 585978 115494 586046
rect 114874 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 115494 585978
rect 114874 568350 115494 585922
rect 114874 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 115494 568350
rect 114874 568226 115494 568294
rect 114874 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 115494 568226
rect 114874 568102 115494 568170
rect 114874 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 115494 568102
rect 114874 567978 115494 568046
rect 114874 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 115494 567978
rect 114874 550350 115494 567922
rect 114874 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 115494 550350
rect 114874 550226 115494 550294
rect 114874 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 115494 550226
rect 114874 550102 115494 550170
rect 114874 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 115494 550102
rect 114874 549978 115494 550046
rect 114874 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 115494 549978
rect 114874 532350 115494 549922
rect 114874 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 115494 532350
rect 114874 532226 115494 532294
rect 114874 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 115494 532226
rect 114874 532102 115494 532170
rect 114874 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 115494 532102
rect 114874 531978 115494 532046
rect 114874 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 115494 531978
rect 114874 514350 115494 531922
rect 114874 514294 114970 514350
rect 115026 514294 115094 514350
rect 115150 514294 115218 514350
rect 115274 514294 115342 514350
rect 115398 514294 115494 514350
rect 114874 514226 115494 514294
rect 114874 514170 114970 514226
rect 115026 514170 115094 514226
rect 115150 514170 115218 514226
rect 115274 514170 115342 514226
rect 115398 514170 115494 514226
rect 114874 514102 115494 514170
rect 114874 514046 114970 514102
rect 115026 514046 115094 514102
rect 115150 514046 115218 514102
rect 115274 514046 115342 514102
rect 115398 514046 115494 514102
rect 114874 513978 115494 514046
rect 114874 513922 114970 513978
rect 115026 513922 115094 513978
rect 115150 513922 115218 513978
rect 115274 513922 115342 513978
rect 115398 513922 115494 513978
rect 114874 496350 115494 513922
rect 114874 496294 114970 496350
rect 115026 496294 115094 496350
rect 115150 496294 115218 496350
rect 115274 496294 115342 496350
rect 115398 496294 115494 496350
rect 114874 496226 115494 496294
rect 114874 496170 114970 496226
rect 115026 496170 115094 496226
rect 115150 496170 115218 496226
rect 115274 496170 115342 496226
rect 115398 496170 115494 496226
rect 114874 496102 115494 496170
rect 114874 496046 114970 496102
rect 115026 496046 115094 496102
rect 115150 496046 115218 496102
rect 115274 496046 115342 496102
rect 115398 496046 115494 496102
rect 114874 495978 115494 496046
rect 114874 495922 114970 495978
rect 115026 495922 115094 495978
rect 115150 495922 115218 495978
rect 115274 495922 115342 495978
rect 115398 495922 115494 495978
rect 114874 478350 115494 495922
rect 114874 478294 114970 478350
rect 115026 478294 115094 478350
rect 115150 478294 115218 478350
rect 115274 478294 115342 478350
rect 115398 478294 115494 478350
rect 114874 478226 115494 478294
rect 114874 478170 114970 478226
rect 115026 478170 115094 478226
rect 115150 478170 115218 478226
rect 115274 478170 115342 478226
rect 115398 478170 115494 478226
rect 114874 478102 115494 478170
rect 114874 478046 114970 478102
rect 115026 478046 115094 478102
rect 115150 478046 115218 478102
rect 115274 478046 115342 478102
rect 115398 478046 115494 478102
rect 114874 477978 115494 478046
rect 114874 477922 114970 477978
rect 115026 477922 115094 477978
rect 115150 477922 115218 477978
rect 115274 477922 115342 477978
rect 115398 477922 115494 477978
rect 114874 460350 115494 477922
rect 114874 460294 114970 460350
rect 115026 460294 115094 460350
rect 115150 460294 115218 460350
rect 115274 460294 115342 460350
rect 115398 460294 115494 460350
rect 114874 460226 115494 460294
rect 114874 460170 114970 460226
rect 115026 460170 115094 460226
rect 115150 460170 115218 460226
rect 115274 460170 115342 460226
rect 115398 460170 115494 460226
rect 114874 460102 115494 460170
rect 114874 460046 114970 460102
rect 115026 460046 115094 460102
rect 115150 460046 115218 460102
rect 115274 460046 115342 460102
rect 115398 460046 115494 460102
rect 114874 459978 115494 460046
rect 114874 459922 114970 459978
rect 115026 459922 115094 459978
rect 115150 459922 115218 459978
rect 115274 459922 115342 459978
rect 115398 459922 115494 459978
rect 114874 442350 115494 459922
rect 114874 442294 114970 442350
rect 115026 442294 115094 442350
rect 115150 442294 115218 442350
rect 115274 442294 115342 442350
rect 115398 442294 115494 442350
rect 114874 442226 115494 442294
rect 114874 442170 114970 442226
rect 115026 442170 115094 442226
rect 115150 442170 115218 442226
rect 115274 442170 115342 442226
rect 115398 442170 115494 442226
rect 114874 442102 115494 442170
rect 114874 442046 114970 442102
rect 115026 442046 115094 442102
rect 115150 442046 115218 442102
rect 115274 442046 115342 442102
rect 115398 442046 115494 442102
rect 114874 441978 115494 442046
rect 114874 441922 114970 441978
rect 115026 441922 115094 441978
rect 115150 441922 115218 441978
rect 115274 441922 115342 441978
rect 115398 441922 115494 441978
rect 114874 424350 115494 441922
rect 114874 424294 114970 424350
rect 115026 424294 115094 424350
rect 115150 424294 115218 424350
rect 115274 424294 115342 424350
rect 115398 424294 115494 424350
rect 114874 424226 115494 424294
rect 114874 424170 114970 424226
rect 115026 424170 115094 424226
rect 115150 424170 115218 424226
rect 115274 424170 115342 424226
rect 115398 424170 115494 424226
rect 114874 424102 115494 424170
rect 114874 424046 114970 424102
rect 115026 424046 115094 424102
rect 115150 424046 115218 424102
rect 115274 424046 115342 424102
rect 115398 424046 115494 424102
rect 114874 423978 115494 424046
rect 114874 423922 114970 423978
rect 115026 423922 115094 423978
rect 115150 423922 115218 423978
rect 115274 423922 115342 423978
rect 115398 423922 115494 423978
rect 114874 406350 115494 423922
rect 114874 406294 114970 406350
rect 115026 406294 115094 406350
rect 115150 406294 115218 406350
rect 115274 406294 115342 406350
rect 115398 406294 115494 406350
rect 114874 406226 115494 406294
rect 114874 406170 114970 406226
rect 115026 406170 115094 406226
rect 115150 406170 115218 406226
rect 115274 406170 115342 406226
rect 115398 406170 115494 406226
rect 114874 406102 115494 406170
rect 114874 406046 114970 406102
rect 115026 406046 115094 406102
rect 115150 406046 115218 406102
rect 115274 406046 115342 406102
rect 115398 406046 115494 406102
rect 114874 405978 115494 406046
rect 114874 405922 114970 405978
rect 115026 405922 115094 405978
rect 115150 405922 115218 405978
rect 115274 405922 115342 405978
rect 115398 405922 115494 405978
rect 114874 388350 115494 405922
rect 114874 388294 114970 388350
rect 115026 388294 115094 388350
rect 115150 388294 115218 388350
rect 115274 388294 115342 388350
rect 115398 388294 115494 388350
rect 114874 388226 115494 388294
rect 114874 388170 114970 388226
rect 115026 388170 115094 388226
rect 115150 388170 115218 388226
rect 115274 388170 115342 388226
rect 115398 388170 115494 388226
rect 114874 388102 115494 388170
rect 114874 388046 114970 388102
rect 115026 388046 115094 388102
rect 115150 388046 115218 388102
rect 115274 388046 115342 388102
rect 115398 388046 115494 388102
rect 114874 387978 115494 388046
rect 114874 387922 114970 387978
rect 115026 387922 115094 387978
rect 115150 387922 115218 387978
rect 115274 387922 115342 387978
rect 115398 387922 115494 387978
rect 114874 370350 115494 387922
rect 114874 370294 114970 370350
rect 115026 370294 115094 370350
rect 115150 370294 115218 370350
rect 115274 370294 115342 370350
rect 115398 370294 115494 370350
rect 114874 370226 115494 370294
rect 114874 370170 114970 370226
rect 115026 370170 115094 370226
rect 115150 370170 115218 370226
rect 115274 370170 115342 370226
rect 115398 370170 115494 370226
rect 114874 370102 115494 370170
rect 114874 370046 114970 370102
rect 115026 370046 115094 370102
rect 115150 370046 115218 370102
rect 115274 370046 115342 370102
rect 115398 370046 115494 370102
rect 114874 369978 115494 370046
rect 114874 369922 114970 369978
rect 115026 369922 115094 369978
rect 115150 369922 115218 369978
rect 115274 369922 115342 369978
rect 115398 369922 115494 369978
rect 114874 352350 115494 369922
rect 114874 352294 114970 352350
rect 115026 352294 115094 352350
rect 115150 352294 115218 352350
rect 115274 352294 115342 352350
rect 115398 352294 115494 352350
rect 114874 352226 115494 352294
rect 114874 352170 114970 352226
rect 115026 352170 115094 352226
rect 115150 352170 115218 352226
rect 115274 352170 115342 352226
rect 115398 352170 115494 352226
rect 114874 352102 115494 352170
rect 114874 352046 114970 352102
rect 115026 352046 115094 352102
rect 115150 352046 115218 352102
rect 115274 352046 115342 352102
rect 115398 352046 115494 352102
rect 114874 351978 115494 352046
rect 114874 351922 114970 351978
rect 115026 351922 115094 351978
rect 115150 351922 115218 351978
rect 115274 351922 115342 351978
rect 115398 351922 115494 351978
rect 114874 334350 115494 351922
rect 114874 334294 114970 334350
rect 115026 334294 115094 334350
rect 115150 334294 115218 334350
rect 115274 334294 115342 334350
rect 115398 334294 115494 334350
rect 114874 334226 115494 334294
rect 114874 334170 114970 334226
rect 115026 334170 115094 334226
rect 115150 334170 115218 334226
rect 115274 334170 115342 334226
rect 115398 334170 115494 334226
rect 114874 334102 115494 334170
rect 114874 334046 114970 334102
rect 115026 334046 115094 334102
rect 115150 334046 115218 334102
rect 115274 334046 115342 334102
rect 115398 334046 115494 334102
rect 114874 333978 115494 334046
rect 114874 333922 114970 333978
rect 115026 333922 115094 333978
rect 115150 333922 115218 333978
rect 115274 333922 115342 333978
rect 115398 333922 115494 333978
rect 114874 316350 115494 333922
rect 114874 316294 114970 316350
rect 115026 316294 115094 316350
rect 115150 316294 115218 316350
rect 115274 316294 115342 316350
rect 115398 316294 115494 316350
rect 114874 316226 115494 316294
rect 114874 316170 114970 316226
rect 115026 316170 115094 316226
rect 115150 316170 115218 316226
rect 115274 316170 115342 316226
rect 115398 316170 115494 316226
rect 114874 316102 115494 316170
rect 114874 316046 114970 316102
rect 115026 316046 115094 316102
rect 115150 316046 115218 316102
rect 115274 316046 115342 316102
rect 115398 316046 115494 316102
rect 114874 315978 115494 316046
rect 114874 315922 114970 315978
rect 115026 315922 115094 315978
rect 115150 315922 115218 315978
rect 115274 315922 115342 315978
rect 115398 315922 115494 315978
rect 114874 298350 115494 315922
rect 114874 298294 114970 298350
rect 115026 298294 115094 298350
rect 115150 298294 115218 298350
rect 115274 298294 115342 298350
rect 115398 298294 115494 298350
rect 114874 298226 115494 298294
rect 114874 298170 114970 298226
rect 115026 298170 115094 298226
rect 115150 298170 115218 298226
rect 115274 298170 115342 298226
rect 115398 298170 115494 298226
rect 114874 298102 115494 298170
rect 114874 298046 114970 298102
rect 115026 298046 115094 298102
rect 115150 298046 115218 298102
rect 115274 298046 115342 298102
rect 115398 298046 115494 298102
rect 114874 297978 115494 298046
rect 114874 297922 114970 297978
rect 115026 297922 115094 297978
rect 115150 297922 115218 297978
rect 115274 297922 115342 297978
rect 115398 297922 115494 297978
rect 114874 280350 115494 297922
rect 114874 280294 114970 280350
rect 115026 280294 115094 280350
rect 115150 280294 115218 280350
rect 115274 280294 115342 280350
rect 115398 280294 115494 280350
rect 114874 280226 115494 280294
rect 114874 280170 114970 280226
rect 115026 280170 115094 280226
rect 115150 280170 115218 280226
rect 115274 280170 115342 280226
rect 115398 280170 115494 280226
rect 114874 280102 115494 280170
rect 114874 280046 114970 280102
rect 115026 280046 115094 280102
rect 115150 280046 115218 280102
rect 115274 280046 115342 280102
rect 115398 280046 115494 280102
rect 114874 279978 115494 280046
rect 114874 279922 114970 279978
rect 115026 279922 115094 279978
rect 115150 279922 115218 279978
rect 115274 279922 115342 279978
rect 115398 279922 115494 279978
rect 114874 262350 115494 279922
rect 114874 262294 114970 262350
rect 115026 262294 115094 262350
rect 115150 262294 115218 262350
rect 115274 262294 115342 262350
rect 115398 262294 115494 262350
rect 114874 262226 115494 262294
rect 114874 262170 114970 262226
rect 115026 262170 115094 262226
rect 115150 262170 115218 262226
rect 115274 262170 115342 262226
rect 115398 262170 115494 262226
rect 114874 262102 115494 262170
rect 114874 262046 114970 262102
rect 115026 262046 115094 262102
rect 115150 262046 115218 262102
rect 115274 262046 115342 262102
rect 115398 262046 115494 262102
rect 114874 261978 115494 262046
rect 114874 261922 114970 261978
rect 115026 261922 115094 261978
rect 115150 261922 115218 261978
rect 115274 261922 115342 261978
rect 115398 261922 115494 261978
rect 114874 244350 115494 261922
rect 114874 244294 114970 244350
rect 115026 244294 115094 244350
rect 115150 244294 115218 244350
rect 115274 244294 115342 244350
rect 115398 244294 115494 244350
rect 114874 244226 115494 244294
rect 114874 244170 114970 244226
rect 115026 244170 115094 244226
rect 115150 244170 115218 244226
rect 115274 244170 115342 244226
rect 115398 244170 115494 244226
rect 114874 244102 115494 244170
rect 114874 244046 114970 244102
rect 115026 244046 115094 244102
rect 115150 244046 115218 244102
rect 115274 244046 115342 244102
rect 115398 244046 115494 244102
rect 114874 243978 115494 244046
rect 114874 243922 114970 243978
rect 115026 243922 115094 243978
rect 115150 243922 115218 243978
rect 115274 243922 115342 243978
rect 115398 243922 115494 243978
rect 114874 226350 115494 243922
rect 114874 226294 114970 226350
rect 115026 226294 115094 226350
rect 115150 226294 115218 226350
rect 115274 226294 115342 226350
rect 115398 226294 115494 226350
rect 114874 226226 115494 226294
rect 114874 226170 114970 226226
rect 115026 226170 115094 226226
rect 115150 226170 115218 226226
rect 115274 226170 115342 226226
rect 115398 226170 115494 226226
rect 114874 226102 115494 226170
rect 114874 226046 114970 226102
rect 115026 226046 115094 226102
rect 115150 226046 115218 226102
rect 115274 226046 115342 226102
rect 115398 226046 115494 226102
rect 114874 225978 115494 226046
rect 114874 225922 114970 225978
rect 115026 225922 115094 225978
rect 115150 225922 115218 225978
rect 115274 225922 115342 225978
rect 115398 225922 115494 225978
rect 114874 208350 115494 225922
rect 114874 208294 114970 208350
rect 115026 208294 115094 208350
rect 115150 208294 115218 208350
rect 115274 208294 115342 208350
rect 115398 208294 115494 208350
rect 114874 208226 115494 208294
rect 114874 208170 114970 208226
rect 115026 208170 115094 208226
rect 115150 208170 115218 208226
rect 115274 208170 115342 208226
rect 115398 208170 115494 208226
rect 114874 208102 115494 208170
rect 114874 208046 114970 208102
rect 115026 208046 115094 208102
rect 115150 208046 115218 208102
rect 115274 208046 115342 208102
rect 115398 208046 115494 208102
rect 114874 207978 115494 208046
rect 114874 207922 114970 207978
rect 115026 207922 115094 207978
rect 115150 207922 115218 207978
rect 115274 207922 115342 207978
rect 115398 207922 115494 207978
rect 114874 190350 115494 207922
rect 114874 190294 114970 190350
rect 115026 190294 115094 190350
rect 115150 190294 115218 190350
rect 115274 190294 115342 190350
rect 115398 190294 115494 190350
rect 114874 190226 115494 190294
rect 114874 190170 114970 190226
rect 115026 190170 115094 190226
rect 115150 190170 115218 190226
rect 115274 190170 115342 190226
rect 115398 190170 115494 190226
rect 114874 190102 115494 190170
rect 114874 190046 114970 190102
rect 115026 190046 115094 190102
rect 115150 190046 115218 190102
rect 115274 190046 115342 190102
rect 115398 190046 115494 190102
rect 114874 189978 115494 190046
rect 114874 189922 114970 189978
rect 115026 189922 115094 189978
rect 115150 189922 115218 189978
rect 115274 189922 115342 189978
rect 115398 189922 115494 189978
rect 114874 172350 115494 189922
rect 114874 172294 114970 172350
rect 115026 172294 115094 172350
rect 115150 172294 115218 172350
rect 115274 172294 115342 172350
rect 115398 172294 115494 172350
rect 114874 172226 115494 172294
rect 114874 172170 114970 172226
rect 115026 172170 115094 172226
rect 115150 172170 115218 172226
rect 115274 172170 115342 172226
rect 115398 172170 115494 172226
rect 114874 172102 115494 172170
rect 114874 172046 114970 172102
rect 115026 172046 115094 172102
rect 115150 172046 115218 172102
rect 115274 172046 115342 172102
rect 115398 172046 115494 172102
rect 114874 171978 115494 172046
rect 114874 171922 114970 171978
rect 115026 171922 115094 171978
rect 115150 171922 115218 171978
rect 115274 171922 115342 171978
rect 115398 171922 115494 171978
rect 114874 154350 115494 171922
rect 114874 154294 114970 154350
rect 115026 154294 115094 154350
rect 115150 154294 115218 154350
rect 115274 154294 115342 154350
rect 115398 154294 115494 154350
rect 114874 154226 115494 154294
rect 114874 154170 114970 154226
rect 115026 154170 115094 154226
rect 115150 154170 115218 154226
rect 115274 154170 115342 154226
rect 115398 154170 115494 154226
rect 114874 154102 115494 154170
rect 114874 154046 114970 154102
rect 115026 154046 115094 154102
rect 115150 154046 115218 154102
rect 115274 154046 115342 154102
rect 115398 154046 115494 154102
rect 114874 153978 115494 154046
rect 114874 153922 114970 153978
rect 115026 153922 115094 153978
rect 115150 153922 115218 153978
rect 115274 153922 115342 153978
rect 115398 153922 115494 153978
rect 114874 136350 115494 153922
rect 114874 136294 114970 136350
rect 115026 136294 115094 136350
rect 115150 136294 115218 136350
rect 115274 136294 115342 136350
rect 115398 136294 115494 136350
rect 114874 136226 115494 136294
rect 114874 136170 114970 136226
rect 115026 136170 115094 136226
rect 115150 136170 115218 136226
rect 115274 136170 115342 136226
rect 115398 136170 115494 136226
rect 114874 136102 115494 136170
rect 114874 136046 114970 136102
rect 115026 136046 115094 136102
rect 115150 136046 115218 136102
rect 115274 136046 115342 136102
rect 115398 136046 115494 136102
rect 114874 135978 115494 136046
rect 114874 135922 114970 135978
rect 115026 135922 115094 135978
rect 115150 135922 115218 135978
rect 115274 135922 115342 135978
rect 115398 135922 115494 135978
rect 114874 118350 115494 135922
rect 114874 118294 114970 118350
rect 115026 118294 115094 118350
rect 115150 118294 115218 118350
rect 115274 118294 115342 118350
rect 115398 118294 115494 118350
rect 114874 118226 115494 118294
rect 114874 118170 114970 118226
rect 115026 118170 115094 118226
rect 115150 118170 115218 118226
rect 115274 118170 115342 118226
rect 115398 118170 115494 118226
rect 114874 118102 115494 118170
rect 114874 118046 114970 118102
rect 115026 118046 115094 118102
rect 115150 118046 115218 118102
rect 115274 118046 115342 118102
rect 115398 118046 115494 118102
rect 114874 117978 115494 118046
rect 114874 117922 114970 117978
rect 115026 117922 115094 117978
rect 115150 117922 115218 117978
rect 115274 117922 115342 117978
rect 115398 117922 115494 117978
rect 114874 100350 115494 117922
rect 114874 100294 114970 100350
rect 115026 100294 115094 100350
rect 115150 100294 115218 100350
rect 115274 100294 115342 100350
rect 115398 100294 115494 100350
rect 114874 100226 115494 100294
rect 114874 100170 114970 100226
rect 115026 100170 115094 100226
rect 115150 100170 115218 100226
rect 115274 100170 115342 100226
rect 115398 100170 115494 100226
rect 114874 100102 115494 100170
rect 114874 100046 114970 100102
rect 115026 100046 115094 100102
rect 115150 100046 115218 100102
rect 115274 100046 115342 100102
rect 115398 100046 115494 100102
rect 114874 99978 115494 100046
rect 114874 99922 114970 99978
rect 115026 99922 115094 99978
rect 115150 99922 115218 99978
rect 115274 99922 115342 99978
rect 115398 99922 115494 99978
rect 114874 82350 115494 99922
rect 114874 82294 114970 82350
rect 115026 82294 115094 82350
rect 115150 82294 115218 82350
rect 115274 82294 115342 82350
rect 115398 82294 115494 82350
rect 114874 82226 115494 82294
rect 114874 82170 114970 82226
rect 115026 82170 115094 82226
rect 115150 82170 115218 82226
rect 115274 82170 115342 82226
rect 115398 82170 115494 82226
rect 114874 82102 115494 82170
rect 114874 82046 114970 82102
rect 115026 82046 115094 82102
rect 115150 82046 115218 82102
rect 115274 82046 115342 82102
rect 115398 82046 115494 82102
rect 114874 81978 115494 82046
rect 114874 81922 114970 81978
rect 115026 81922 115094 81978
rect 115150 81922 115218 81978
rect 115274 81922 115342 81978
rect 115398 81922 115494 81978
rect 114874 64350 115494 81922
rect 114874 64294 114970 64350
rect 115026 64294 115094 64350
rect 115150 64294 115218 64350
rect 115274 64294 115342 64350
rect 115398 64294 115494 64350
rect 114874 64226 115494 64294
rect 114874 64170 114970 64226
rect 115026 64170 115094 64226
rect 115150 64170 115218 64226
rect 115274 64170 115342 64226
rect 115398 64170 115494 64226
rect 114874 64102 115494 64170
rect 114874 64046 114970 64102
rect 115026 64046 115094 64102
rect 115150 64046 115218 64102
rect 115274 64046 115342 64102
rect 115398 64046 115494 64102
rect 114874 63978 115494 64046
rect 114874 63922 114970 63978
rect 115026 63922 115094 63978
rect 115150 63922 115218 63978
rect 115274 63922 115342 63978
rect 115398 63922 115494 63978
rect 114874 46350 115494 63922
rect 114874 46294 114970 46350
rect 115026 46294 115094 46350
rect 115150 46294 115218 46350
rect 115274 46294 115342 46350
rect 115398 46294 115494 46350
rect 114874 46226 115494 46294
rect 114874 46170 114970 46226
rect 115026 46170 115094 46226
rect 115150 46170 115218 46226
rect 115274 46170 115342 46226
rect 115398 46170 115494 46226
rect 114874 46102 115494 46170
rect 114874 46046 114970 46102
rect 115026 46046 115094 46102
rect 115150 46046 115218 46102
rect 115274 46046 115342 46102
rect 115398 46046 115494 46102
rect 114874 45978 115494 46046
rect 114874 45922 114970 45978
rect 115026 45922 115094 45978
rect 115150 45922 115218 45978
rect 115274 45922 115342 45978
rect 115398 45922 115494 45978
rect 114874 28350 115494 45922
rect 114874 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 115494 28350
rect 114874 28226 115494 28294
rect 114874 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 115494 28226
rect 114874 28102 115494 28170
rect 114874 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 115494 28102
rect 114874 27978 115494 28046
rect 114874 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 115494 27978
rect 114874 10350 115494 27922
rect 114874 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 115494 10350
rect 114874 10226 115494 10294
rect 114874 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 115494 10226
rect 114874 10102 115494 10170
rect 114874 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 115494 10102
rect 114874 9978 115494 10046
rect 114874 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 115494 9978
rect 114874 -1120 115494 9922
rect 114874 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 115494 -1120
rect 114874 -1244 115494 -1176
rect 114874 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 115494 -1244
rect 114874 -1368 115494 -1300
rect 114874 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 115494 -1368
rect 114874 -1492 115494 -1424
rect 114874 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 115494 -1492
rect 114874 -1644 115494 -1548
rect 129154 597212 129774 598268
rect 129154 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 129774 597212
rect 129154 597088 129774 597156
rect 129154 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 129774 597088
rect 129154 596964 129774 597032
rect 129154 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 129774 596964
rect 129154 596840 129774 596908
rect 129154 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 129774 596840
rect 129154 580350 129774 596784
rect 129154 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 129774 580350
rect 129154 580226 129774 580294
rect 129154 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 129774 580226
rect 129154 580102 129774 580170
rect 129154 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 129774 580102
rect 129154 579978 129774 580046
rect 129154 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 129774 579978
rect 129154 562350 129774 579922
rect 129154 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 129774 562350
rect 129154 562226 129774 562294
rect 129154 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 129774 562226
rect 129154 562102 129774 562170
rect 129154 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 129774 562102
rect 129154 561978 129774 562046
rect 129154 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 129774 561978
rect 129154 544350 129774 561922
rect 129154 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 129774 544350
rect 129154 544226 129774 544294
rect 129154 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 129774 544226
rect 129154 544102 129774 544170
rect 129154 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 129774 544102
rect 129154 543978 129774 544046
rect 129154 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 129774 543978
rect 129154 526350 129774 543922
rect 129154 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 129774 526350
rect 129154 526226 129774 526294
rect 129154 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 129774 526226
rect 129154 526102 129774 526170
rect 129154 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 129774 526102
rect 129154 525978 129774 526046
rect 129154 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 129774 525978
rect 129154 508350 129774 525922
rect 129154 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 129774 508350
rect 129154 508226 129774 508294
rect 129154 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 129774 508226
rect 129154 508102 129774 508170
rect 129154 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 129774 508102
rect 129154 507978 129774 508046
rect 129154 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 129774 507978
rect 129154 490350 129774 507922
rect 129154 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 129774 490350
rect 129154 490226 129774 490294
rect 129154 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 129774 490226
rect 129154 490102 129774 490170
rect 129154 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 129774 490102
rect 129154 489978 129774 490046
rect 129154 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 129774 489978
rect 129154 472350 129774 489922
rect 129154 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 129774 472350
rect 129154 472226 129774 472294
rect 129154 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 129774 472226
rect 129154 472102 129774 472170
rect 129154 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 129774 472102
rect 129154 471978 129774 472046
rect 129154 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 129774 471978
rect 129154 454350 129774 471922
rect 129154 454294 129250 454350
rect 129306 454294 129374 454350
rect 129430 454294 129498 454350
rect 129554 454294 129622 454350
rect 129678 454294 129774 454350
rect 129154 454226 129774 454294
rect 129154 454170 129250 454226
rect 129306 454170 129374 454226
rect 129430 454170 129498 454226
rect 129554 454170 129622 454226
rect 129678 454170 129774 454226
rect 129154 454102 129774 454170
rect 129154 454046 129250 454102
rect 129306 454046 129374 454102
rect 129430 454046 129498 454102
rect 129554 454046 129622 454102
rect 129678 454046 129774 454102
rect 129154 453978 129774 454046
rect 129154 453922 129250 453978
rect 129306 453922 129374 453978
rect 129430 453922 129498 453978
rect 129554 453922 129622 453978
rect 129678 453922 129774 453978
rect 129154 436350 129774 453922
rect 129154 436294 129250 436350
rect 129306 436294 129374 436350
rect 129430 436294 129498 436350
rect 129554 436294 129622 436350
rect 129678 436294 129774 436350
rect 129154 436226 129774 436294
rect 129154 436170 129250 436226
rect 129306 436170 129374 436226
rect 129430 436170 129498 436226
rect 129554 436170 129622 436226
rect 129678 436170 129774 436226
rect 129154 436102 129774 436170
rect 129154 436046 129250 436102
rect 129306 436046 129374 436102
rect 129430 436046 129498 436102
rect 129554 436046 129622 436102
rect 129678 436046 129774 436102
rect 129154 435978 129774 436046
rect 129154 435922 129250 435978
rect 129306 435922 129374 435978
rect 129430 435922 129498 435978
rect 129554 435922 129622 435978
rect 129678 435922 129774 435978
rect 129154 418350 129774 435922
rect 129154 418294 129250 418350
rect 129306 418294 129374 418350
rect 129430 418294 129498 418350
rect 129554 418294 129622 418350
rect 129678 418294 129774 418350
rect 129154 418226 129774 418294
rect 129154 418170 129250 418226
rect 129306 418170 129374 418226
rect 129430 418170 129498 418226
rect 129554 418170 129622 418226
rect 129678 418170 129774 418226
rect 129154 418102 129774 418170
rect 129154 418046 129250 418102
rect 129306 418046 129374 418102
rect 129430 418046 129498 418102
rect 129554 418046 129622 418102
rect 129678 418046 129774 418102
rect 129154 417978 129774 418046
rect 129154 417922 129250 417978
rect 129306 417922 129374 417978
rect 129430 417922 129498 417978
rect 129554 417922 129622 417978
rect 129678 417922 129774 417978
rect 129154 400350 129774 417922
rect 129154 400294 129250 400350
rect 129306 400294 129374 400350
rect 129430 400294 129498 400350
rect 129554 400294 129622 400350
rect 129678 400294 129774 400350
rect 129154 400226 129774 400294
rect 129154 400170 129250 400226
rect 129306 400170 129374 400226
rect 129430 400170 129498 400226
rect 129554 400170 129622 400226
rect 129678 400170 129774 400226
rect 129154 400102 129774 400170
rect 129154 400046 129250 400102
rect 129306 400046 129374 400102
rect 129430 400046 129498 400102
rect 129554 400046 129622 400102
rect 129678 400046 129774 400102
rect 129154 399978 129774 400046
rect 129154 399922 129250 399978
rect 129306 399922 129374 399978
rect 129430 399922 129498 399978
rect 129554 399922 129622 399978
rect 129678 399922 129774 399978
rect 129154 382350 129774 399922
rect 129154 382294 129250 382350
rect 129306 382294 129374 382350
rect 129430 382294 129498 382350
rect 129554 382294 129622 382350
rect 129678 382294 129774 382350
rect 129154 382226 129774 382294
rect 129154 382170 129250 382226
rect 129306 382170 129374 382226
rect 129430 382170 129498 382226
rect 129554 382170 129622 382226
rect 129678 382170 129774 382226
rect 129154 382102 129774 382170
rect 129154 382046 129250 382102
rect 129306 382046 129374 382102
rect 129430 382046 129498 382102
rect 129554 382046 129622 382102
rect 129678 382046 129774 382102
rect 129154 381978 129774 382046
rect 129154 381922 129250 381978
rect 129306 381922 129374 381978
rect 129430 381922 129498 381978
rect 129554 381922 129622 381978
rect 129678 381922 129774 381978
rect 129154 364350 129774 381922
rect 129154 364294 129250 364350
rect 129306 364294 129374 364350
rect 129430 364294 129498 364350
rect 129554 364294 129622 364350
rect 129678 364294 129774 364350
rect 129154 364226 129774 364294
rect 129154 364170 129250 364226
rect 129306 364170 129374 364226
rect 129430 364170 129498 364226
rect 129554 364170 129622 364226
rect 129678 364170 129774 364226
rect 129154 364102 129774 364170
rect 129154 364046 129250 364102
rect 129306 364046 129374 364102
rect 129430 364046 129498 364102
rect 129554 364046 129622 364102
rect 129678 364046 129774 364102
rect 129154 363978 129774 364046
rect 129154 363922 129250 363978
rect 129306 363922 129374 363978
rect 129430 363922 129498 363978
rect 129554 363922 129622 363978
rect 129678 363922 129774 363978
rect 129154 346350 129774 363922
rect 129154 346294 129250 346350
rect 129306 346294 129374 346350
rect 129430 346294 129498 346350
rect 129554 346294 129622 346350
rect 129678 346294 129774 346350
rect 129154 346226 129774 346294
rect 129154 346170 129250 346226
rect 129306 346170 129374 346226
rect 129430 346170 129498 346226
rect 129554 346170 129622 346226
rect 129678 346170 129774 346226
rect 129154 346102 129774 346170
rect 129154 346046 129250 346102
rect 129306 346046 129374 346102
rect 129430 346046 129498 346102
rect 129554 346046 129622 346102
rect 129678 346046 129774 346102
rect 129154 345978 129774 346046
rect 129154 345922 129250 345978
rect 129306 345922 129374 345978
rect 129430 345922 129498 345978
rect 129554 345922 129622 345978
rect 129678 345922 129774 345978
rect 129154 328350 129774 345922
rect 129154 328294 129250 328350
rect 129306 328294 129374 328350
rect 129430 328294 129498 328350
rect 129554 328294 129622 328350
rect 129678 328294 129774 328350
rect 129154 328226 129774 328294
rect 129154 328170 129250 328226
rect 129306 328170 129374 328226
rect 129430 328170 129498 328226
rect 129554 328170 129622 328226
rect 129678 328170 129774 328226
rect 129154 328102 129774 328170
rect 129154 328046 129250 328102
rect 129306 328046 129374 328102
rect 129430 328046 129498 328102
rect 129554 328046 129622 328102
rect 129678 328046 129774 328102
rect 129154 327978 129774 328046
rect 129154 327922 129250 327978
rect 129306 327922 129374 327978
rect 129430 327922 129498 327978
rect 129554 327922 129622 327978
rect 129678 327922 129774 327978
rect 129154 310350 129774 327922
rect 129154 310294 129250 310350
rect 129306 310294 129374 310350
rect 129430 310294 129498 310350
rect 129554 310294 129622 310350
rect 129678 310294 129774 310350
rect 129154 310226 129774 310294
rect 129154 310170 129250 310226
rect 129306 310170 129374 310226
rect 129430 310170 129498 310226
rect 129554 310170 129622 310226
rect 129678 310170 129774 310226
rect 129154 310102 129774 310170
rect 129154 310046 129250 310102
rect 129306 310046 129374 310102
rect 129430 310046 129498 310102
rect 129554 310046 129622 310102
rect 129678 310046 129774 310102
rect 129154 309978 129774 310046
rect 129154 309922 129250 309978
rect 129306 309922 129374 309978
rect 129430 309922 129498 309978
rect 129554 309922 129622 309978
rect 129678 309922 129774 309978
rect 129154 292350 129774 309922
rect 129154 292294 129250 292350
rect 129306 292294 129374 292350
rect 129430 292294 129498 292350
rect 129554 292294 129622 292350
rect 129678 292294 129774 292350
rect 129154 292226 129774 292294
rect 129154 292170 129250 292226
rect 129306 292170 129374 292226
rect 129430 292170 129498 292226
rect 129554 292170 129622 292226
rect 129678 292170 129774 292226
rect 129154 292102 129774 292170
rect 129154 292046 129250 292102
rect 129306 292046 129374 292102
rect 129430 292046 129498 292102
rect 129554 292046 129622 292102
rect 129678 292046 129774 292102
rect 129154 291978 129774 292046
rect 129154 291922 129250 291978
rect 129306 291922 129374 291978
rect 129430 291922 129498 291978
rect 129554 291922 129622 291978
rect 129678 291922 129774 291978
rect 129154 274350 129774 291922
rect 129154 274294 129250 274350
rect 129306 274294 129374 274350
rect 129430 274294 129498 274350
rect 129554 274294 129622 274350
rect 129678 274294 129774 274350
rect 129154 274226 129774 274294
rect 129154 274170 129250 274226
rect 129306 274170 129374 274226
rect 129430 274170 129498 274226
rect 129554 274170 129622 274226
rect 129678 274170 129774 274226
rect 129154 274102 129774 274170
rect 129154 274046 129250 274102
rect 129306 274046 129374 274102
rect 129430 274046 129498 274102
rect 129554 274046 129622 274102
rect 129678 274046 129774 274102
rect 129154 273978 129774 274046
rect 129154 273922 129250 273978
rect 129306 273922 129374 273978
rect 129430 273922 129498 273978
rect 129554 273922 129622 273978
rect 129678 273922 129774 273978
rect 129154 256350 129774 273922
rect 129154 256294 129250 256350
rect 129306 256294 129374 256350
rect 129430 256294 129498 256350
rect 129554 256294 129622 256350
rect 129678 256294 129774 256350
rect 129154 256226 129774 256294
rect 129154 256170 129250 256226
rect 129306 256170 129374 256226
rect 129430 256170 129498 256226
rect 129554 256170 129622 256226
rect 129678 256170 129774 256226
rect 129154 256102 129774 256170
rect 129154 256046 129250 256102
rect 129306 256046 129374 256102
rect 129430 256046 129498 256102
rect 129554 256046 129622 256102
rect 129678 256046 129774 256102
rect 129154 255978 129774 256046
rect 129154 255922 129250 255978
rect 129306 255922 129374 255978
rect 129430 255922 129498 255978
rect 129554 255922 129622 255978
rect 129678 255922 129774 255978
rect 129154 238350 129774 255922
rect 129154 238294 129250 238350
rect 129306 238294 129374 238350
rect 129430 238294 129498 238350
rect 129554 238294 129622 238350
rect 129678 238294 129774 238350
rect 129154 238226 129774 238294
rect 129154 238170 129250 238226
rect 129306 238170 129374 238226
rect 129430 238170 129498 238226
rect 129554 238170 129622 238226
rect 129678 238170 129774 238226
rect 129154 238102 129774 238170
rect 129154 238046 129250 238102
rect 129306 238046 129374 238102
rect 129430 238046 129498 238102
rect 129554 238046 129622 238102
rect 129678 238046 129774 238102
rect 129154 237978 129774 238046
rect 129154 237922 129250 237978
rect 129306 237922 129374 237978
rect 129430 237922 129498 237978
rect 129554 237922 129622 237978
rect 129678 237922 129774 237978
rect 129154 220350 129774 237922
rect 129154 220294 129250 220350
rect 129306 220294 129374 220350
rect 129430 220294 129498 220350
rect 129554 220294 129622 220350
rect 129678 220294 129774 220350
rect 129154 220226 129774 220294
rect 129154 220170 129250 220226
rect 129306 220170 129374 220226
rect 129430 220170 129498 220226
rect 129554 220170 129622 220226
rect 129678 220170 129774 220226
rect 129154 220102 129774 220170
rect 129154 220046 129250 220102
rect 129306 220046 129374 220102
rect 129430 220046 129498 220102
rect 129554 220046 129622 220102
rect 129678 220046 129774 220102
rect 129154 219978 129774 220046
rect 129154 219922 129250 219978
rect 129306 219922 129374 219978
rect 129430 219922 129498 219978
rect 129554 219922 129622 219978
rect 129678 219922 129774 219978
rect 129154 202350 129774 219922
rect 129154 202294 129250 202350
rect 129306 202294 129374 202350
rect 129430 202294 129498 202350
rect 129554 202294 129622 202350
rect 129678 202294 129774 202350
rect 129154 202226 129774 202294
rect 129154 202170 129250 202226
rect 129306 202170 129374 202226
rect 129430 202170 129498 202226
rect 129554 202170 129622 202226
rect 129678 202170 129774 202226
rect 129154 202102 129774 202170
rect 129154 202046 129250 202102
rect 129306 202046 129374 202102
rect 129430 202046 129498 202102
rect 129554 202046 129622 202102
rect 129678 202046 129774 202102
rect 129154 201978 129774 202046
rect 129154 201922 129250 201978
rect 129306 201922 129374 201978
rect 129430 201922 129498 201978
rect 129554 201922 129622 201978
rect 129678 201922 129774 201978
rect 129154 184350 129774 201922
rect 129154 184294 129250 184350
rect 129306 184294 129374 184350
rect 129430 184294 129498 184350
rect 129554 184294 129622 184350
rect 129678 184294 129774 184350
rect 129154 184226 129774 184294
rect 129154 184170 129250 184226
rect 129306 184170 129374 184226
rect 129430 184170 129498 184226
rect 129554 184170 129622 184226
rect 129678 184170 129774 184226
rect 129154 184102 129774 184170
rect 129154 184046 129250 184102
rect 129306 184046 129374 184102
rect 129430 184046 129498 184102
rect 129554 184046 129622 184102
rect 129678 184046 129774 184102
rect 129154 183978 129774 184046
rect 129154 183922 129250 183978
rect 129306 183922 129374 183978
rect 129430 183922 129498 183978
rect 129554 183922 129622 183978
rect 129678 183922 129774 183978
rect 129154 166350 129774 183922
rect 129154 166294 129250 166350
rect 129306 166294 129374 166350
rect 129430 166294 129498 166350
rect 129554 166294 129622 166350
rect 129678 166294 129774 166350
rect 129154 166226 129774 166294
rect 129154 166170 129250 166226
rect 129306 166170 129374 166226
rect 129430 166170 129498 166226
rect 129554 166170 129622 166226
rect 129678 166170 129774 166226
rect 129154 166102 129774 166170
rect 129154 166046 129250 166102
rect 129306 166046 129374 166102
rect 129430 166046 129498 166102
rect 129554 166046 129622 166102
rect 129678 166046 129774 166102
rect 129154 165978 129774 166046
rect 129154 165922 129250 165978
rect 129306 165922 129374 165978
rect 129430 165922 129498 165978
rect 129554 165922 129622 165978
rect 129678 165922 129774 165978
rect 129154 148350 129774 165922
rect 129154 148294 129250 148350
rect 129306 148294 129374 148350
rect 129430 148294 129498 148350
rect 129554 148294 129622 148350
rect 129678 148294 129774 148350
rect 129154 148226 129774 148294
rect 129154 148170 129250 148226
rect 129306 148170 129374 148226
rect 129430 148170 129498 148226
rect 129554 148170 129622 148226
rect 129678 148170 129774 148226
rect 129154 148102 129774 148170
rect 129154 148046 129250 148102
rect 129306 148046 129374 148102
rect 129430 148046 129498 148102
rect 129554 148046 129622 148102
rect 129678 148046 129774 148102
rect 129154 147978 129774 148046
rect 129154 147922 129250 147978
rect 129306 147922 129374 147978
rect 129430 147922 129498 147978
rect 129554 147922 129622 147978
rect 129678 147922 129774 147978
rect 129154 130350 129774 147922
rect 129154 130294 129250 130350
rect 129306 130294 129374 130350
rect 129430 130294 129498 130350
rect 129554 130294 129622 130350
rect 129678 130294 129774 130350
rect 129154 130226 129774 130294
rect 129154 130170 129250 130226
rect 129306 130170 129374 130226
rect 129430 130170 129498 130226
rect 129554 130170 129622 130226
rect 129678 130170 129774 130226
rect 129154 130102 129774 130170
rect 129154 130046 129250 130102
rect 129306 130046 129374 130102
rect 129430 130046 129498 130102
rect 129554 130046 129622 130102
rect 129678 130046 129774 130102
rect 129154 129978 129774 130046
rect 129154 129922 129250 129978
rect 129306 129922 129374 129978
rect 129430 129922 129498 129978
rect 129554 129922 129622 129978
rect 129678 129922 129774 129978
rect 129154 112350 129774 129922
rect 129154 112294 129250 112350
rect 129306 112294 129374 112350
rect 129430 112294 129498 112350
rect 129554 112294 129622 112350
rect 129678 112294 129774 112350
rect 129154 112226 129774 112294
rect 129154 112170 129250 112226
rect 129306 112170 129374 112226
rect 129430 112170 129498 112226
rect 129554 112170 129622 112226
rect 129678 112170 129774 112226
rect 129154 112102 129774 112170
rect 129154 112046 129250 112102
rect 129306 112046 129374 112102
rect 129430 112046 129498 112102
rect 129554 112046 129622 112102
rect 129678 112046 129774 112102
rect 129154 111978 129774 112046
rect 129154 111922 129250 111978
rect 129306 111922 129374 111978
rect 129430 111922 129498 111978
rect 129554 111922 129622 111978
rect 129678 111922 129774 111978
rect 129154 94350 129774 111922
rect 129154 94294 129250 94350
rect 129306 94294 129374 94350
rect 129430 94294 129498 94350
rect 129554 94294 129622 94350
rect 129678 94294 129774 94350
rect 129154 94226 129774 94294
rect 129154 94170 129250 94226
rect 129306 94170 129374 94226
rect 129430 94170 129498 94226
rect 129554 94170 129622 94226
rect 129678 94170 129774 94226
rect 129154 94102 129774 94170
rect 129154 94046 129250 94102
rect 129306 94046 129374 94102
rect 129430 94046 129498 94102
rect 129554 94046 129622 94102
rect 129678 94046 129774 94102
rect 129154 93978 129774 94046
rect 129154 93922 129250 93978
rect 129306 93922 129374 93978
rect 129430 93922 129498 93978
rect 129554 93922 129622 93978
rect 129678 93922 129774 93978
rect 129154 76350 129774 93922
rect 129154 76294 129250 76350
rect 129306 76294 129374 76350
rect 129430 76294 129498 76350
rect 129554 76294 129622 76350
rect 129678 76294 129774 76350
rect 129154 76226 129774 76294
rect 129154 76170 129250 76226
rect 129306 76170 129374 76226
rect 129430 76170 129498 76226
rect 129554 76170 129622 76226
rect 129678 76170 129774 76226
rect 129154 76102 129774 76170
rect 129154 76046 129250 76102
rect 129306 76046 129374 76102
rect 129430 76046 129498 76102
rect 129554 76046 129622 76102
rect 129678 76046 129774 76102
rect 129154 75978 129774 76046
rect 129154 75922 129250 75978
rect 129306 75922 129374 75978
rect 129430 75922 129498 75978
rect 129554 75922 129622 75978
rect 129678 75922 129774 75978
rect 129154 58350 129774 75922
rect 129154 58294 129250 58350
rect 129306 58294 129374 58350
rect 129430 58294 129498 58350
rect 129554 58294 129622 58350
rect 129678 58294 129774 58350
rect 129154 58226 129774 58294
rect 129154 58170 129250 58226
rect 129306 58170 129374 58226
rect 129430 58170 129498 58226
rect 129554 58170 129622 58226
rect 129678 58170 129774 58226
rect 129154 58102 129774 58170
rect 129154 58046 129250 58102
rect 129306 58046 129374 58102
rect 129430 58046 129498 58102
rect 129554 58046 129622 58102
rect 129678 58046 129774 58102
rect 129154 57978 129774 58046
rect 129154 57922 129250 57978
rect 129306 57922 129374 57978
rect 129430 57922 129498 57978
rect 129554 57922 129622 57978
rect 129678 57922 129774 57978
rect 129154 40350 129774 57922
rect 129154 40294 129250 40350
rect 129306 40294 129374 40350
rect 129430 40294 129498 40350
rect 129554 40294 129622 40350
rect 129678 40294 129774 40350
rect 129154 40226 129774 40294
rect 129154 40170 129250 40226
rect 129306 40170 129374 40226
rect 129430 40170 129498 40226
rect 129554 40170 129622 40226
rect 129678 40170 129774 40226
rect 129154 40102 129774 40170
rect 129154 40046 129250 40102
rect 129306 40046 129374 40102
rect 129430 40046 129498 40102
rect 129554 40046 129622 40102
rect 129678 40046 129774 40102
rect 129154 39978 129774 40046
rect 129154 39922 129250 39978
rect 129306 39922 129374 39978
rect 129430 39922 129498 39978
rect 129554 39922 129622 39978
rect 129678 39922 129774 39978
rect 129154 22350 129774 39922
rect 129154 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 129774 22350
rect 129154 22226 129774 22294
rect 129154 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 129774 22226
rect 129154 22102 129774 22170
rect 129154 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 129774 22102
rect 129154 21978 129774 22046
rect 129154 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 129774 21978
rect 129154 4350 129774 21922
rect 129154 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 129774 4350
rect 129154 4226 129774 4294
rect 129154 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 129774 4226
rect 129154 4102 129774 4170
rect 129154 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 129774 4102
rect 129154 3978 129774 4046
rect 129154 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 129774 3978
rect 129154 -160 129774 3922
rect 129154 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 129774 -160
rect 129154 -284 129774 -216
rect 129154 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 129774 -284
rect 129154 -408 129774 -340
rect 129154 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 129774 -408
rect 129154 -532 129774 -464
rect 129154 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 129774 -532
rect 129154 -1644 129774 -588
rect 132874 598172 133494 598268
rect 132874 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 133494 598172
rect 132874 598048 133494 598116
rect 132874 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 133494 598048
rect 132874 597924 133494 597992
rect 132874 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 133494 597924
rect 132874 597800 133494 597868
rect 132874 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 133494 597800
rect 132874 586350 133494 597744
rect 132874 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 133494 586350
rect 132874 586226 133494 586294
rect 132874 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 133494 586226
rect 132874 586102 133494 586170
rect 132874 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 133494 586102
rect 132874 585978 133494 586046
rect 132874 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 133494 585978
rect 132874 568350 133494 585922
rect 132874 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 133494 568350
rect 132874 568226 133494 568294
rect 132874 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 133494 568226
rect 132874 568102 133494 568170
rect 132874 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 133494 568102
rect 132874 567978 133494 568046
rect 132874 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 133494 567978
rect 132874 550350 133494 567922
rect 132874 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 133494 550350
rect 132874 550226 133494 550294
rect 132874 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 133494 550226
rect 132874 550102 133494 550170
rect 132874 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 133494 550102
rect 132874 549978 133494 550046
rect 132874 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 133494 549978
rect 132874 532350 133494 549922
rect 132874 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 133494 532350
rect 132874 532226 133494 532294
rect 132874 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 133494 532226
rect 132874 532102 133494 532170
rect 132874 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 133494 532102
rect 132874 531978 133494 532046
rect 132874 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 133494 531978
rect 132874 514350 133494 531922
rect 132874 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 133494 514350
rect 132874 514226 133494 514294
rect 132874 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 133494 514226
rect 132874 514102 133494 514170
rect 132874 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 133494 514102
rect 132874 513978 133494 514046
rect 132874 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 133494 513978
rect 132874 496350 133494 513922
rect 132874 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 133494 496350
rect 132874 496226 133494 496294
rect 132874 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 133494 496226
rect 132874 496102 133494 496170
rect 132874 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 133494 496102
rect 132874 495978 133494 496046
rect 132874 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 133494 495978
rect 132874 478350 133494 495922
rect 132874 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 133494 478350
rect 132874 478226 133494 478294
rect 132874 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 133494 478226
rect 132874 478102 133494 478170
rect 132874 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 133494 478102
rect 132874 477978 133494 478046
rect 132874 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 133494 477978
rect 132874 460350 133494 477922
rect 132874 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 133494 460350
rect 132874 460226 133494 460294
rect 132874 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 133494 460226
rect 132874 460102 133494 460170
rect 132874 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 133494 460102
rect 132874 459978 133494 460046
rect 132874 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 133494 459978
rect 132874 442350 133494 459922
rect 132874 442294 132970 442350
rect 133026 442294 133094 442350
rect 133150 442294 133218 442350
rect 133274 442294 133342 442350
rect 133398 442294 133494 442350
rect 132874 442226 133494 442294
rect 132874 442170 132970 442226
rect 133026 442170 133094 442226
rect 133150 442170 133218 442226
rect 133274 442170 133342 442226
rect 133398 442170 133494 442226
rect 132874 442102 133494 442170
rect 132874 442046 132970 442102
rect 133026 442046 133094 442102
rect 133150 442046 133218 442102
rect 133274 442046 133342 442102
rect 133398 442046 133494 442102
rect 132874 441978 133494 442046
rect 132874 441922 132970 441978
rect 133026 441922 133094 441978
rect 133150 441922 133218 441978
rect 133274 441922 133342 441978
rect 133398 441922 133494 441978
rect 132874 424350 133494 441922
rect 132874 424294 132970 424350
rect 133026 424294 133094 424350
rect 133150 424294 133218 424350
rect 133274 424294 133342 424350
rect 133398 424294 133494 424350
rect 132874 424226 133494 424294
rect 132874 424170 132970 424226
rect 133026 424170 133094 424226
rect 133150 424170 133218 424226
rect 133274 424170 133342 424226
rect 133398 424170 133494 424226
rect 132874 424102 133494 424170
rect 132874 424046 132970 424102
rect 133026 424046 133094 424102
rect 133150 424046 133218 424102
rect 133274 424046 133342 424102
rect 133398 424046 133494 424102
rect 132874 423978 133494 424046
rect 132874 423922 132970 423978
rect 133026 423922 133094 423978
rect 133150 423922 133218 423978
rect 133274 423922 133342 423978
rect 133398 423922 133494 423978
rect 132874 406350 133494 423922
rect 132874 406294 132970 406350
rect 133026 406294 133094 406350
rect 133150 406294 133218 406350
rect 133274 406294 133342 406350
rect 133398 406294 133494 406350
rect 132874 406226 133494 406294
rect 132874 406170 132970 406226
rect 133026 406170 133094 406226
rect 133150 406170 133218 406226
rect 133274 406170 133342 406226
rect 133398 406170 133494 406226
rect 132874 406102 133494 406170
rect 132874 406046 132970 406102
rect 133026 406046 133094 406102
rect 133150 406046 133218 406102
rect 133274 406046 133342 406102
rect 133398 406046 133494 406102
rect 132874 405978 133494 406046
rect 132874 405922 132970 405978
rect 133026 405922 133094 405978
rect 133150 405922 133218 405978
rect 133274 405922 133342 405978
rect 133398 405922 133494 405978
rect 132874 388350 133494 405922
rect 132874 388294 132970 388350
rect 133026 388294 133094 388350
rect 133150 388294 133218 388350
rect 133274 388294 133342 388350
rect 133398 388294 133494 388350
rect 132874 388226 133494 388294
rect 132874 388170 132970 388226
rect 133026 388170 133094 388226
rect 133150 388170 133218 388226
rect 133274 388170 133342 388226
rect 133398 388170 133494 388226
rect 132874 388102 133494 388170
rect 132874 388046 132970 388102
rect 133026 388046 133094 388102
rect 133150 388046 133218 388102
rect 133274 388046 133342 388102
rect 133398 388046 133494 388102
rect 132874 387978 133494 388046
rect 132874 387922 132970 387978
rect 133026 387922 133094 387978
rect 133150 387922 133218 387978
rect 133274 387922 133342 387978
rect 133398 387922 133494 387978
rect 132874 370350 133494 387922
rect 132874 370294 132970 370350
rect 133026 370294 133094 370350
rect 133150 370294 133218 370350
rect 133274 370294 133342 370350
rect 133398 370294 133494 370350
rect 132874 370226 133494 370294
rect 132874 370170 132970 370226
rect 133026 370170 133094 370226
rect 133150 370170 133218 370226
rect 133274 370170 133342 370226
rect 133398 370170 133494 370226
rect 132874 370102 133494 370170
rect 132874 370046 132970 370102
rect 133026 370046 133094 370102
rect 133150 370046 133218 370102
rect 133274 370046 133342 370102
rect 133398 370046 133494 370102
rect 132874 369978 133494 370046
rect 132874 369922 132970 369978
rect 133026 369922 133094 369978
rect 133150 369922 133218 369978
rect 133274 369922 133342 369978
rect 133398 369922 133494 369978
rect 132874 352350 133494 369922
rect 132874 352294 132970 352350
rect 133026 352294 133094 352350
rect 133150 352294 133218 352350
rect 133274 352294 133342 352350
rect 133398 352294 133494 352350
rect 132874 352226 133494 352294
rect 132874 352170 132970 352226
rect 133026 352170 133094 352226
rect 133150 352170 133218 352226
rect 133274 352170 133342 352226
rect 133398 352170 133494 352226
rect 132874 352102 133494 352170
rect 132874 352046 132970 352102
rect 133026 352046 133094 352102
rect 133150 352046 133218 352102
rect 133274 352046 133342 352102
rect 133398 352046 133494 352102
rect 132874 351978 133494 352046
rect 132874 351922 132970 351978
rect 133026 351922 133094 351978
rect 133150 351922 133218 351978
rect 133274 351922 133342 351978
rect 133398 351922 133494 351978
rect 132874 334350 133494 351922
rect 132874 334294 132970 334350
rect 133026 334294 133094 334350
rect 133150 334294 133218 334350
rect 133274 334294 133342 334350
rect 133398 334294 133494 334350
rect 132874 334226 133494 334294
rect 132874 334170 132970 334226
rect 133026 334170 133094 334226
rect 133150 334170 133218 334226
rect 133274 334170 133342 334226
rect 133398 334170 133494 334226
rect 132874 334102 133494 334170
rect 132874 334046 132970 334102
rect 133026 334046 133094 334102
rect 133150 334046 133218 334102
rect 133274 334046 133342 334102
rect 133398 334046 133494 334102
rect 132874 333978 133494 334046
rect 132874 333922 132970 333978
rect 133026 333922 133094 333978
rect 133150 333922 133218 333978
rect 133274 333922 133342 333978
rect 133398 333922 133494 333978
rect 132874 316350 133494 333922
rect 132874 316294 132970 316350
rect 133026 316294 133094 316350
rect 133150 316294 133218 316350
rect 133274 316294 133342 316350
rect 133398 316294 133494 316350
rect 132874 316226 133494 316294
rect 132874 316170 132970 316226
rect 133026 316170 133094 316226
rect 133150 316170 133218 316226
rect 133274 316170 133342 316226
rect 133398 316170 133494 316226
rect 132874 316102 133494 316170
rect 132874 316046 132970 316102
rect 133026 316046 133094 316102
rect 133150 316046 133218 316102
rect 133274 316046 133342 316102
rect 133398 316046 133494 316102
rect 132874 315978 133494 316046
rect 132874 315922 132970 315978
rect 133026 315922 133094 315978
rect 133150 315922 133218 315978
rect 133274 315922 133342 315978
rect 133398 315922 133494 315978
rect 132874 298350 133494 315922
rect 132874 298294 132970 298350
rect 133026 298294 133094 298350
rect 133150 298294 133218 298350
rect 133274 298294 133342 298350
rect 133398 298294 133494 298350
rect 132874 298226 133494 298294
rect 132874 298170 132970 298226
rect 133026 298170 133094 298226
rect 133150 298170 133218 298226
rect 133274 298170 133342 298226
rect 133398 298170 133494 298226
rect 132874 298102 133494 298170
rect 132874 298046 132970 298102
rect 133026 298046 133094 298102
rect 133150 298046 133218 298102
rect 133274 298046 133342 298102
rect 133398 298046 133494 298102
rect 132874 297978 133494 298046
rect 132874 297922 132970 297978
rect 133026 297922 133094 297978
rect 133150 297922 133218 297978
rect 133274 297922 133342 297978
rect 133398 297922 133494 297978
rect 132874 280350 133494 297922
rect 132874 280294 132970 280350
rect 133026 280294 133094 280350
rect 133150 280294 133218 280350
rect 133274 280294 133342 280350
rect 133398 280294 133494 280350
rect 132874 280226 133494 280294
rect 132874 280170 132970 280226
rect 133026 280170 133094 280226
rect 133150 280170 133218 280226
rect 133274 280170 133342 280226
rect 133398 280170 133494 280226
rect 132874 280102 133494 280170
rect 132874 280046 132970 280102
rect 133026 280046 133094 280102
rect 133150 280046 133218 280102
rect 133274 280046 133342 280102
rect 133398 280046 133494 280102
rect 132874 279978 133494 280046
rect 132874 279922 132970 279978
rect 133026 279922 133094 279978
rect 133150 279922 133218 279978
rect 133274 279922 133342 279978
rect 133398 279922 133494 279978
rect 132874 262350 133494 279922
rect 132874 262294 132970 262350
rect 133026 262294 133094 262350
rect 133150 262294 133218 262350
rect 133274 262294 133342 262350
rect 133398 262294 133494 262350
rect 132874 262226 133494 262294
rect 132874 262170 132970 262226
rect 133026 262170 133094 262226
rect 133150 262170 133218 262226
rect 133274 262170 133342 262226
rect 133398 262170 133494 262226
rect 132874 262102 133494 262170
rect 132874 262046 132970 262102
rect 133026 262046 133094 262102
rect 133150 262046 133218 262102
rect 133274 262046 133342 262102
rect 133398 262046 133494 262102
rect 132874 261978 133494 262046
rect 132874 261922 132970 261978
rect 133026 261922 133094 261978
rect 133150 261922 133218 261978
rect 133274 261922 133342 261978
rect 133398 261922 133494 261978
rect 132874 244350 133494 261922
rect 132874 244294 132970 244350
rect 133026 244294 133094 244350
rect 133150 244294 133218 244350
rect 133274 244294 133342 244350
rect 133398 244294 133494 244350
rect 132874 244226 133494 244294
rect 132874 244170 132970 244226
rect 133026 244170 133094 244226
rect 133150 244170 133218 244226
rect 133274 244170 133342 244226
rect 133398 244170 133494 244226
rect 132874 244102 133494 244170
rect 132874 244046 132970 244102
rect 133026 244046 133094 244102
rect 133150 244046 133218 244102
rect 133274 244046 133342 244102
rect 133398 244046 133494 244102
rect 132874 243978 133494 244046
rect 132874 243922 132970 243978
rect 133026 243922 133094 243978
rect 133150 243922 133218 243978
rect 133274 243922 133342 243978
rect 133398 243922 133494 243978
rect 132874 226350 133494 243922
rect 132874 226294 132970 226350
rect 133026 226294 133094 226350
rect 133150 226294 133218 226350
rect 133274 226294 133342 226350
rect 133398 226294 133494 226350
rect 132874 226226 133494 226294
rect 132874 226170 132970 226226
rect 133026 226170 133094 226226
rect 133150 226170 133218 226226
rect 133274 226170 133342 226226
rect 133398 226170 133494 226226
rect 132874 226102 133494 226170
rect 132874 226046 132970 226102
rect 133026 226046 133094 226102
rect 133150 226046 133218 226102
rect 133274 226046 133342 226102
rect 133398 226046 133494 226102
rect 132874 225978 133494 226046
rect 132874 225922 132970 225978
rect 133026 225922 133094 225978
rect 133150 225922 133218 225978
rect 133274 225922 133342 225978
rect 133398 225922 133494 225978
rect 132874 208350 133494 225922
rect 132874 208294 132970 208350
rect 133026 208294 133094 208350
rect 133150 208294 133218 208350
rect 133274 208294 133342 208350
rect 133398 208294 133494 208350
rect 132874 208226 133494 208294
rect 132874 208170 132970 208226
rect 133026 208170 133094 208226
rect 133150 208170 133218 208226
rect 133274 208170 133342 208226
rect 133398 208170 133494 208226
rect 132874 208102 133494 208170
rect 132874 208046 132970 208102
rect 133026 208046 133094 208102
rect 133150 208046 133218 208102
rect 133274 208046 133342 208102
rect 133398 208046 133494 208102
rect 132874 207978 133494 208046
rect 132874 207922 132970 207978
rect 133026 207922 133094 207978
rect 133150 207922 133218 207978
rect 133274 207922 133342 207978
rect 133398 207922 133494 207978
rect 132874 190350 133494 207922
rect 132874 190294 132970 190350
rect 133026 190294 133094 190350
rect 133150 190294 133218 190350
rect 133274 190294 133342 190350
rect 133398 190294 133494 190350
rect 132874 190226 133494 190294
rect 132874 190170 132970 190226
rect 133026 190170 133094 190226
rect 133150 190170 133218 190226
rect 133274 190170 133342 190226
rect 133398 190170 133494 190226
rect 132874 190102 133494 190170
rect 132874 190046 132970 190102
rect 133026 190046 133094 190102
rect 133150 190046 133218 190102
rect 133274 190046 133342 190102
rect 133398 190046 133494 190102
rect 132874 189978 133494 190046
rect 132874 189922 132970 189978
rect 133026 189922 133094 189978
rect 133150 189922 133218 189978
rect 133274 189922 133342 189978
rect 133398 189922 133494 189978
rect 132874 172350 133494 189922
rect 132874 172294 132970 172350
rect 133026 172294 133094 172350
rect 133150 172294 133218 172350
rect 133274 172294 133342 172350
rect 133398 172294 133494 172350
rect 132874 172226 133494 172294
rect 132874 172170 132970 172226
rect 133026 172170 133094 172226
rect 133150 172170 133218 172226
rect 133274 172170 133342 172226
rect 133398 172170 133494 172226
rect 132874 172102 133494 172170
rect 132874 172046 132970 172102
rect 133026 172046 133094 172102
rect 133150 172046 133218 172102
rect 133274 172046 133342 172102
rect 133398 172046 133494 172102
rect 132874 171978 133494 172046
rect 132874 171922 132970 171978
rect 133026 171922 133094 171978
rect 133150 171922 133218 171978
rect 133274 171922 133342 171978
rect 133398 171922 133494 171978
rect 132874 154350 133494 171922
rect 132874 154294 132970 154350
rect 133026 154294 133094 154350
rect 133150 154294 133218 154350
rect 133274 154294 133342 154350
rect 133398 154294 133494 154350
rect 132874 154226 133494 154294
rect 132874 154170 132970 154226
rect 133026 154170 133094 154226
rect 133150 154170 133218 154226
rect 133274 154170 133342 154226
rect 133398 154170 133494 154226
rect 132874 154102 133494 154170
rect 132874 154046 132970 154102
rect 133026 154046 133094 154102
rect 133150 154046 133218 154102
rect 133274 154046 133342 154102
rect 133398 154046 133494 154102
rect 132874 153978 133494 154046
rect 132874 153922 132970 153978
rect 133026 153922 133094 153978
rect 133150 153922 133218 153978
rect 133274 153922 133342 153978
rect 133398 153922 133494 153978
rect 132874 136350 133494 153922
rect 132874 136294 132970 136350
rect 133026 136294 133094 136350
rect 133150 136294 133218 136350
rect 133274 136294 133342 136350
rect 133398 136294 133494 136350
rect 132874 136226 133494 136294
rect 132874 136170 132970 136226
rect 133026 136170 133094 136226
rect 133150 136170 133218 136226
rect 133274 136170 133342 136226
rect 133398 136170 133494 136226
rect 132874 136102 133494 136170
rect 132874 136046 132970 136102
rect 133026 136046 133094 136102
rect 133150 136046 133218 136102
rect 133274 136046 133342 136102
rect 133398 136046 133494 136102
rect 132874 135978 133494 136046
rect 132874 135922 132970 135978
rect 133026 135922 133094 135978
rect 133150 135922 133218 135978
rect 133274 135922 133342 135978
rect 133398 135922 133494 135978
rect 132874 118350 133494 135922
rect 132874 118294 132970 118350
rect 133026 118294 133094 118350
rect 133150 118294 133218 118350
rect 133274 118294 133342 118350
rect 133398 118294 133494 118350
rect 132874 118226 133494 118294
rect 132874 118170 132970 118226
rect 133026 118170 133094 118226
rect 133150 118170 133218 118226
rect 133274 118170 133342 118226
rect 133398 118170 133494 118226
rect 132874 118102 133494 118170
rect 132874 118046 132970 118102
rect 133026 118046 133094 118102
rect 133150 118046 133218 118102
rect 133274 118046 133342 118102
rect 133398 118046 133494 118102
rect 132874 117978 133494 118046
rect 132874 117922 132970 117978
rect 133026 117922 133094 117978
rect 133150 117922 133218 117978
rect 133274 117922 133342 117978
rect 133398 117922 133494 117978
rect 132874 100350 133494 117922
rect 132874 100294 132970 100350
rect 133026 100294 133094 100350
rect 133150 100294 133218 100350
rect 133274 100294 133342 100350
rect 133398 100294 133494 100350
rect 132874 100226 133494 100294
rect 132874 100170 132970 100226
rect 133026 100170 133094 100226
rect 133150 100170 133218 100226
rect 133274 100170 133342 100226
rect 133398 100170 133494 100226
rect 132874 100102 133494 100170
rect 132874 100046 132970 100102
rect 133026 100046 133094 100102
rect 133150 100046 133218 100102
rect 133274 100046 133342 100102
rect 133398 100046 133494 100102
rect 132874 99978 133494 100046
rect 132874 99922 132970 99978
rect 133026 99922 133094 99978
rect 133150 99922 133218 99978
rect 133274 99922 133342 99978
rect 133398 99922 133494 99978
rect 132874 82350 133494 99922
rect 132874 82294 132970 82350
rect 133026 82294 133094 82350
rect 133150 82294 133218 82350
rect 133274 82294 133342 82350
rect 133398 82294 133494 82350
rect 132874 82226 133494 82294
rect 132874 82170 132970 82226
rect 133026 82170 133094 82226
rect 133150 82170 133218 82226
rect 133274 82170 133342 82226
rect 133398 82170 133494 82226
rect 132874 82102 133494 82170
rect 132874 82046 132970 82102
rect 133026 82046 133094 82102
rect 133150 82046 133218 82102
rect 133274 82046 133342 82102
rect 133398 82046 133494 82102
rect 132874 81978 133494 82046
rect 132874 81922 132970 81978
rect 133026 81922 133094 81978
rect 133150 81922 133218 81978
rect 133274 81922 133342 81978
rect 133398 81922 133494 81978
rect 132874 64350 133494 81922
rect 132874 64294 132970 64350
rect 133026 64294 133094 64350
rect 133150 64294 133218 64350
rect 133274 64294 133342 64350
rect 133398 64294 133494 64350
rect 132874 64226 133494 64294
rect 132874 64170 132970 64226
rect 133026 64170 133094 64226
rect 133150 64170 133218 64226
rect 133274 64170 133342 64226
rect 133398 64170 133494 64226
rect 132874 64102 133494 64170
rect 132874 64046 132970 64102
rect 133026 64046 133094 64102
rect 133150 64046 133218 64102
rect 133274 64046 133342 64102
rect 133398 64046 133494 64102
rect 132874 63978 133494 64046
rect 132874 63922 132970 63978
rect 133026 63922 133094 63978
rect 133150 63922 133218 63978
rect 133274 63922 133342 63978
rect 133398 63922 133494 63978
rect 132874 46350 133494 63922
rect 132874 46294 132970 46350
rect 133026 46294 133094 46350
rect 133150 46294 133218 46350
rect 133274 46294 133342 46350
rect 133398 46294 133494 46350
rect 132874 46226 133494 46294
rect 132874 46170 132970 46226
rect 133026 46170 133094 46226
rect 133150 46170 133218 46226
rect 133274 46170 133342 46226
rect 133398 46170 133494 46226
rect 132874 46102 133494 46170
rect 132874 46046 132970 46102
rect 133026 46046 133094 46102
rect 133150 46046 133218 46102
rect 133274 46046 133342 46102
rect 133398 46046 133494 46102
rect 132874 45978 133494 46046
rect 132874 45922 132970 45978
rect 133026 45922 133094 45978
rect 133150 45922 133218 45978
rect 133274 45922 133342 45978
rect 133398 45922 133494 45978
rect 132874 28350 133494 45922
rect 132874 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 133494 28350
rect 132874 28226 133494 28294
rect 132874 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 133494 28226
rect 132874 28102 133494 28170
rect 132874 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 133494 28102
rect 132874 27978 133494 28046
rect 132874 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 133494 27978
rect 132874 10350 133494 27922
rect 132874 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 133494 10350
rect 132874 10226 133494 10294
rect 132874 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 133494 10226
rect 132874 10102 133494 10170
rect 132874 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 133494 10102
rect 132874 9978 133494 10046
rect 132874 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 133494 9978
rect 132874 -1120 133494 9922
rect 132874 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 133494 -1120
rect 132874 -1244 133494 -1176
rect 132874 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 133494 -1244
rect 132874 -1368 133494 -1300
rect 132874 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 133494 -1368
rect 132874 -1492 133494 -1424
rect 132874 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 133494 -1492
rect 132874 -1644 133494 -1548
rect 147154 597212 147774 598268
rect 147154 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 147774 597212
rect 147154 597088 147774 597156
rect 147154 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 147774 597088
rect 147154 596964 147774 597032
rect 147154 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 147774 596964
rect 147154 596840 147774 596908
rect 147154 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 147774 596840
rect 147154 580350 147774 596784
rect 147154 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 147774 580350
rect 147154 580226 147774 580294
rect 147154 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 147774 580226
rect 147154 580102 147774 580170
rect 147154 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 147774 580102
rect 147154 579978 147774 580046
rect 147154 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 147774 579978
rect 147154 562350 147774 579922
rect 147154 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 147774 562350
rect 147154 562226 147774 562294
rect 147154 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 147774 562226
rect 147154 562102 147774 562170
rect 147154 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 147774 562102
rect 147154 561978 147774 562046
rect 147154 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 147774 561978
rect 147154 544350 147774 561922
rect 147154 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 147774 544350
rect 147154 544226 147774 544294
rect 147154 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 147774 544226
rect 147154 544102 147774 544170
rect 147154 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 147774 544102
rect 147154 543978 147774 544046
rect 147154 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 147774 543978
rect 147154 526350 147774 543922
rect 147154 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 147774 526350
rect 147154 526226 147774 526294
rect 147154 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 147774 526226
rect 147154 526102 147774 526170
rect 147154 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 147774 526102
rect 147154 525978 147774 526046
rect 147154 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 147774 525978
rect 147154 508350 147774 525922
rect 147154 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 147774 508350
rect 147154 508226 147774 508294
rect 147154 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 147774 508226
rect 147154 508102 147774 508170
rect 147154 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 147774 508102
rect 147154 507978 147774 508046
rect 147154 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 147774 507978
rect 147154 490350 147774 507922
rect 147154 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 147774 490350
rect 147154 490226 147774 490294
rect 147154 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 147774 490226
rect 147154 490102 147774 490170
rect 147154 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 147774 490102
rect 147154 489978 147774 490046
rect 147154 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 147774 489978
rect 147154 472350 147774 489922
rect 147154 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 147774 472350
rect 147154 472226 147774 472294
rect 147154 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 147774 472226
rect 147154 472102 147774 472170
rect 147154 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 147774 472102
rect 147154 471978 147774 472046
rect 147154 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 147774 471978
rect 147154 454350 147774 471922
rect 147154 454294 147250 454350
rect 147306 454294 147374 454350
rect 147430 454294 147498 454350
rect 147554 454294 147622 454350
rect 147678 454294 147774 454350
rect 147154 454226 147774 454294
rect 147154 454170 147250 454226
rect 147306 454170 147374 454226
rect 147430 454170 147498 454226
rect 147554 454170 147622 454226
rect 147678 454170 147774 454226
rect 147154 454102 147774 454170
rect 147154 454046 147250 454102
rect 147306 454046 147374 454102
rect 147430 454046 147498 454102
rect 147554 454046 147622 454102
rect 147678 454046 147774 454102
rect 147154 453978 147774 454046
rect 147154 453922 147250 453978
rect 147306 453922 147374 453978
rect 147430 453922 147498 453978
rect 147554 453922 147622 453978
rect 147678 453922 147774 453978
rect 147154 436350 147774 453922
rect 147154 436294 147250 436350
rect 147306 436294 147374 436350
rect 147430 436294 147498 436350
rect 147554 436294 147622 436350
rect 147678 436294 147774 436350
rect 147154 436226 147774 436294
rect 147154 436170 147250 436226
rect 147306 436170 147374 436226
rect 147430 436170 147498 436226
rect 147554 436170 147622 436226
rect 147678 436170 147774 436226
rect 147154 436102 147774 436170
rect 147154 436046 147250 436102
rect 147306 436046 147374 436102
rect 147430 436046 147498 436102
rect 147554 436046 147622 436102
rect 147678 436046 147774 436102
rect 147154 435978 147774 436046
rect 147154 435922 147250 435978
rect 147306 435922 147374 435978
rect 147430 435922 147498 435978
rect 147554 435922 147622 435978
rect 147678 435922 147774 435978
rect 147154 418350 147774 435922
rect 147154 418294 147250 418350
rect 147306 418294 147374 418350
rect 147430 418294 147498 418350
rect 147554 418294 147622 418350
rect 147678 418294 147774 418350
rect 147154 418226 147774 418294
rect 147154 418170 147250 418226
rect 147306 418170 147374 418226
rect 147430 418170 147498 418226
rect 147554 418170 147622 418226
rect 147678 418170 147774 418226
rect 147154 418102 147774 418170
rect 147154 418046 147250 418102
rect 147306 418046 147374 418102
rect 147430 418046 147498 418102
rect 147554 418046 147622 418102
rect 147678 418046 147774 418102
rect 147154 417978 147774 418046
rect 147154 417922 147250 417978
rect 147306 417922 147374 417978
rect 147430 417922 147498 417978
rect 147554 417922 147622 417978
rect 147678 417922 147774 417978
rect 147154 400350 147774 417922
rect 147154 400294 147250 400350
rect 147306 400294 147374 400350
rect 147430 400294 147498 400350
rect 147554 400294 147622 400350
rect 147678 400294 147774 400350
rect 147154 400226 147774 400294
rect 147154 400170 147250 400226
rect 147306 400170 147374 400226
rect 147430 400170 147498 400226
rect 147554 400170 147622 400226
rect 147678 400170 147774 400226
rect 147154 400102 147774 400170
rect 147154 400046 147250 400102
rect 147306 400046 147374 400102
rect 147430 400046 147498 400102
rect 147554 400046 147622 400102
rect 147678 400046 147774 400102
rect 147154 399978 147774 400046
rect 147154 399922 147250 399978
rect 147306 399922 147374 399978
rect 147430 399922 147498 399978
rect 147554 399922 147622 399978
rect 147678 399922 147774 399978
rect 147154 382350 147774 399922
rect 147154 382294 147250 382350
rect 147306 382294 147374 382350
rect 147430 382294 147498 382350
rect 147554 382294 147622 382350
rect 147678 382294 147774 382350
rect 147154 382226 147774 382294
rect 147154 382170 147250 382226
rect 147306 382170 147374 382226
rect 147430 382170 147498 382226
rect 147554 382170 147622 382226
rect 147678 382170 147774 382226
rect 147154 382102 147774 382170
rect 147154 382046 147250 382102
rect 147306 382046 147374 382102
rect 147430 382046 147498 382102
rect 147554 382046 147622 382102
rect 147678 382046 147774 382102
rect 147154 381978 147774 382046
rect 147154 381922 147250 381978
rect 147306 381922 147374 381978
rect 147430 381922 147498 381978
rect 147554 381922 147622 381978
rect 147678 381922 147774 381978
rect 147154 364350 147774 381922
rect 147154 364294 147250 364350
rect 147306 364294 147374 364350
rect 147430 364294 147498 364350
rect 147554 364294 147622 364350
rect 147678 364294 147774 364350
rect 147154 364226 147774 364294
rect 147154 364170 147250 364226
rect 147306 364170 147374 364226
rect 147430 364170 147498 364226
rect 147554 364170 147622 364226
rect 147678 364170 147774 364226
rect 147154 364102 147774 364170
rect 147154 364046 147250 364102
rect 147306 364046 147374 364102
rect 147430 364046 147498 364102
rect 147554 364046 147622 364102
rect 147678 364046 147774 364102
rect 147154 363978 147774 364046
rect 147154 363922 147250 363978
rect 147306 363922 147374 363978
rect 147430 363922 147498 363978
rect 147554 363922 147622 363978
rect 147678 363922 147774 363978
rect 147154 346350 147774 363922
rect 147154 346294 147250 346350
rect 147306 346294 147374 346350
rect 147430 346294 147498 346350
rect 147554 346294 147622 346350
rect 147678 346294 147774 346350
rect 147154 346226 147774 346294
rect 147154 346170 147250 346226
rect 147306 346170 147374 346226
rect 147430 346170 147498 346226
rect 147554 346170 147622 346226
rect 147678 346170 147774 346226
rect 147154 346102 147774 346170
rect 147154 346046 147250 346102
rect 147306 346046 147374 346102
rect 147430 346046 147498 346102
rect 147554 346046 147622 346102
rect 147678 346046 147774 346102
rect 147154 345978 147774 346046
rect 147154 345922 147250 345978
rect 147306 345922 147374 345978
rect 147430 345922 147498 345978
rect 147554 345922 147622 345978
rect 147678 345922 147774 345978
rect 147154 328350 147774 345922
rect 147154 328294 147250 328350
rect 147306 328294 147374 328350
rect 147430 328294 147498 328350
rect 147554 328294 147622 328350
rect 147678 328294 147774 328350
rect 147154 328226 147774 328294
rect 147154 328170 147250 328226
rect 147306 328170 147374 328226
rect 147430 328170 147498 328226
rect 147554 328170 147622 328226
rect 147678 328170 147774 328226
rect 147154 328102 147774 328170
rect 147154 328046 147250 328102
rect 147306 328046 147374 328102
rect 147430 328046 147498 328102
rect 147554 328046 147622 328102
rect 147678 328046 147774 328102
rect 147154 327978 147774 328046
rect 147154 327922 147250 327978
rect 147306 327922 147374 327978
rect 147430 327922 147498 327978
rect 147554 327922 147622 327978
rect 147678 327922 147774 327978
rect 147154 310350 147774 327922
rect 147154 310294 147250 310350
rect 147306 310294 147374 310350
rect 147430 310294 147498 310350
rect 147554 310294 147622 310350
rect 147678 310294 147774 310350
rect 147154 310226 147774 310294
rect 147154 310170 147250 310226
rect 147306 310170 147374 310226
rect 147430 310170 147498 310226
rect 147554 310170 147622 310226
rect 147678 310170 147774 310226
rect 147154 310102 147774 310170
rect 147154 310046 147250 310102
rect 147306 310046 147374 310102
rect 147430 310046 147498 310102
rect 147554 310046 147622 310102
rect 147678 310046 147774 310102
rect 147154 309978 147774 310046
rect 147154 309922 147250 309978
rect 147306 309922 147374 309978
rect 147430 309922 147498 309978
rect 147554 309922 147622 309978
rect 147678 309922 147774 309978
rect 147154 292350 147774 309922
rect 147154 292294 147250 292350
rect 147306 292294 147374 292350
rect 147430 292294 147498 292350
rect 147554 292294 147622 292350
rect 147678 292294 147774 292350
rect 147154 292226 147774 292294
rect 147154 292170 147250 292226
rect 147306 292170 147374 292226
rect 147430 292170 147498 292226
rect 147554 292170 147622 292226
rect 147678 292170 147774 292226
rect 147154 292102 147774 292170
rect 147154 292046 147250 292102
rect 147306 292046 147374 292102
rect 147430 292046 147498 292102
rect 147554 292046 147622 292102
rect 147678 292046 147774 292102
rect 147154 291978 147774 292046
rect 147154 291922 147250 291978
rect 147306 291922 147374 291978
rect 147430 291922 147498 291978
rect 147554 291922 147622 291978
rect 147678 291922 147774 291978
rect 147154 274350 147774 291922
rect 147154 274294 147250 274350
rect 147306 274294 147374 274350
rect 147430 274294 147498 274350
rect 147554 274294 147622 274350
rect 147678 274294 147774 274350
rect 147154 274226 147774 274294
rect 147154 274170 147250 274226
rect 147306 274170 147374 274226
rect 147430 274170 147498 274226
rect 147554 274170 147622 274226
rect 147678 274170 147774 274226
rect 147154 274102 147774 274170
rect 147154 274046 147250 274102
rect 147306 274046 147374 274102
rect 147430 274046 147498 274102
rect 147554 274046 147622 274102
rect 147678 274046 147774 274102
rect 147154 273978 147774 274046
rect 147154 273922 147250 273978
rect 147306 273922 147374 273978
rect 147430 273922 147498 273978
rect 147554 273922 147622 273978
rect 147678 273922 147774 273978
rect 147154 256350 147774 273922
rect 147154 256294 147250 256350
rect 147306 256294 147374 256350
rect 147430 256294 147498 256350
rect 147554 256294 147622 256350
rect 147678 256294 147774 256350
rect 147154 256226 147774 256294
rect 147154 256170 147250 256226
rect 147306 256170 147374 256226
rect 147430 256170 147498 256226
rect 147554 256170 147622 256226
rect 147678 256170 147774 256226
rect 147154 256102 147774 256170
rect 147154 256046 147250 256102
rect 147306 256046 147374 256102
rect 147430 256046 147498 256102
rect 147554 256046 147622 256102
rect 147678 256046 147774 256102
rect 147154 255978 147774 256046
rect 147154 255922 147250 255978
rect 147306 255922 147374 255978
rect 147430 255922 147498 255978
rect 147554 255922 147622 255978
rect 147678 255922 147774 255978
rect 147154 238350 147774 255922
rect 147154 238294 147250 238350
rect 147306 238294 147374 238350
rect 147430 238294 147498 238350
rect 147554 238294 147622 238350
rect 147678 238294 147774 238350
rect 147154 238226 147774 238294
rect 147154 238170 147250 238226
rect 147306 238170 147374 238226
rect 147430 238170 147498 238226
rect 147554 238170 147622 238226
rect 147678 238170 147774 238226
rect 147154 238102 147774 238170
rect 147154 238046 147250 238102
rect 147306 238046 147374 238102
rect 147430 238046 147498 238102
rect 147554 238046 147622 238102
rect 147678 238046 147774 238102
rect 147154 237978 147774 238046
rect 147154 237922 147250 237978
rect 147306 237922 147374 237978
rect 147430 237922 147498 237978
rect 147554 237922 147622 237978
rect 147678 237922 147774 237978
rect 147154 220350 147774 237922
rect 147154 220294 147250 220350
rect 147306 220294 147374 220350
rect 147430 220294 147498 220350
rect 147554 220294 147622 220350
rect 147678 220294 147774 220350
rect 147154 220226 147774 220294
rect 147154 220170 147250 220226
rect 147306 220170 147374 220226
rect 147430 220170 147498 220226
rect 147554 220170 147622 220226
rect 147678 220170 147774 220226
rect 147154 220102 147774 220170
rect 147154 220046 147250 220102
rect 147306 220046 147374 220102
rect 147430 220046 147498 220102
rect 147554 220046 147622 220102
rect 147678 220046 147774 220102
rect 147154 219978 147774 220046
rect 147154 219922 147250 219978
rect 147306 219922 147374 219978
rect 147430 219922 147498 219978
rect 147554 219922 147622 219978
rect 147678 219922 147774 219978
rect 147154 202350 147774 219922
rect 147154 202294 147250 202350
rect 147306 202294 147374 202350
rect 147430 202294 147498 202350
rect 147554 202294 147622 202350
rect 147678 202294 147774 202350
rect 147154 202226 147774 202294
rect 147154 202170 147250 202226
rect 147306 202170 147374 202226
rect 147430 202170 147498 202226
rect 147554 202170 147622 202226
rect 147678 202170 147774 202226
rect 147154 202102 147774 202170
rect 147154 202046 147250 202102
rect 147306 202046 147374 202102
rect 147430 202046 147498 202102
rect 147554 202046 147622 202102
rect 147678 202046 147774 202102
rect 147154 201978 147774 202046
rect 147154 201922 147250 201978
rect 147306 201922 147374 201978
rect 147430 201922 147498 201978
rect 147554 201922 147622 201978
rect 147678 201922 147774 201978
rect 147154 184350 147774 201922
rect 147154 184294 147250 184350
rect 147306 184294 147374 184350
rect 147430 184294 147498 184350
rect 147554 184294 147622 184350
rect 147678 184294 147774 184350
rect 147154 184226 147774 184294
rect 147154 184170 147250 184226
rect 147306 184170 147374 184226
rect 147430 184170 147498 184226
rect 147554 184170 147622 184226
rect 147678 184170 147774 184226
rect 147154 184102 147774 184170
rect 147154 184046 147250 184102
rect 147306 184046 147374 184102
rect 147430 184046 147498 184102
rect 147554 184046 147622 184102
rect 147678 184046 147774 184102
rect 147154 183978 147774 184046
rect 147154 183922 147250 183978
rect 147306 183922 147374 183978
rect 147430 183922 147498 183978
rect 147554 183922 147622 183978
rect 147678 183922 147774 183978
rect 147154 166350 147774 183922
rect 147154 166294 147250 166350
rect 147306 166294 147374 166350
rect 147430 166294 147498 166350
rect 147554 166294 147622 166350
rect 147678 166294 147774 166350
rect 147154 166226 147774 166294
rect 147154 166170 147250 166226
rect 147306 166170 147374 166226
rect 147430 166170 147498 166226
rect 147554 166170 147622 166226
rect 147678 166170 147774 166226
rect 147154 166102 147774 166170
rect 147154 166046 147250 166102
rect 147306 166046 147374 166102
rect 147430 166046 147498 166102
rect 147554 166046 147622 166102
rect 147678 166046 147774 166102
rect 147154 165978 147774 166046
rect 147154 165922 147250 165978
rect 147306 165922 147374 165978
rect 147430 165922 147498 165978
rect 147554 165922 147622 165978
rect 147678 165922 147774 165978
rect 147154 148350 147774 165922
rect 147154 148294 147250 148350
rect 147306 148294 147374 148350
rect 147430 148294 147498 148350
rect 147554 148294 147622 148350
rect 147678 148294 147774 148350
rect 147154 148226 147774 148294
rect 147154 148170 147250 148226
rect 147306 148170 147374 148226
rect 147430 148170 147498 148226
rect 147554 148170 147622 148226
rect 147678 148170 147774 148226
rect 147154 148102 147774 148170
rect 147154 148046 147250 148102
rect 147306 148046 147374 148102
rect 147430 148046 147498 148102
rect 147554 148046 147622 148102
rect 147678 148046 147774 148102
rect 147154 147978 147774 148046
rect 147154 147922 147250 147978
rect 147306 147922 147374 147978
rect 147430 147922 147498 147978
rect 147554 147922 147622 147978
rect 147678 147922 147774 147978
rect 147154 130350 147774 147922
rect 147154 130294 147250 130350
rect 147306 130294 147374 130350
rect 147430 130294 147498 130350
rect 147554 130294 147622 130350
rect 147678 130294 147774 130350
rect 147154 130226 147774 130294
rect 147154 130170 147250 130226
rect 147306 130170 147374 130226
rect 147430 130170 147498 130226
rect 147554 130170 147622 130226
rect 147678 130170 147774 130226
rect 147154 130102 147774 130170
rect 147154 130046 147250 130102
rect 147306 130046 147374 130102
rect 147430 130046 147498 130102
rect 147554 130046 147622 130102
rect 147678 130046 147774 130102
rect 147154 129978 147774 130046
rect 147154 129922 147250 129978
rect 147306 129922 147374 129978
rect 147430 129922 147498 129978
rect 147554 129922 147622 129978
rect 147678 129922 147774 129978
rect 147154 112350 147774 129922
rect 147154 112294 147250 112350
rect 147306 112294 147374 112350
rect 147430 112294 147498 112350
rect 147554 112294 147622 112350
rect 147678 112294 147774 112350
rect 147154 112226 147774 112294
rect 147154 112170 147250 112226
rect 147306 112170 147374 112226
rect 147430 112170 147498 112226
rect 147554 112170 147622 112226
rect 147678 112170 147774 112226
rect 147154 112102 147774 112170
rect 147154 112046 147250 112102
rect 147306 112046 147374 112102
rect 147430 112046 147498 112102
rect 147554 112046 147622 112102
rect 147678 112046 147774 112102
rect 147154 111978 147774 112046
rect 147154 111922 147250 111978
rect 147306 111922 147374 111978
rect 147430 111922 147498 111978
rect 147554 111922 147622 111978
rect 147678 111922 147774 111978
rect 147154 94350 147774 111922
rect 147154 94294 147250 94350
rect 147306 94294 147374 94350
rect 147430 94294 147498 94350
rect 147554 94294 147622 94350
rect 147678 94294 147774 94350
rect 147154 94226 147774 94294
rect 147154 94170 147250 94226
rect 147306 94170 147374 94226
rect 147430 94170 147498 94226
rect 147554 94170 147622 94226
rect 147678 94170 147774 94226
rect 147154 94102 147774 94170
rect 147154 94046 147250 94102
rect 147306 94046 147374 94102
rect 147430 94046 147498 94102
rect 147554 94046 147622 94102
rect 147678 94046 147774 94102
rect 147154 93978 147774 94046
rect 147154 93922 147250 93978
rect 147306 93922 147374 93978
rect 147430 93922 147498 93978
rect 147554 93922 147622 93978
rect 147678 93922 147774 93978
rect 147154 76350 147774 93922
rect 147154 76294 147250 76350
rect 147306 76294 147374 76350
rect 147430 76294 147498 76350
rect 147554 76294 147622 76350
rect 147678 76294 147774 76350
rect 147154 76226 147774 76294
rect 147154 76170 147250 76226
rect 147306 76170 147374 76226
rect 147430 76170 147498 76226
rect 147554 76170 147622 76226
rect 147678 76170 147774 76226
rect 147154 76102 147774 76170
rect 147154 76046 147250 76102
rect 147306 76046 147374 76102
rect 147430 76046 147498 76102
rect 147554 76046 147622 76102
rect 147678 76046 147774 76102
rect 147154 75978 147774 76046
rect 147154 75922 147250 75978
rect 147306 75922 147374 75978
rect 147430 75922 147498 75978
rect 147554 75922 147622 75978
rect 147678 75922 147774 75978
rect 147154 58350 147774 75922
rect 147154 58294 147250 58350
rect 147306 58294 147374 58350
rect 147430 58294 147498 58350
rect 147554 58294 147622 58350
rect 147678 58294 147774 58350
rect 147154 58226 147774 58294
rect 147154 58170 147250 58226
rect 147306 58170 147374 58226
rect 147430 58170 147498 58226
rect 147554 58170 147622 58226
rect 147678 58170 147774 58226
rect 147154 58102 147774 58170
rect 147154 58046 147250 58102
rect 147306 58046 147374 58102
rect 147430 58046 147498 58102
rect 147554 58046 147622 58102
rect 147678 58046 147774 58102
rect 147154 57978 147774 58046
rect 147154 57922 147250 57978
rect 147306 57922 147374 57978
rect 147430 57922 147498 57978
rect 147554 57922 147622 57978
rect 147678 57922 147774 57978
rect 147154 40350 147774 57922
rect 147154 40294 147250 40350
rect 147306 40294 147374 40350
rect 147430 40294 147498 40350
rect 147554 40294 147622 40350
rect 147678 40294 147774 40350
rect 147154 40226 147774 40294
rect 147154 40170 147250 40226
rect 147306 40170 147374 40226
rect 147430 40170 147498 40226
rect 147554 40170 147622 40226
rect 147678 40170 147774 40226
rect 147154 40102 147774 40170
rect 147154 40046 147250 40102
rect 147306 40046 147374 40102
rect 147430 40046 147498 40102
rect 147554 40046 147622 40102
rect 147678 40046 147774 40102
rect 147154 39978 147774 40046
rect 147154 39922 147250 39978
rect 147306 39922 147374 39978
rect 147430 39922 147498 39978
rect 147554 39922 147622 39978
rect 147678 39922 147774 39978
rect 147154 22350 147774 39922
rect 147154 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 147774 22350
rect 147154 22226 147774 22294
rect 147154 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 147774 22226
rect 147154 22102 147774 22170
rect 147154 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 147774 22102
rect 147154 21978 147774 22046
rect 147154 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 147774 21978
rect 147154 4350 147774 21922
rect 147154 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 147774 4350
rect 147154 4226 147774 4294
rect 147154 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 147774 4226
rect 147154 4102 147774 4170
rect 147154 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 147774 4102
rect 147154 3978 147774 4046
rect 147154 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 147774 3978
rect 147154 -160 147774 3922
rect 147154 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 147774 -160
rect 147154 -284 147774 -216
rect 147154 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 147774 -284
rect 147154 -408 147774 -340
rect 147154 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 147774 -408
rect 147154 -532 147774 -464
rect 147154 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 147774 -532
rect 147154 -1644 147774 -588
rect 150874 598172 151494 598268
rect 150874 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 151494 598172
rect 150874 598048 151494 598116
rect 150874 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 151494 598048
rect 150874 597924 151494 597992
rect 150874 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 151494 597924
rect 150874 597800 151494 597868
rect 150874 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 151494 597800
rect 150874 586350 151494 597744
rect 150874 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 151494 586350
rect 150874 586226 151494 586294
rect 150874 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 151494 586226
rect 150874 586102 151494 586170
rect 150874 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 151494 586102
rect 150874 585978 151494 586046
rect 150874 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 151494 585978
rect 150874 568350 151494 585922
rect 150874 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 151494 568350
rect 150874 568226 151494 568294
rect 150874 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 151494 568226
rect 150874 568102 151494 568170
rect 150874 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 151494 568102
rect 150874 567978 151494 568046
rect 150874 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 151494 567978
rect 150874 550350 151494 567922
rect 150874 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 151494 550350
rect 150874 550226 151494 550294
rect 150874 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 151494 550226
rect 150874 550102 151494 550170
rect 150874 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 151494 550102
rect 150874 549978 151494 550046
rect 150874 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 151494 549978
rect 150874 532350 151494 549922
rect 150874 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 151494 532350
rect 150874 532226 151494 532294
rect 150874 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 151494 532226
rect 150874 532102 151494 532170
rect 150874 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 151494 532102
rect 150874 531978 151494 532046
rect 150874 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 151494 531978
rect 150874 514350 151494 531922
rect 150874 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 151494 514350
rect 150874 514226 151494 514294
rect 150874 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 151494 514226
rect 150874 514102 151494 514170
rect 150874 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 151494 514102
rect 150874 513978 151494 514046
rect 150874 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 151494 513978
rect 150874 496350 151494 513922
rect 150874 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 151494 496350
rect 150874 496226 151494 496294
rect 150874 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 151494 496226
rect 150874 496102 151494 496170
rect 150874 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 151494 496102
rect 150874 495978 151494 496046
rect 150874 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 151494 495978
rect 150874 478350 151494 495922
rect 150874 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 151494 478350
rect 150874 478226 151494 478294
rect 150874 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 151494 478226
rect 150874 478102 151494 478170
rect 150874 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 151494 478102
rect 150874 477978 151494 478046
rect 150874 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 151494 477978
rect 150874 460350 151494 477922
rect 150874 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 151494 460350
rect 150874 460226 151494 460294
rect 150874 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 151494 460226
rect 150874 460102 151494 460170
rect 150874 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 151494 460102
rect 150874 459978 151494 460046
rect 150874 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 151494 459978
rect 150874 442350 151494 459922
rect 150874 442294 150970 442350
rect 151026 442294 151094 442350
rect 151150 442294 151218 442350
rect 151274 442294 151342 442350
rect 151398 442294 151494 442350
rect 150874 442226 151494 442294
rect 150874 442170 150970 442226
rect 151026 442170 151094 442226
rect 151150 442170 151218 442226
rect 151274 442170 151342 442226
rect 151398 442170 151494 442226
rect 150874 442102 151494 442170
rect 150874 442046 150970 442102
rect 151026 442046 151094 442102
rect 151150 442046 151218 442102
rect 151274 442046 151342 442102
rect 151398 442046 151494 442102
rect 150874 441978 151494 442046
rect 150874 441922 150970 441978
rect 151026 441922 151094 441978
rect 151150 441922 151218 441978
rect 151274 441922 151342 441978
rect 151398 441922 151494 441978
rect 150874 424350 151494 441922
rect 150874 424294 150970 424350
rect 151026 424294 151094 424350
rect 151150 424294 151218 424350
rect 151274 424294 151342 424350
rect 151398 424294 151494 424350
rect 150874 424226 151494 424294
rect 150874 424170 150970 424226
rect 151026 424170 151094 424226
rect 151150 424170 151218 424226
rect 151274 424170 151342 424226
rect 151398 424170 151494 424226
rect 150874 424102 151494 424170
rect 150874 424046 150970 424102
rect 151026 424046 151094 424102
rect 151150 424046 151218 424102
rect 151274 424046 151342 424102
rect 151398 424046 151494 424102
rect 150874 423978 151494 424046
rect 150874 423922 150970 423978
rect 151026 423922 151094 423978
rect 151150 423922 151218 423978
rect 151274 423922 151342 423978
rect 151398 423922 151494 423978
rect 150874 406350 151494 423922
rect 150874 406294 150970 406350
rect 151026 406294 151094 406350
rect 151150 406294 151218 406350
rect 151274 406294 151342 406350
rect 151398 406294 151494 406350
rect 150874 406226 151494 406294
rect 150874 406170 150970 406226
rect 151026 406170 151094 406226
rect 151150 406170 151218 406226
rect 151274 406170 151342 406226
rect 151398 406170 151494 406226
rect 150874 406102 151494 406170
rect 150874 406046 150970 406102
rect 151026 406046 151094 406102
rect 151150 406046 151218 406102
rect 151274 406046 151342 406102
rect 151398 406046 151494 406102
rect 150874 405978 151494 406046
rect 150874 405922 150970 405978
rect 151026 405922 151094 405978
rect 151150 405922 151218 405978
rect 151274 405922 151342 405978
rect 151398 405922 151494 405978
rect 150874 388350 151494 405922
rect 150874 388294 150970 388350
rect 151026 388294 151094 388350
rect 151150 388294 151218 388350
rect 151274 388294 151342 388350
rect 151398 388294 151494 388350
rect 150874 388226 151494 388294
rect 150874 388170 150970 388226
rect 151026 388170 151094 388226
rect 151150 388170 151218 388226
rect 151274 388170 151342 388226
rect 151398 388170 151494 388226
rect 150874 388102 151494 388170
rect 150874 388046 150970 388102
rect 151026 388046 151094 388102
rect 151150 388046 151218 388102
rect 151274 388046 151342 388102
rect 151398 388046 151494 388102
rect 150874 387978 151494 388046
rect 150874 387922 150970 387978
rect 151026 387922 151094 387978
rect 151150 387922 151218 387978
rect 151274 387922 151342 387978
rect 151398 387922 151494 387978
rect 150874 370350 151494 387922
rect 150874 370294 150970 370350
rect 151026 370294 151094 370350
rect 151150 370294 151218 370350
rect 151274 370294 151342 370350
rect 151398 370294 151494 370350
rect 150874 370226 151494 370294
rect 150874 370170 150970 370226
rect 151026 370170 151094 370226
rect 151150 370170 151218 370226
rect 151274 370170 151342 370226
rect 151398 370170 151494 370226
rect 150874 370102 151494 370170
rect 150874 370046 150970 370102
rect 151026 370046 151094 370102
rect 151150 370046 151218 370102
rect 151274 370046 151342 370102
rect 151398 370046 151494 370102
rect 150874 369978 151494 370046
rect 150874 369922 150970 369978
rect 151026 369922 151094 369978
rect 151150 369922 151218 369978
rect 151274 369922 151342 369978
rect 151398 369922 151494 369978
rect 150874 352350 151494 369922
rect 150874 352294 150970 352350
rect 151026 352294 151094 352350
rect 151150 352294 151218 352350
rect 151274 352294 151342 352350
rect 151398 352294 151494 352350
rect 150874 352226 151494 352294
rect 150874 352170 150970 352226
rect 151026 352170 151094 352226
rect 151150 352170 151218 352226
rect 151274 352170 151342 352226
rect 151398 352170 151494 352226
rect 150874 352102 151494 352170
rect 150874 352046 150970 352102
rect 151026 352046 151094 352102
rect 151150 352046 151218 352102
rect 151274 352046 151342 352102
rect 151398 352046 151494 352102
rect 150874 351978 151494 352046
rect 150874 351922 150970 351978
rect 151026 351922 151094 351978
rect 151150 351922 151218 351978
rect 151274 351922 151342 351978
rect 151398 351922 151494 351978
rect 150874 334350 151494 351922
rect 150874 334294 150970 334350
rect 151026 334294 151094 334350
rect 151150 334294 151218 334350
rect 151274 334294 151342 334350
rect 151398 334294 151494 334350
rect 150874 334226 151494 334294
rect 150874 334170 150970 334226
rect 151026 334170 151094 334226
rect 151150 334170 151218 334226
rect 151274 334170 151342 334226
rect 151398 334170 151494 334226
rect 150874 334102 151494 334170
rect 150874 334046 150970 334102
rect 151026 334046 151094 334102
rect 151150 334046 151218 334102
rect 151274 334046 151342 334102
rect 151398 334046 151494 334102
rect 150874 333978 151494 334046
rect 150874 333922 150970 333978
rect 151026 333922 151094 333978
rect 151150 333922 151218 333978
rect 151274 333922 151342 333978
rect 151398 333922 151494 333978
rect 150874 316350 151494 333922
rect 150874 316294 150970 316350
rect 151026 316294 151094 316350
rect 151150 316294 151218 316350
rect 151274 316294 151342 316350
rect 151398 316294 151494 316350
rect 150874 316226 151494 316294
rect 150874 316170 150970 316226
rect 151026 316170 151094 316226
rect 151150 316170 151218 316226
rect 151274 316170 151342 316226
rect 151398 316170 151494 316226
rect 150874 316102 151494 316170
rect 150874 316046 150970 316102
rect 151026 316046 151094 316102
rect 151150 316046 151218 316102
rect 151274 316046 151342 316102
rect 151398 316046 151494 316102
rect 150874 315978 151494 316046
rect 150874 315922 150970 315978
rect 151026 315922 151094 315978
rect 151150 315922 151218 315978
rect 151274 315922 151342 315978
rect 151398 315922 151494 315978
rect 150874 298350 151494 315922
rect 150874 298294 150970 298350
rect 151026 298294 151094 298350
rect 151150 298294 151218 298350
rect 151274 298294 151342 298350
rect 151398 298294 151494 298350
rect 150874 298226 151494 298294
rect 150874 298170 150970 298226
rect 151026 298170 151094 298226
rect 151150 298170 151218 298226
rect 151274 298170 151342 298226
rect 151398 298170 151494 298226
rect 150874 298102 151494 298170
rect 150874 298046 150970 298102
rect 151026 298046 151094 298102
rect 151150 298046 151218 298102
rect 151274 298046 151342 298102
rect 151398 298046 151494 298102
rect 150874 297978 151494 298046
rect 150874 297922 150970 297978
rect 151026 297922 151094 297978
rect 151150 297922 151218 297978
rect 151274 297922 151342 297978
rect 151398 297922 151494 297978
rect 150874 280350 151494 297922
rect 150874 280294 150970 280350
rect 151026 280294 151094 280350
rect 151150 280294 151218 280350
rect 151274 280294 151342 280350
rect 151398 280294 151494 280350
rect 150874 280226 151494 280294
rect 150874 280170 150970 280226
rect 151026 280170 151094 280226
rect 151150 280170 151218 280226
rect 151274 280170 151342 280226
rect 151398 280170 151494 280226
rect 150874 280102 151494 280170
rect 150874 280046 150970 280102
rect 151026 280046 151094 280102
rect 151150 280046 151218 280102
rect 151274 280046 151342 280102
rect 151398 280046 151494 280102
rect 150874 279978 151494 280046
rect 150874 279922 150970 279978
rect 151026 279922 151094 279978
rect 151150 279922 151218 279978
rect 151274 279922 151342 279978
rect 151398 279922 151494 279978
rect 150874 262350 151494 279922
rect 150874 262294 150970 262350
rect 151026 262294 151094 262350
rect 151150 262294 151218 262350
rect 151274 262294 151342 262350
rect 151398 262294 151494 262350
rect 150874 262226 151494 262294
rect 150874 262170 150970 262226
rect 151026 262170 151094 262226
rect 151150 262170 151218 262226
rect 151274 262170 151342 262226
rect 151398 262170 151494 262226
rect 150874 262102 151494 262170
rect 150874 262046 150970 262102
rect 151026 262046 151094 262102
rect 151150 262046 151218 262102
rect 151274 262046 151342 262102
rect 151398 262046 151494 262102
rect 150874 261978 151494 262046
rect 150874 261922 150970 261978
rect 151026 261922 151094 261978
rect 151150 261922 151218 261978
rect 151274 261922 151342 261978
rect 151398 261922 151494 261978
rect 150874 244350 151494 261922
rect 150874 244294 150970 244350
rect 151026 244294 151094 244350
rect 151150 244294 151218 244350
rect 151274 244294 151342 244350
rect 151398 244294 151494 244350
rect 150874 244226 151494 244294
rect 150874 244170 150970 244226
rect 151026 244170 151094 244226
rect 151150 244170 151218 244226
rect 151274 244170 151342 244226
rect 151398 244170 151494 244226
rect 150874 244102 151494 244170
rect 150874 244046 150970 244102
rect 151026 244046 151094 244102
rect 151150 244046 151218 244102
rect 151274 244046 151342 244102
rect 151398 244046 151494 244102
rect 150874 243978 151494 244046
rect 150874 243922 150970 243978
rect 151026 243922 151094 243978
rect 151150 243922 151218 243978
rect 151274 243922 151342 243978
rect 151398 243922 151494 243978
rect 150874 226350 151494 243922
rect 150874 226294 150970 226350
rect 151026 226294 151094 226350
rect 151150 226294 151218 226350
rect 151274 226294 151342 226350
rect 151398 226294 151494 226350
rect 150874 226226 151494 226294
rect 150874 226170 150970 226226
rect 151026 226170 151094 226226
rect 151150 226170 151218 226226
rect 151274 226170 151342 226226
rect 151398 226170 151494 226226
rect 150874 226102 151494 226170
rect 150874 226046 150970 226102
rect 151026 226046 151094 226102
rect 151150 226046 151218 226102
rect 151274 226046 151342 226102
rect 151398 226046 151494 226102
rect 150874 225978 151494 226046
rect 150874 225922 150970 225978
rect 151026 225922 151094 225978
rect 151150 225922 151218 225978
rect 151274 225922 151342 225978
rect 151398 225922 151494 225978
rect 150874 208350 151494 225922
rect 150874 208294 150970 208350
rect 151026 208294 151094 208350
rect 151150 208294 151218 208350
rect 151274 208294 151342 208350
rect 151398 208294 151494 208350
rect 150874 208226 151494 208294
rect 150874 208170 150970 208226
rect 151026 208170 151094 208226
rect 151150 208170 151218 208226
rect 151274 208170 151342 208226
rect 151398 208170 151494 208226
rect 150874 208102 151494 208170
rect 150874 208046 150970 208102
rect 151026 208046 151094 208102
rect 151150 208046 151218 208102
rect 151274 208046 151342 208102
rect 151398 208046 151494 208102
rect 150874 207978 151494 208046
rect 150874 207922 150970 207978
rect 151026 207922 151094 207978
rect 151150 207922 151218 207978
rect 151274 207922 151342 207978
rect 151398 207922 151494 207978
rect 150874 190350 151494 207922
rect 150874 190294 150970 190350
rect 151026 190294 151094 190350
rect 151150 190294 151218 190350
rect 151274 190294 151342 190350
rect 151398 190294 151494 190350
rect 150874 190226 151494 190294
rect 150874 190170 150970 190226
rect 151026 190170 151094 190226
rect 151150 190170 151218 190226
rect 151274 190170 151342 190226
rect 151398 190170 151494 190226
rect 150874 190102 151494 190170
rect 150874 190046 150970 190102
rect 151026 190046 151094 190102
rect 151150 190046 151218 190102
rect 151274 190046 151342 190102
rect 151398 190046 151494 190102
rect 150874 189978 151494 190046
rect 150874 189922 150970 189978
rect 151026 189922 151094 189978
rect 151150 189922 151218 189978
rect 151274 189922 151342 189978
rect 151398 189922 151494 189978
rect 150874 172350 151494 189922
rect 150874 172294 150970 172350
rect 151026 172294 151094 172350
rect 151150 172294 151218 172350
rect 151274 172294 151342 172350
rect 151398 172294 151494 172350
rect 150874 172226 151494 172294
rect 150874 172170 150970 172226
rect 151026 172170 151094 172226
rect 151150 172170 151218 172226
rect 151274 172170 151342 172226
rect 151398 172170 151494 172226
rect 150874 172102 151494 172170
rect 150874 172046 150970 172102
rect 151026 172046 151094 172102
rect 151150 172046 151218 172102
rect 151274 172046 151342 172102
rect 151398 172046 151494 172102
rect 150874 171978 151494 172046
rect 150874 171922 150970 171978
rect 151026 171922 151094 171978
rect 151150 171922 151218 171978
rect 151274 171922 151342 171978
rect 151398 171922 151494 171978
rect 150874 154350 151494 171922
rect 150874 154294 150970 154350
rect 151026 154294 151094 154350
rect 151150 154294 151218 154350
rect 151274 154294 151342 154350
rect 151398 154294 151494 154350
rect 150874 154226 151494 154294
rect 150874 154170 150970 154226
rect 151026 154170 151094 154226
rect 151150 154170 151218 154226
rect 151274 154170 151342 154226
rect 151398 154170 151494 154226
rect 150874 154102 151494 154170
rect 150874 154046 150970 154102
rect 151026 154046 151094 154102
rect 151150 154046 151218 154102
rect 151274 154046 151342 154102
rect 151398 154046 151494 154102
rect 150874 153978 151494 154046
rect 150874 153922 150970 153978
rect 151026 153922 151094 153978
rect 151150 153922 151218 153978
rect 151274 153922 151342 153978
rect 151398 153922 151494 153978
rect 150874 136350 151494 153922
rect 150874 136294 150970 136350
rect 151026 136294 151094 136350
rect 151150 136294 151218 136350
rect 151274 136294 151342 136350
rect 151398 136294 151494 136350
rect 150874 136226 151494 136294
rect 150874 136170 150970 136226
rect 151026 136170 151094 136226
rect 151150 136170 151218 136226
rect 151274 136170 151342 136226
rect 151398 136170 151494 136226
rect 150874 136102 151494 136170
rect 150874 136046 150970 136102
rect 151026 136046 151094 136102
rect 151150 136046 151218 136102
rect 151274 136046 151342 136102
rect 151398 136046 151494 136102
rect 150874 135978 151494 136046
rect 150874 135922 150970 135978
rect 151026 135922 151094 135978
rect 151150 135922 151218 135978
rect 151274 135922 151342 135978
rect 151398 135922 151494 135978
rect 150874 118350 151494 135922
rect 150874 118294 150970 118350
rect 151026 118294 151094 118350
rect 151150 118294 151218 118350
rect 151274 118294 151342 118350
rect 151398 118294 151494 118350
rect 150874 118226 151494 118294
rect 150874 118170 150970 118226
rect 151026 118170 151094 118226
rect 151150 118170 151218 118226
rect 151274 118170 151342 118226
rect 151398 118170 151494 118226
rect 150874 118102 151494 118170
rect 150874 118046 150970 118102
rect 151026 118046 151094 118102
rect 151150 118046 151218 118102
rect 151274 118046 151342 118102
rect 151398 118046 151494 118102
rect 150874 117978 151494 118046
rect 150874 117922 150970 117978
rect 151026 117922 151094 117978
rect 151150 117922 151218 117978
rect 151274 117922 151342 117978
rect 151398 117922 151494 117978
rect 150874 100350 151494 117922
rect 150874 100294 150970 100350
rect 151026 100294 151094 100350
rect 151150 100294 151218 100350
rect 151274 100294 151342 100350
rect 151398 100294 151494 100350
rect 150874 100226 151494 100294
rect 150874 100170 150970 100226
rect 151026 100170 151094 100226
rect 151150 100170 151218 100226
rect 151274 100170 151342 100226
rect 151398 100170 151494 100226
rect 150874 100102 151494 100170
rect 150874 100046 150970 100102
rect 151026 100046 151094 100102
rect 151150 100046 151218 100102
rect 151274 100046 151342 100102
rect 151398 100046 151494 100102
rect 150874 99978 151494 100046
rect 150874 99922 150970 99978
rect 151026 99922 151094 99978
rect 151150 99922 151218 99978
rect 151274 99922 151342 99978
rect 151398 99922 151494 99978
rect 150874 82350 151494 99922
rect 150874 82294 150970 82350
rect 151026 82294 151094 82350
rect 151150 82294 151218 82350
rect 151274 82294 151342 82350
rect 151398 82294 151494 82350
rect 150874 82226 151494 82294
rect 150874 82170 150970 82226
rect 151026 82170 151094 82226
rect 151150 82170 151218 82226
rect 151274 82170 151342 82226
rect 151398 82170 151494 82226
rect 150874 82102 151494 82170
rect 150874 82046 150970 82102
rect 151026 82046 151094 82102
rect 151150 82046 151218 82102
rect 151274 82046 151342 82102
rect 151398 82046 151494 82102
rect 150874 81978 151494 82046
rect 150874 81922 150970 81978
rect 151026 81922 151094 81978
rect 151150 81922 151218 81978
rect 151274 81922 151342 81978
rect 151398 81922 151494 81978
rect 150874 64350 151494 81922
rect 150874 64294 150970 64350
rect 151026 64294 151094 64350
rect 151150 64294 151218 64350
rect 151274 64294 151342 64350
rect 151398 64294 151494 64350
rect 150874 64226 151494 64294
rect 150874 64170 150970 64226
rect 151026 64170 151094 64226
rect 151150 64170 151218 64226
rect 151274 64170 151342 64226
rect 151398 64170 151494 64226
rect 150874 64102 151494 64170
rect 150874 64046 150970 64102
rect 151026 64046 151094 64102
rect 151150 64046 151218 64102
rect 151274 64046 151342 64102
rect 151398 64046 151494 64102
rect 150874 63978 151494 64046
rect 150874 63922 150970 63978
rect 151026 63922 151094 63978
rect 151150 63922 151218 63978
rect 151274 63922 151342 63978
rect 151398 63922 151494 63978
rect 150874 46350 151494 63922
rect 150874 46294 150970 46350
rect 151026 46294 151094 46350
rect 151150 46294 151218 46350
rect 151274 46294 151342 46350
rect 151398 46294 151494 46350
rect 150874 46226 151494 46294
rect 150874 46170 150970 46226
rect 151026 46170 151094 46226
rect 151150 46170 151218 46226
rect 151274 46170 151342 46226
rect 151398 46170 151494 46226
rect 150874 46102 151494 46170
rect 150874 46046 150970 46102
rect 151026 46046 151094 46102
rect 151150 46046 151218 46102
rect 151274 46046 151342 46102
rect 151398 46046 151494 46102
rect 150874 45978 151494 46046
rect 150874 45922 150970 45978
rect 151026 45922 151094 45978
rect 151150 45922 151218 45978
rect 151274 45922 151342 45978
rect 151398 45922 151494 45978
rect 150874 28350 151494 45922
rect 150874 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 151494 28350
rect 150874 28226 151494 28294
rect 150874 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 151494 28226
rect 150874 28102 151494 28170
rect 150874 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 151494 28102
rect 150874 27978 151494 28046
rect 150874 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 151494 27978
rect 150874 10350 151494 27922
rect 150874 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 151494 10350
rect 150874 10226 151494 10294
rect 150874 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 151494 10226
rect 150874 10102 151494 10170
rect 150874 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 151494 10102
rect 150874 9978 151494 10046
rect 150874 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 151494 9978
rect 150874 -1120 151494 9922
rect 150874 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 151494 -1120
rect 150874 -1244 151494 -1176
rect 150874 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 151494 -1244
rect 150874 -1368 151494 -1300
rect 150874 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 151494 -1368
rect 150874 -1492 151494 -1424
rect 150874 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 151494 -1492
rect 150874 -1644 151494 -1548
rect 165154 597212 165774 598268
rect 165154 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 165774 597212
rect 165154 597088 165774 597156
rect 165154 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 165774 597088
rect 165154 596964 165774 597032
rect 165154 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 165774 596964
rect 165154 596840 165774 596908
rect 165154 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 165774 596840
rect 165154 580350 165774 596784
rect 165154 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 165774 580350
rect 165154 580226 165774 580294
rect 165154 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 165774 580226
rect 165154 580102 165774 580170
rect 165154 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 165774 580102
rect 165154 579978 165774 580046
rect 165154 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 165774 579978
rect 165154 562350 165774 579922
rect 165154 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 165774 562350
rect 165154 562226 165774 562294
rect 165154 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 165774 562226
rect 165154 562102 165774 562170
rect 165154 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 165774 562102
rect 165154 561978 165774 562046
rect 165154 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 165774 561978
rect 165154 544350 165774 561922
rect 165154 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 165774 544350
rect 165154 544226 165774 544294
rect 165154 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 165774 544226
rect 165154 544102 165774 544170
rect 165154 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 165774 544102
rect 165154 543978 165774 544046
rect 165154 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 165774 543978
rect 165154 526350 165774 543922
rect 165154 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 165774 526350
rect 165154 526226 165774 526294
rect 165154 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 165774 526226
rect 165154 526102 165774 526170
rect 165154 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 165774 526102
rect 165154 525978 165774 526046
rect 165154 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 165774 525978
rect 165154 508350 165774 525922
rect 165154 508294 165250 508350
rect 165306 508294 165374 508350
rect 165430 508294 165498 508350
rect 165554 508294 165622 508350
rect 165678 508294 165774 508350
rect 165154 508226 165774 508294
rect 165154 508170 165250 508226
rect 165306 508170 165374 508226
rect 165430 508170 165498 508226
rect 165554 508170 165622 508226
rect 165678 508170 165774 508226
rect 165154 508102 165774 508170
rect 165154 508046 165250 508102
rect 165306 508046 165374 508102
rect 165430 508046 165498 508102
rect 165554 508046 165622 508102
rect 165678 508046 165774 508102
rect 165154 507978 165774 508046
rect 165154 507922 165250 507978
rect 165306 507922 165374 507978
rect 165430 507922 165498 507978
rect 165554 507922 165622 507978
rect 165678 507922 165774 507978
rect 165154 490350 165774 507922
rect 165154 490294 165250 490350
rect 165306 490294 165374 490350
rect 165430 490294 165498 490350
rect 165554 490294 165622 490350
rect 165678 490294 165774 490350
rect 165154 490226 165774 490294
rect 165154 490170 165250 490226
rect 165306 490170 165374 490226
rect 165430 490170 165498 490226
rect 165554 490170 165622 490226
rect 165678 490170 165774 490226
rect 165154 490102 165774 490170
rect 165154 490046 165250 490102
rect 165306 490046 165374 490102
rect 165430 490046 165498 490102
rect 165554 490046 165622 490102
rect 165678 490046 165774 490102
rect 165154 489978 165774 490046
rect 165154 489922 165250 489978
rect 165306 489922 165374 489978
rect 165430 489922 165498 489978
rect 165554 489922 165622 489978
rect 165678 489922 165774 489978
rect 165154 472350 165774 489922
rect 165154 472294 165250 472350
rect 165306 472294 165374 472350
rect 165430 472294 165498 472350
rect 165554 472294 165622 472350
rect 165678 472294 165774 472350
rect 165154 472226 165774 472294
rect 165154 472170 165250 472226
rect 165306 472170 165374 472226
rect 165430 472170 165498 472226
rect 165554 472170 165622 472226
rect 165678 472170 165774 472226
rect 165154 472102 165774 472170
rect 165154 472046 165250 472102
rect 165306 472046 165374 472102
rect 165430 472046 165498 472102
rect 165554 472046 165622 472102
rect 165678 472046 165774 472102
rect 165154 471978 165774 472046
rect 165154 471922 165250 471978
rect 165306 471922 165374 471978
rect 165430 471922 165498 471978
rect 165554 471922 165622 471978
rect 165678 471922 165774 471978
rect 165154 454350 165774 471922
rect 165154 454294 165250 454350
rect 165306 454294 165374 454350
rect 165430 454294 165498 454350
rect 165554 454294 165622 454350
rect 165678 454294 165774 454350
rect 165154 454226 165774 454294
rect 165154 454170 165250 454226
rect 165306 454170 165374 454226
rect 165430 454170 165498 454226
rect 165554 454170 165622 454226
rect 165678 454170 165774 454226
rect 165154 454102 165774 454170
rect 165154 454046 165250 454102
rect 165306 454046 165374 454102
rect 165430 454046 165498 454102
rect 165554 454046 165622 454102
rect 165678 454046 165774 454102
rect 165154 453978 165774 454046
rect 165154 453922 165250 453978
rect 165306 453922 165374 453978
rect 165430 453922 165498 453978
rect 165554 453922 165622 453978
rect 165678 453922 165774 453978
rect 165154 436350 165774 453922
rect 165154 436294 165250 436350
rect 165306 436294 165374 436350
rect 165430 436294 165498 436350
rect 165554 436294 165622 436350
rect 165678 436294 165774 436350
rect 165154 436226 165774 436294
rect 165154 436170 165250 436226
rect 165306 436170 165374 436226
rect 165430 436170 165498 436226
rect 165554 436170 165622 436226
rect 165678 436170 165774 436226
rect 165154 436102 165774 436170
rect 165154 436046 165250 436102
rect 165306 436046 165374 436102
rect 165430 436046 165498 436102
rect 165554 436046 165622 436102
rect 165678 436046 165774 436102
rect 165154 435978 165774 436046
rect 165154 435922 165250 435978
rect 165306 435922 165374 435978
rect 165430 435922 165498 435978
rect 165554 435922 165622 435978
rect 165678 435922 165774 435978
rect 165154 418350 165774 435922
rect 165154 418294 165250 418350
rect 165306 418294 165374 418350
rect 165430 418294 165498 418350
rect 165554 418294 165622 418350
rect 165678 418294 165774 418350
rect 165154 418226 165774 418294
rect 165154 418170 165250 418226
rect 165306 418170 165374 418226
rect 165430 418170 165498 418226
rect 165554 418170 165622 418226
rect 165678 418170 165774 418226
rect 165154 418102 165774 418170
rect 165154 418046 165250 418102
rect 165306 418046 165374 418102
rect 165430 418046 165498 418102
rect 165554 418046 165622 418102
rect 165678 418046 165774 418102
rect 165154 417978 165774 418046
rect 165154 417922 165250 417978
rect 165306 417922 165374 417978
rect 165430 417922 165498 417978
rect 165554 417922 165622 417978
rect 165678 417922 165774 417978
rect 165154 400350 165774 417922
rect 165154 400294 165250 400350
rect 165306 400294 165374 400350
rect 165430 400294 165498 400350
rect 165554 400294 165622 400350
rect 165678 400294 165774 400350
rect 165154 400226 165774 400294
rect 165154 400170 165250 400226
rect 165306 400170 165374 400226
rect 165430 400170 165498 400226
rect 165554 400170 165622 400226
rect 165678 400170 165774 400226
rect 165154 400102 165774 400170
rect 165154 400046 165250 400102
rect 165306 400046 165374 400102
rect 165430 400046 165498 400102
rect 165554 400046 165622 400102
rect 165678 400046 165774 400102
rect 165154 399978 165774 400046
rect 165154 399922 165250 399978
rect 165306 399922 165374 399978
rect 165430 399922 165498 399978
rect 165554 399922 165622 399978
rect 165678 399922 165774 399978
rect 165154 382350 165774 399922
rect 165154 382294 165250 382350
rect 165306 382294 165374 382350
rect 165430 382294 165498 382350
rect 165554 382294 165622 382350
rect 165678 382294 165774 382350
rect 165154 382226 165774 382294
rect 165154 382170 165250 382226
rect 165306 382170 165374 382226
rect 165430 382170 165498 382226
rect 165554 382170 165622 382226
rect 165678 382170 165774 382226
rect 165154 382102 165774 382170
rect 165154 382046 165250 382102
rect 165306 382046 165374 382102
rect 165430 382046 165498 382102
rect 165554 382046 165622 382102
rect 165678 382046 165774 382102
rect 165154 381978 165774 382046
rect 165154 381922 165250 381978
rect 165306 381922 165374 381978
rect 165430 381922 165498 381978
rect 165554 381922 165622 381978
rect 165678 381922 165774 381978
rect 165154 364350 165774 381922
rect 165154 364294 165250 364350
rect 165306 364294 165374 364350
rect 165430 364294 165498 364350
rect 165554 364294 165622 364350
rect 165678 364294 165774 364350
rect 165154 364226 165774 364294
rect 165154 364170 165250 364226
rect 165306 364170 165374 364226
rect 165430 364170 165498 364226
rect 165554 364170 165622 364226
rect 165678 364170 165774 364226
rect 165154 364102 165774 364170
rect 165154 364046 165250 364102
rect 165306 364046 165374 364102
rect 165430 364046 165498 364102
rect 165554 364046 165622 364102
rect 165678 364046 165774 364102
rect 165154 363978 165774 364046
rect 165154 363922 165250 363978
rect 165306 363922 165374 363978
rect 165430 363922 165498 363978
rect 165554 363922 165622 363978
rect 165678 363922 165774 363978
rect 165154 346350 165774 363922
rect 165154 346294 165250 346350
rect 165306 346294 165374 346350
rect 165430 346294 165498 346350
rect 165554 346294 165622 346350
rect 165678 346294 165774 346350
rect 165154 346226 165774 346294
rect 165154 346170 165250 346226
rect 165306 346170 165374 346226
rect 165430 346170 165498 346226
rect 165554 346170 165622 346226
rect 165678 346170 165774 346226
rect 165154 346102 165774 346170
rect 165154 346046 165250 346102
rect 165306 346046 165374 346102
rect 165430 346046 165498 346102
rect 165554 346046 165622 346102
rect 165678 346046 165774 346102
rect 165154 345978 165774 346046
rect 165154 345922 165250 345978
rect 165306 345922 165374 345978
rect 165430 345922 165498 345978
rect 165554 345922 165622 345978
rect 165678 345922 165774 345978
rect 165154 328350 165774 345922
rect 165154 328294 165250 328350
rect 165306 328294 165374 328350
rect 165430 328294 165498 328350
rect 165554 328294 165622 328350
rect 165678 328294 165774 328350
rect 165154 328226 165774 328294
rect 165154 328170 165250 328226
rect 165306 328170 165374 328226
rect 165430 328170 165498 328226
rect 165554 328170 165622 328226
rect 165678 328170 165774 328226
rect 165154 328102 165774 328170
rect 165154 328046 165250 328102
rect 165306 328046 165374 328102
rect 165430 328046 165498 328102
rect 165554 328046 165622 328102
rect 165678 328046 165774 328102
rect 165154 327978 165774 328046
rect 165154 327922 165250 327978
rect 165306 327922 165374 327978
rect 165430 327922 165498 327978
rect 165554 327922 165622 327978
rect 165678 327922 165774 327978
rect 165154 310350 165774 327922
rect 165154 310294 165250 310350
rect 165306 310294 165374 310350
rect 165430 310294 165498 310350
rect 165554 310294 165622 310350
rect 165678 310294 165774 310350
rect 165154 310226 165774 310294
rect 165154 310170 165250 310226
rect 165306 310170 165374 310226
rect 165430 310170 165498 310226
rect 165554 310170 165622 310226
rect 165678 310170 165774 310226
rect 165154 310102 165774 310170
rect 165154 310046 165250 310102
rect 165306 310046 165374 310102
rect 165430 310046 165498 310102
rect 165554 310046 165622 310102
rect 165678 310046 165774 310102
rect 165154 309978 165774 310046
rect 165154 309922 165250 309978
rect 165306 309922 165374 309978
rect 165430 309922 165498 309978
rect 165554 309922 165622 309978
rect 165678 309922 165774 309978
rect 165154 292350 165774 309922
rect 165154 292294 165250 292350
rect 165306 292294 165374 292350
rect 165430 292294 165498 292350
rect 165554 292294 165622 292350
rect 165678 292294 165774 292350
rect 165154 292226 165774 292294
rect 165154 292170 165250 292226
rect 165306 292170 165374 292226
rect 165430 292170 165498 292226
rect 165554 292170 165622 292226
rect 165678 292170 165774 292226
rect 165154 292102 165774 292170
rect 165154 292046 165250 292102
rect 165306 292046 165374 292102
rect 165430 292046 165498 292102
rect 165554 292046 165622 292102
rect 165678 292046 165774 292102
rect 165154 291978 165774 292046
rect 165154 291922 165250 291978
rect 165306 291922 165374 291978
rect 165430 291922 165498 291978
rect 165554 291922 165622 291978
rect 165678 291922 165774 291978
rect 165154 274350 165774 291922
rect 165154 274294 165250 274350
rect 165306 274294 165374 274350
rect 165430 274294 165498 274350
rect 165554 274294 165622 274350
rect 165678 274294 165774 274350
rect 165154 274226 165774 274294
rect 165154 274170 165250 274226
rect 165306 274170 165374 274226
rect 165430 274170 165498 274226
rect 165554 274170 165622 274226
rect 165678 274170 165774 274226
rect 165154 274102 165774 274170
rect 165154 274046 165250 274102
rect 165306 274046 165374 274102
rect 165430 274046 165498 274102
rect 165554 274046 165622 274102
rect 165678 274046 165774 274102
rect 165154 273978 165774 274046
rect 165154 273922 165250 273978
rect 165306 273922 165374 273978
rect 165430 273922 165498 273978
rect 165554 273922 165622 273978
rect 165678 273922 165774 273978
rect 165154 256350 165774 273922
rect 165154 256294 165250 256350
rect 165306 256294 165374 256350
rect 165430 256294 165498 256350
rect 165554 256294 165622 256350
rect 165678 256294 165774 256350
rect 165154 256226 165774 256294
rect 165154 256170 165250 256226
rect 165306 256170 165374 256226
rect 165430 256170 165498 256226
rect 165554 256170 165622 256226
rect 165678 256170 165774 256226
rect 165154 256102 165774 256170
rect 165154 256046 165250 256102
rect 165306 256046 165374 256102
rect 165430 256046 165498 256102
rect 165554 256046 165622 256102
rect 165678 256046 165774 256102
rect 165154 255978 165774 256046
rect 165154 255922 165250 255978
rect 165306 255922 165374 255978
rect 165430 255922 165498 255978
rect 165554 255922 165622 255978
rect 165678 255922 165774 255978
rect 165154 238350 165774 255922
rect 165154 238294 165250 238350
rect 165306 238294 165374 238350
rect 165430 238294 165498 238350
rect 165554 238294 165622 238350
rect 165678 238294 165774 238350
rect 165154 238226 165774 238294
rect 165154 238170 165250 238226
rect 165306 238170 165374 238226
rect 165430 238170 165498 238226
rect 165554 238170 165622 238226
rect 165678 238170 165774 238226
rect 165154 238102 165774 238170
rect 165154 238046 165250 238102
rect 165306 238046 165374 238102
rect 165430 238046 165498 238102
rect 165554 238046 165622 238102
rect 165678 238046 165774 238102
rect 165154 237978 165774 238046
rect 165154 237922 165250 237978
rect 165306 237922 165374 237978
rect 165430 237922 165498 237978
rect 165554 237922 165622 237978
rect 165678 237922 165774 237978
rect 165154 220350 165774 237922
rect 165154 220294 165250 220350
rect 165306 220294 165374 220350
rect 165430 220294 165498 220350
rect 165554 220294 165622 220350
rect 165678 220294 165774 220350
rect 165154 220226 165774 220294
rect 165154 220170 165250 220226
rect 165306 220170 165374 220226
rect 165430 220170 165498 220226
rect 165554 220170 165622 220226
rect 165678 220170 165774 220226
rect 165154 220102 165774 220170
rect 165154 220046 165250 220102
rect 165306 220046 165374 220102
rect 165430 220046 165498 220102
rect 165554 220046 165622 220102
rect 165678 220046 165774 220102
rect 165154 219978 165774 220046
rect 165154 219922 165250 219978
rect 165306 219922 165374 219978
rect 165430 219922 165498 219978
rect 165554 219922 165622 219978
rect 165678 219922 165774 219978
rect 165154 202350 165774 219922
rect 165154 202294 165250 202350
rect 165306 202294 165374 202350
rect 165430 202294 165498 202350
rect 165554 202294 165622 202350
rect 165678 202294 165774 202350
rect 165154 202226 165774 202294
rect 165154 202170 165250 202226
rect 165306 202170 165374 202226
rect 165430 202170 165498 202226
rect 165554 202170 165622 202226
rect 165678 202170 165774 202226
rect 165154 202102 165774 202170
rect 165154 202046 165250 202102
rect 165306 202046 165374 202102
rect 165430 202046 165498 202102
rect 165554 202046 165622 202102
rect 165678 202046 165774 202102
rect 165154 201978 165774 202046
rect 165154 201922 165250 201978
rect 165306 201922 165374 201978
rect 165430 201922 165498 201978
rect 165554 201922 165622 201978
rect 165678 201922 165774 201978
rect 165154 184350 165774 201922
rect 165154 184294 165250 184350
rect 165306 184294 165374 184350
rect 165430 184294 165498 184350
rect 165554 184294 165622 184350
rect 165678 184294 165774 184350
rect 165154 184226 165774 184294
rect 165154 184170 165250 184226
rect 165306 184170 165374 184226
rect 165430 184170 165498 184226
rect 165554 184170 165622 184226
rect 165678 184170 165774 184226
rect 165154 184102 165774 184170
rect 165154 184046 165250 184102
rect 165306 184046 165374 184102
rect 165430 184046 165498 184102
rect 165554 184046 165622 184102
rect 165678 184046 165774 184102
rect 165154 183978 165774 184046
rect 165154 183922 165250 183978
rect 165306 183922 165374 183978
rect 165430 183922 165498 183978
rect 165554 183922 165622 183978
rect 165678 183922 165774 183978
rect 165154 166350 165774 183922
rect 165154 166294 165250 166350
rect 165306 166294 165374 166350
rect 165430 166294 165498 166350
rect 165554 166294 165622 166350
rect 165678 166294 165774 166350
rect 165154 166226 165774 166294
rect 165154 166170 165250 166226
rect 165306 166170 165374 166226
rect 165430 166170 165498 166226
rect 165554 166170 165622 166226
rect 165678 166170 165774 166226
rect 165154 166102 165774 166170
rect 165154 166046 165250 166102
rect 165306 166046 165374 166102
rect 165430 166046 165498 166102
rect 165554 166046 165622 166102
rect 165678 166046 165774 166102
rect 165154 165978 165774 166046
rect 165154 165922 165250 165978
rect 165306 165922 165374 165978
rect 165430 165922 165498 165978
rect 165554 165922 165622 165978
rect 165678 165922 165774 165978
rect 165154 148350 165774 165922
rect 165154 148294 165250 148350
rect 165306 148294 165374 148350
rect 165430 148294 165498 148350
rect 165554 148294 165622 148350
rect 165678 148294 165774 148350
rect 165154 148226 165774 148294
rect 165154 148170 165250 148226
rect 165306 148170 165374 148226
rect 165430 148170 165498 148226
rect 165554 148170 165622 148226
rect 165678 148170 165774 148226
rect 165154 148102 165774 148170
rect 165154 148046 165250 148102
rect 165306 148046 165374 148102
rect 165430 148046 165498 148102
rect 165554 148046 165622 148102
rect 165678 148046 165774 148102
rect 165154 147978 165774 148046
rect 165154 147922 165250 147978
rect 165306 147922 165374 147978
rect 165430 147922 165498 147978
rect 165554 147922 165622 147978
rect 165678 147922 165774 147978
rect 165154 130350 165774 147922
rect 165154 130294 165250 130350
rect 165306 130294 165374 130350
rect 165430 130294 165498 130350
rect 165554 130294 165622 130350
rect 165678 130294 165774 130350
rect 165154 130226 165774 130294
rect 165154 130170 165250 130226
rect 165306 130170 165374 130226
rect 165430 130170 165498 130226
rect 165554 130170 165622 130226
rect 165678 130170 165774 130226
rect 165154 130102 165774 130170
rect 165154 130046 165250 130102
rect 165306 130046 165374 130102
rect 165430 130046 165498 130102
rect 165554 130046 165622 130102
rect 165678 130046 165774 130102
rect 165154 129978 165774 130046
rect 165154 129922 165250 129978
rect 165306 129922 165374 129978
rect 165430 129922 165498 129978
rect 165554 129922 165622 129978
rect 165678 129922 165774 129978
rect 165154 112350 165774 129922
rect 165154 112294 165250 112350
rect 165306 112294 165374 112350
rect 165430 112294 165498 112350
rect 165554 112294 165622 112350
rect 165678 112294 165774 112350
rect 165154 112226 165774 112294
rect 165154 112170 165250 112226
rect 165306 112170 165374 112226
rect 165430 112170 165498 112226
rect 165554 112170 165622 112226
rect 165678 112170 165774 112226
rect 165154 112102 165774 112170
rect 165154 112046 165250 112102
rect 165306 112046 165374 112102
rect 165430 112046 165498 112102
rect 165554 112046 165622 112102
rect 165678 112046 165774 112102
rect 165154 111978 165774 112046
rect 165154 111922 165250 111978
rect 165306 111922 165374 111978
rect 165430 111922 165498 111978
rect 165554 111922 165622 111978
rect 165678 111922 165774 111978
rect 165154 94350 165774 111922
rect 165154 94294 165250 94350
rect 165306 94294 165374 94350
rect 165430 94294 165498 94350
rect 165554 94294 165622 94350
rect 165678 94294 165774 94350
rect 165154 94226 165774 94294
rect 165154 94170 165250 94226
rect 165306 94170 165374 94226
rect 165430 94170 165498 94226
rect 165554 94170 165622 94226
rect 165678 94170 165774 94226
rect 165154 94102 165774 94170
rect 165154 94046 165250 94102
rect 165306 94046 165374 94102
rect 165430 94046 165498 94102
rect 165554 94046 165622 94102
rect 165678 94046 165774 94102
rect 165154 93978 165774 94046
rect 165154 93922 165250 93978
rect 165306 93922 165374 93978
rect 165430 93922 165498 93978
rect 165554 93922 165622 93978
rect 165678 93922 165774 93978
rect 165154 76350 165774 93922
rect 165154 76294 165250 76350
rect 165306 76294 165374 76350
rect 165430 76294 165498 76350
rect 165554 76294 165622 76350
rect 165678 76294 165774 76350
rect 165154 76226 165774 76294
rect 165154 76170 165250 76226
rect 165306 76170 165374 76226
rect 165430 76170 165498 76226
rect 165554 76170 165622 76226
rect 165678 76170 165774 76226
rect 165154 76102 165774 76170
rect 165154 76046 165250 76102
rect 165306 76046 165374 76102
rect 165430 76046 165498 76102
rect 165554 76046 165622 76102
rect 165678 76046 165774 76102
rect 165154 75978 165774 76046
rect 165154 75922 165250 75978
rect 165306 75922 165374 75978
rect 165430 75922 165498 75978
rect 165554 75922 165622 75978
rect 165678 75922 165774 75978
rect 165154 58350 165774 75922
rect 165154 58294 165250 58350
rect 165306 58294 165374 58350
rect 165430 58294 165498 58350
rect 165554 58294 165622 58350
rect 165678 58294 165774 58350
rect 165154 58226 165774 58294
rect 165154 58170 165250 58226
rect 165306 58170 165374 58226
rect 165430 58170 165498 58226
rect 165554 58170 165622 58226
rect 165678 58170 165774 58226
rect 165154 58102 165774 58170
rect 165154 58046 165250 58102
rect 165306 58046 165374 58102
rect 165430 58046 165498 58102
rect 165554 58046 165622 58102
rect 165678 58046 165774 58102
rect 165154 57978 165774 58046
rect 165154 57922 165250 57978
rect 165306 57922 165374 57978
rect 165430 57922 165498 57978
rect 165554 57922 165622 57978
rect 165678 57922 165774 57978
rect 165154 40350 165774 57922
rect 165154 40294 165250 40350
rect 165306 40294 165374 40350
rect 165430 40294 165498 40350
rect 165554 40294 165622 40350
rect 165678 40294 165774 40350
rect 165154 40226 165774 40294
rect 165154 40170 165250 40226
rect 165306 40170 165374 40226
rect 165430 40170 165498 40226
rect 165554 40170 165622 40226
rect 165678 40170 165774 40226
rect 165154 40102 165774 40170
rect 165154 40046 165250 40102
rect 165306 40046 165374 40102
rect 165430 40046 165498 40102
rect 165554 40046 165622 40102
rect 165678 40046 165774 40102
rect 165154 39978 165774 40046
rect 165154 39922 165250 39978
rect 165306 39922 165374 39978
rect 165430 39922 165498 39978
rect 165554 39922 165622 39978
rect 165678 39922 165774 39978
rect 165154 22350 165774 39922
rect 165154 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 165774 22350
rect 165154 22226 165774 22294
rect 165154 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 165774 22226
rect 165154 22102 165774 22170
rect 165154 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 165774 22102
rect 165154 21978 165774 22046
rect 165154 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 165774 21978
rect 165154 4350 165774 21922
rect 165154 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 165774 4350
rect 165154 4226 165774 4294
rect 165154 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 165774 4226
rect 165154 4102 165774 4170
rect 165154 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 165774 4102
rect 165154 3978 165774 4046
rect 165154 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 165774 3978
rect 165154 -160 165774 3922
rect 165154 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 165774 -160
rect 165154 -284 165774 -216
rect 165154 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 165774 -284
rect 165154 -408 165774 -340
rect 165154 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 165774 -408
rect 165154 -532 165774 -464
rect 165154 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 165774 -532
rect 165154 -1644 165774 -588
rect 168874 598172 169494 598268
rect 168874 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 169494 598172
rect 168874 598048 169494 598116
rect 168874 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 169494 598048
rect 168874 597924 169494 597992
rect 168874 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 169494 597924
rect 168874 597800 169494 597868
rect 168874 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 169494 597800
rect 168874 586350 169494 597744
rect 168874 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 169494 586350
rect 168874 586226 169494 586294
rect 168874 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 169494 586226
rect 168874 586102 169494 586170
rect 168874 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 169494 586102
rect 168874 585978 169494 586046
rect 168874 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 169494 585978
rect 168874 568350 169494 585922
rect 168874 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 169494 568350
rect 168874 568226 169494 568294
rect 168874 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 169494 568226
rect 168874 568102 169494 568170
rect 168874 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 169494 568102
rect 168874 567978 169494 568046
rect 168874 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 169494 567978
rect 168874 550350 169494 567922
rect 168874 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 169494 550350
rect 168874 550226 169494 550294
rect 168874 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 169494 550226
rect 168874 550102 169494 550170
rect 168874 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 169494 550102
rect 168874 549978 169494 550046
rect 168874 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 169494 549978
rect 168874 532350 169494 549922
rect 168874 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 169494 532350
rect 168874 532226 169494 532294
rect 168874 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 169494 532226
rect 168874 532102 169494 532170
rect 168874 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 169494 532102
rect 168874 531978 169494 532046
rect 168874 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 169494 531978
rect 168874 514350 169494 531922
rect 168874 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 169494 514350
rect 168874 514226 169494 514294
rect 168874 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 169494 514226
rect 168874 514102 169494 514170
rect 168874 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 169494 514102
rect 168874 513978 169494 514046
rect 168874 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 169494 513978
rect 168874 496350 169494 513922
rect 168874 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 169494 496350
rect 168874 496226 169494 496294
rect 168874 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 169494 496226
rect 168874 496102 169494 496170
rect 168874 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 169494 496102
rect 168874 495978 169494 496046
rect 168874 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 169494 495978
rect 168874 478350 169494 495922
rect 168874 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 169494 478350
rect 168874 478226 169494 478294
rect 168874 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 169494 478226
rect 168874 478102 169494 478170
rect 168874 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 169494 478102
rect 168874 477978 169494 478046
rect 168874 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 169494 477978
rect 168874 460350 169494 477922
rect 168874 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 169494 460350
rect 168874 460226 169494 460294
rect 168874 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 169494 460226
rect 168874 460102 169494 460170
rect 168874 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 169494 460102
rect 168874 459978 169494 460046
rect 168874 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 169494 459978
rect 168874 442350 169494 459922
rect 168874 442294 168970 442350
rect 169026 442294 169094 442350
rect 169150 442294 169218 442350
rect 169274 442294 169342 442350
rect 169398 442294 169494 442350
rect 168874 442226 169494 442294
rect 168874 442170 168970 442226
rect 169026 442170 169094 442226
rect 169150 442170 169218 442226
rect 169274 442170 169342 442226
rect 169398 442170 169494 442226
rect 168874 442102 169494 442170
rect 168874 442046 168970 442102
rect 169026 442046 169094 442102
rect 169150 442046 169218 442102
rect 169274 442046 169342 442102
rect 169398 442046 169494 442102
rect 168874 441978 169494 442046
rect 168874 441922 168970 441978
rect 169026 441922 169094 441978
rect 169150 441922 169218 441978
rect 169274 441922 169342 441978
rect 169398 441922 169494 441978
rect 168874 424350 169494 441922
rect 168874 424294 168970 424350
rect 169026 424294 169094 424350
rect 169150 424294 169218 424350
rect 169274 424294 169342 424350
rect 169398 424294 169494 424350
rect 168874 424226 169494 424294
rect 168874 424170 168970 424226
rect 169026 424170 169094 424226
rect 169150 424170 169218 424226
rect 169274 424170 169342 424226
rect 169398 424170 169494 424226
rect 168874 424102 169494 424170
rect 168874 424046 168970 424102
rect 169026 424046 169094 424102
rect 169150 424046 169218 424102
rect 169274 424046 169342 424102
rect 169398 424046 169494 424102
rect 168874 423978 169494 424046
rect 168874 423922 168970 423978
rect 169026 423922 169094 423978
rect 169150 423922 169218 423978
rect 169274 423922 169342 423978
rect 169398 423922 169494 423978
rect 168874 406350 169494 423922
rect 168874 406294 168970 406350
rect 169026 406294 169094 406350
rect 169150 406294 169218 406350
rect 169274 406294 169342 406350
rect 169398 406294 169494 406350
rect 168874 406226 169494 406294
rect 168874 406170 168970 406226
rect 169026 406170 169094 406226
rect 169150 406170 169218 406226
rect 169274 406170 169342 406226
rect 169398 406170 169494 406226
rect 168874 406102 169494 406170
rect 168874 406046 168970 406102
rect 169026 406046 169094 406102
rect 169150 406046 169218 406102
rect 169274 406046 169342 406102
rect 169398 406046 169494 406102
rect 168874 405978 169494 406046
rect 168874 405922 168970 405978
rect 169026 405922 169094 405978
rect 169150 405922 169218 405978
rect 169274 405922 169342 405978
rect 169398 405922 169494 405978
rect 168874 388350 169494 405922
rect 168874 388294 168970 388350
rect 169026 388294 169094 388350
rect 169150 388294 169218 388350
rect 169274 388294 169342 388350
rect 169398 388294 169494 388350
rect 168874 388226 169494 388294
rect 168874 388170 168970 388226
rect 169026 388170 169094 388226
rect 169150 388170 169218 388226
rect 169274 388170 169342 388226
rect 169398 388170 169494 388226
rect 168874 388102 169494 388170
rect 168874 388046 168970 388102
rect 169026 388046 169094 388102
rect 169150 388046 169218 388102
rect 169274 388046 169342 388102
rect 169398 388046 169494 388102
rect 168874 387978 169494 388046
rect 168874 387922 168970 387978
rect 169026 387922 169094 387978
rect 169150 387922 169218 387978
rect 169274 387922 169342 387978
rect 169398 387922 169494 387978
rect 168874 370350 169494 387922
rect 168874 370294 168970 370350
rect 169026 370294 169094 370350
rect 169150 370294 169218 370350
rect 169274 370294 169342 370350
rect 169398 370294 169494 370350
rect 168874 370226 169494 370294
rect 168874 370170 168970 370226
rect 169026 370170 169094 370226
rect 169150 370170 169218 370226
rect 169274 370170 169342 370226
rect 169398 370170 169494 370226
rect 168874 370102 169494 370170
rect 168874 370046 168970 370102
rect 169026 370046 169094 370102
rect 169150 370046 169218 370102
rect 169274 370046 169342 370102
rect 169398 370046 169494 370102
rect 168874 369978 169494 370046
rect 168874 369922 168970 369978
rect 169026 369922 169094 369978
rect 169150 369922 169218 369978
rect 169274 369922 169342 369978
rect 169398 369922 169494 369978
rect 168874 352350 169494 369922
rect 168874 352294 168970 352350
rect 169026 352294 169094 352350
rect 169150 352294 169218 352350
rect 169274 352294 169342 352350
rect 169398 352294 169494 352350
rect 168874 352226 169494 352294
rect 168874 352170 168970 352226
rect 169026 352170 169094 352226
rect 169150 352170 169218 352226
rect 169274 352170 169342 352226
rect 169398 352170 169494 352226
rect 168874 352102 169494 352170
rect 168874 352046 168970 352102
rect 169026 352046 169094 352102
rect 169150 352046 169218 352102
rect 169274 352046 169342 352102
rect 169398 352046 169494 352102
rect 168874 351978 169494 352046
rect 168874 351922 168970 351978
rect 169026 351922 169094 351978
rect 169150 351922 169218 351978
rect 169274 351922 169342 351978
rect 169398 351922 169494 351978
rect 168874 334350 169494 351922
rect 168874 334294 168970 334350
rect 169026 334294 169094 334350
rect 169150 334294 169218 334350
rect 169274 334294 169342 334350
rect 169398 334294 169494 334350
rect 168874 334226 169494 334294
rect 168874 334170 168970 334226
rect 169026 334170 169094 334226
rect 169150 334170 169218 334226
rect 169274 334170 169342 334226
rect 169398 334170 169494 334226
rect 168874 334102 169494 334170
rect 168874 334046 168970 334102
rect 169026 334046 169094 334102
rect 169150 334046 169218 334102
rect 169274 334046 169342 334102
rect 169398 334046 169494 334102
rect 168874 333978 169494 334046
rect 168874 333922 168970 333978
rect 169026 333922 169094 333978
rect 169150 333922 169218 333978
rect 169274 333922 169342 333978
rect 169398 333922 169494 333978
rect 168874 316350 169494 333922
rect 168874 316294 168970 316350
rect 169026 316294 169094 316350
rect 169150 316294 169218 316350
rect 169274 316294 169342 316350
rect 169398 316294 169494 316350
rect 168874 316226 169494 316294
rect 168874 316170 168970 316226
rect 169026 316170 169094 316226
rect 169150 316170 169218 316226
rect 169274 316170 169342 316226
rect 169398 316170 169494 316226
rect 168874 316102 169494 316170
rect 168874 316046 168970 316102
rect 169026 316046 169094 316102
rect 169150 316046 169218 316102
rect 169274 316046 169342 316102
rect 169398 316046 169494 316102
rect 168874 315978 169494 316046
rect 168874 315922 168970 315978
rect 169026 315922 169094 315978
rect 169150 315922 169218 315978
rect 169274 315922 169342 315978
rect 169398 315922 169494 315978
rect 168874 298350 169494 315922
rect 168874 298294 168970 298350
rect 169026 298294 169094 298350
rect 169150 298294 169218 298350
rect 169274 298294 169342 298350
rect 169398 298294 169494 298350
rect 168874 298226 169494 298294
rect 168874 298170 168970 298226
rect 169026 298170 169094 298226
rect 169150 298170 169218 298226
rect 169274 298170 169342 298226
rect 169398 298170 169494 298226
rect 168874 298102 169494 298170
rect 168874 298046 168970 298102
rect 169026 298046 169094 298102
rect 169150 298046 169218 298102
rect 169274 298046 169342 298102
rect 169398 298046 169494 298102
rect 168874 297978 169494 298046
rect 168874 297922 168970 297978
rect 169026 297922 169094 297978
rect 169150 297922 169218 297978
rect 169274 297922 169342 297978
rect 169398 297922 169494 297978
rect 168874 280350 169494 297922
rect 168874 280294 168970 280350
rect 169026 280294 169094 280350
rect 169150 280294 169218 280350
rect 169274 280294 169342 280350
rect 169398 280294 169494 280350
rect 168874 280226 169494 280294
rect 168874 280170 168970 280226
rect 169026 280170 169094 280226
rect 169150 280170 169218 280226
rect 169274 280170 169342 280226
rect 169398 280170 169494 280226
rect 168874 280102 169494 280170
rect 168874 280046 168970 280102
rect 169026 280046 169094 280102
rect 169150 280046 169218 280102
rect 169274 280046 169342 280102
rect 169398 280046 169494 280102
rect 168874 279978 169494 280046
rect 168874 279922 168970 279978
rect 169026 279922 169094 279978
rect 169150 279922 169218 279978
rect 169274 279922 169342 279978
rect 169398 279922 169494 279978
rect 168874 262350 169494 279922
rect 168874 262294 168970 262350
rect 169026 262294 169094 262350
rect 169150 262294 169218 262350
rect 169274 262294 169342 262350
rect 169398 262294 169494 262350
rect 168874 262226 169494 262294
rect 168874 262170 168970 262226
rect 169026 262170 169094 262226
rect 169150 262170 169218 262226
rect 169274 262170 169342 262226
rect 169398 262170 169494 262226
rect 168874 262102 169494 262170
rect 168874 262046 168970 262102
rect 169026 262046 169094 262102
rect 169150 262046 169218 262102
rect 169274 262046 169342 262102
rect 169398 262046 169494 262102
rect 168874 261978 169494 262046
rect 168874 261922 168970 261978
rect 169026 261922 169094 261978
rect 169150 261922 169218 261978
rect 169274 261922 169342 261978
rect 169398 261922 169494 261978
rect 168874 244350 169494 261922
rect 168874 244294 168970 244350
rect 169026 244294 169094 244350
rect 169150 244294 169218 244350
rect 169274 244294 169342 244350
rect 169398 244294 169494 244350
rect 168874 244226 169494 244294
rect 168874 244170 168970 244226
rect 169026 244170 169094 244226
rect 169150 244170 169218 244226
rect 169274 244170 169342 244226
rect 169398 244170 169494 244226
rect 168874 244102 169494 244170
rect 168874 244046 168970 244102
rect 169026 244046 169094 244102
rect 169150 244046 169218 244102
rect 169274 244046 169342 244102
rect 169398 244046 169494 244102
rect 168874 243978 169494 244046
rect 168874 243922 168970 243978
rect 169026 243922 169094 243978
rect 169150 243922 169218 243978
rect 169274 243922 169342 243978
rect 169398 243922 169494 243978
rect 168874 226350 169494 243922
rect 168874 226294 168970 226350
rect 169026 226294 169094 226350
rect 169150 226294 169218 226350
rect 169274 226294 169342 226350
rect 169398 226294 169494 226350
rect 168874 226226 169494 226294
rect 168874 226170 168970 226226
rect 169026 226170 169094 226226
rect 169150 226170 169218 226226
rect 169274 226170 169342 226226
rect 169398 226170 169494 226226
rect 168874 226102 169494 226170
rect 168874 226046 168970 226102
rect 169026 226046 169094 226102
rect 169150 226046 169218 226102
rect 169274 226046 169342 226102
rect 169398 226046 169494 226102
rect 168874 225978 169494 226046
rect 168874 225922 168970 225978
rect 169026 225922 169094 225978
rect 169150 225922 169218 225978
rect 169274 225922 169342 225978
rect 169398 225922 169494 225978
rect 168874 208350 169494 225922
rect 168874 208294 168970 208350
rect 169026 208294 169094 208350
rect 169150 208294 169218 208350
rect 169274 208294 169342 208350
rect 169398 208294 169494 208350
rect 168874 208226 169494 208294
rect 168874 208170 168970 208226
rect 169026 208170 169094 208226
rect 169150 208170 169218 208226
rect 169274 208170 169342 208226
rect 169398 208170 169494 208226
rect 168874 208102 169494 208170
rect 168874 208046 168970 208102
rect 169026 208046 169094 208102
rect 169150 208046 169218 208102
rect 169274 208046 169342 208102
rect 169398 208046 169494 208102
rect 168874 207978 169494 208046
rect 168874 207922 168970 207978
rect 169026 207922 169094 207978
rect 169150 207922 169218 207978
rect 169274 207922 169342 207978
rect 169398 207922 169494 207978
rect 168874 190350 169494 207922
rect 168874 190294 168970 190350
rect 169026 190294 169094 190350
rect 169150 190294 169218 190350
rect 169274 190294 169342 190350
rect 169398 190294 169494 190350
rect 168874 190226 169494 190294
rect 168874 190170 168970 190226
rect 169026 190170 169094 190226
rect 169150 190170 169218 190226
rect 169274 190170 169342 190226
rect 169398 190170 169494 190226
rect 168874 190102 169494 190170
rect 168874 190046 168970 190102
rect 169026 190046 169094 190102
rect 169150 190046 169218 190102
rect 169274 190046 169342 190102
rect 169398 190046 169494 190102
rect 168874 189978 169494 190046
rect 168874 189922 168970 189978
rect 169026 189922 169094 189978
rect 169150 189922 169218 189978
rect 169274 189922 169342 189978
rect 169398 189922 169494 189978
rect 168874 172350 169494 189922
rect 168874 172294 168970 172350
rect 169026 172294 169094 172350
rect 169150 172294 169218 172350
rect 169274 172294 169342 172350
rect 169398 172294 169494 172350
rect 168874 172226 169494 172294
rect 168874 172170 168970 172226
rect 169026 172170 169094 172226
rect 169150 172170 169218 172226
rect 169274 172170 169342 172226
rect 169398 172170 169494 172226
rect 168874 172102 169494 172170
rect 168874 172046 168970 172102
rect 169026 172046 169094 172102
rect 169150 172046 169218 172102
rect 169274 172046 169342 172102
rect 169398 172046 169494 172102
rect 168874 171978 169494 172046
rect 168874 171922 168970 171978
rect 169026 171922 169094 171978
rect 169150 171922 169218 171978
rect 169274 171922 169342 171978
rect 169398 171922 169494 171978
rect 168874 154350 169494 171922
rect 168874 154294 168970 154350
rect 169026 154294 169094 154350
rect 169150 154294 169218 154350
rect 169274 154294 169342 154350
rect 169398 154294 169494 154350
rect 168874 154226 169494 154294
rect 168874 154170 168970 154226
rect 169026 154170 169094 154226
rect 169150 154170 169218 154226
rect 169274 154170 169342 154226
rect 169398 154170 169494 154226
rect 168874 154102 169494 154170
rect 168874 154046 168970 154102
rect 169026 154046 169094 154102
rect 169150 154046 169218 154102
rect 169274 154046 169342 154102
rect 169398 154046 169494 154102
rect 168874 153978 169494 154046
rect 168874 153922 168970 153978
rect 169026 153922 169094 153978
rect 169150 153922 169218 153978
rect 169274 153922 169342 153978
rect 169398 153922 169494 153978
rect 168874 136350 169494 153922
rect 168874 136294 168970 136350
rect 169026 136294 169094 136350
rect 169150 136294 169218 136350
rect 169274 136294 169342 136350
rect 169398 136294 169494 136350
rect 168874 136226 169494 136294
rect 168874 136170 168970 136226
rect 169026 136170 169094 136226
rect 169150 136170 169218 136226
rect 169274 136170 169342 136226
rect 169398 136170 169494 136226
rect 168874 136102 169494 136170
rect 168874 136046 168970 136102
rect 169026 136046 169094 136102
rect 169150 136046 169218 136102
rect 169274 136046 169342 136102
rect 169398 136046 169494 136102
rect 168874 135978 169494 136046
rect 168874 135922 168970 135978
rect 169026 135922 169094 135978
rect 169150 135922 169218 135978
rect 169274 135922 169342 135978
rect 169398 135922 169494 135978
rect 168874 118350 169494 135922
rect 168874 118294 168970 118350
rect 169026 118294 169094 118350
rect 169150 118294 169218 118350
rect 169274 118294 169342 118350
rect 169398 118294 169494 118350
rect 168874 118226 169494 118294
rect 168874 118170 168970 118226
rect 169026 118170 169094 118226
rect 169150 118170 169218 118226
rect 169274 118170 169342 118226
rect 169398 118170 169494 118226
rect 168874 118102 169494 118170
rect 168874 118046 168970 118102
rect 169026 118046 169094 118102
rect 169150 118046 169218 118102
rect 169274 118046 169342 118102
rect 169398 118046 169494 118102
rect 168874 117978 169494 118046
rect 168874 117922 168970 117978
rect 169026 117922 169094 117978
rect 169150 117922 169218 117978
rect 169274 117922 169342 117978
rect 169398 117922 169494 117978
rect 168874 100350 169494 117922
rect 168874 100294 168970 100350
rect 169026 100294 169094 100350
rect 169150 100294 169218 100350
rect 169274 100294 169342 100350
rect 169398 100294 169494 100350
rect 168874 100226 169494 100294
rect 168874 100170 168970 100226
rect 169026 100170 169094 100226
rect 169150 100170 169218 100226
rect 169274 100170 169342 100226
rect 169398 100170 169494 100226
rect 168874 100102 169494 100170
rect 168874 100046 168970 100102
rect 169026 100046 169094 100102
rect 169150 100046 169218 100102
rect 169274 100046 169342 100102
rect 169398 100046 169494 100102
rect 168874 99978 169494 100046
rect 168874 99922 168970 99978
rect 169026 99922 169094 99978
rect 169150 99922 169218 99978
rect 169274 99922 169342 99978
rect 169398 99922 169494 99978
rect 168874 82350 169494 99922
rect 168874 82294 168970 82350
rect 169026 82294 169094 82350
rect 169150 82294 169218 82350
rect 169274 82294 169342 82350
rect 169398 82294 169494 82350
rect 168874 82226 169494 82294
rect 168874 82170 168970 82226
rect 169026 82170 169094 82226
rect 169150 82170 169218 82226
rect 169274 82170 169342 82226
rect 169398 82170 169494 82226
rect 168874 82102 169494 82170
rect 168874 82046 168970 82102
rect 169026 82046 169094 82102
rect 169150 82046 169218 82102
rect 169274 82046 169342 82102
rect 169398 82046 169494 82102
rect 168874 81978 169494 82046
rect 168874 81922 168970 81978
rect 169026 81922 169094 81978
rect 169150 81922 169218 81978
rect 169274 81922 169342 81978
rect 169398 81922 169494 81978
rect 168874 64350 169494 81922
rect 168874 64294 168970 64350
rect 169026 64294 169094 64350
rect 169150 64294 169218 64350
rect 169274 64294 169342 64350
rect 169398 64294 169494 64350
rect 168874 64226 169494 64294
rect 168874 64170 168970 64226
rect 169026 64170 169094 64226
rect 169150 64170 169218 64226
rect 169274 64170 169342 64226
rect 169398 64170 169494 64226
rect 168874 64102 169494 64170
rect 168874 64046 168970 64102
rect 169026 64046 169094 64102
rect 169150 64046 169218 64102
rect 169274 64046 169342 64102
rect 169398 64046 169494 64102
rect 168874 63978 169494 64046
rect 168874 63922 168970 63978
rect 169026 63922 169094 63978
rect 169150 63922 169218 63978
rect 169274 63922 169342 63978
rect 169398 63922 169494 63978
rect 168874 46350 169494 63922
rect 168874 46294 168970 46350
rect 169026 46294 169094 46350
rect 169150 46294 169218 46350
rect 169274 46294 169342 46350
rect 169398 46294 169494 46350
rect 168874 46226 169494 46294
rect 168874 46170 168970 46226
rect 169026 46170 169094 46226
rect 169150 46170 169218 46226
rect 169274 46170 169342 46226
rect 169398 46170 169494 46226
rect 168874 46102 169494 46170
rect 168874 46046 168970 46102
rect 169026 46046 169094 46102
rect 169150 46046 169218 46102
rect 169274 46046 169342 46102
rect 169398 46046 169494 46102
rect 168874 45978 169494 46046
rect 168874 45922 168970 45978
rect 169026 45922 169094 45978
rect 169150 45922 169218 45978
rect 169274 45922 169342 45978
rect 169398 45922 169494 45978
rect 168874 28350 169494 45922
rect 168874 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 169494 28350
rect 168874 28226 169494 28294
rect 168874 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 169494 28226
rect 168874 28102 169494 28170
rect 168874 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 169494 28102
rect 168874 27978 169494 28046
rect 168874 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 169494 27978
rect 168874 10350 169494 27922
rect 168874 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 169494 10350
rect 168874 10226 169494 10294
rect 168874 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 169494 10226
rect 168874 10102 169494 10170
rect 168874 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 169494 10102
rect 168874 9978 169494 10046
rect 168874 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 169494 9978
rect 168874 -1120 169494 9922
rect 168874 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 169494 -1120
rect 168874 -1244 169494 -1176
rect 168874 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 169494 -1244
rect 168874 -1368 169494 -1300
rect 168874 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 169494 -1368
rect 168874 -1492 169494 -1424
rect 168874 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 169494 -1492
rect 168874 -1644 169494 -1548
rect 183154 597212 183774 598268
rect 183154 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 183774 597212
rect 183154 597088 183774 597156
rect 183154 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 183774 597088
rect 183154 596964 183774 597032
rect 183154 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 183774 596964
rect 183154 596840 183774 596908
rect 183154 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 183774 596840
rect 183154 580350 183774 596784
rect 183154 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 183774 580350
rect 183154 580226 183774 580294
rect 183154 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 183774 580226
rect 183154 580102 183774 580170
rect 183154 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 183774 580102
rect 183154 579978 183774 580046
rect 183154 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 183774 579978
rect 183154 562350 183774 579922
rect 183154 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 183774 562350
rect 183154 562226 183774 562294
rect 183154 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 183774 562226
rect 183154 562102 183774 562170
rect 183154 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 183774 562102
rect 183154 561978 183774 562046
rect 183154 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 183774 561978
rect 183154 544350 183774 561922
rect 183154 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 183774 544350
rect 183154 544226 183774 544294
rect 183154 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 183774 544226
rect 183154 544102 183774 544170
rect 183154 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 183774 544102
rect 183154 543978 183774 544046
rect 183154 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 183774 543978
rect 183154 526350 183774 543922
rect 183154 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 183774 526350
rect 183154 526226 183774 526294
rect 183154 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 183774 526226
rect 183154 526102 183774 526170
rect 183154 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 183774 526102
rect 183154 525978 183774 526046
rect 183154 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 183774 525978
rect 183154 508350 183774 525922
rect 183154 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 183774 508350
rect 183154 508226 183774 508294
rect 183154 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 183774 508226
rect 183154 508102 183774 508170
rect 183154 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 183774 508102
rect 183154 507978 183774 508046
rect 183154 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 183774 507978
rect 183154 490350 183774 507922
rect 183154 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 183774 490350
rect 183154 490226 183774 490294
rect 183154 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 183774 490226
rect 183154 490102 183774 490170
rect 183154 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 183774 490102
rect 183154 489978 183774 490046
rect 183154 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 183774 489978
rect 183154 472350 183774 489922
rect 183154 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 183774 472350
rect 183154 472226 183774 472294
rect 183154 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 183774 472226
rect 183154 472102 183774 472170
rect 183154 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 183774 472102
rect 183154 471978 183774 472046
rect 183154 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 183774 471978
rect 183154 454350 183774 471922
rect 183154 454294 183250 454350
rect 183306 454294 183374 454350
rect 183430 454294 183498 454350
rect 183554 454294 183622 454350
rect 183678 454294 183774 454350
rect 183154 454226 183774 454294
rect 183154 454170 183250 454226
rect 183306 454170 183374 454226
rect 183430 454170 183498 454226
rect 183554 454170 183622 454226
rect 183678 454170 183774 454226
rect 183154 454102 183774 454170
rect 183154 454046 183250 454102
rect 183306 454046 183374 454102
rect 183430 454046 183498 454102
rect 183554 454046 183622 454102
rect 183678 454046 183774 454102
rect 183154 453978 183774 454046
rect 183154 453922 183250 453978
rect 183306 453922 183374 453978
rect 183430 453922 183498 453978
rect 183554 453922 183622 453978
rect 183678 453922 183774 453978
rect 183154 436350 183774 453922
rect 183154 436294 183250 436350
rect 183306 436294 183374 436350
rect 183430 436294 183498 436350
rect 183554 436294 183622 436350
rect 183678 436294 183774 436350
rect 183154 436226 183774 436294
rect 183154 436170 183250 436226
rect 183306 436170 183374 436226
rect 183430 436170 183498 436226
rect 183554 436170 183622 436226
rect 183678 436170 183774 436226
rect 183154 436102 183774 436170
rect 183154 436046 183250 436102
rect 183306 436046 183374 436102
rect 183430 436046 183498 436102
rect 183554 436046 183622 436102
rect 183678 436046 183774 436102
rect 183154 435978 183774 436046
rect 183154 435922 183250 435978
rect 183306 435922 183374 435978
rect 183430 435922 183498 435978
rect 183554 435922 183622 435978
rect 183678 435922 183774 435978
rect 183154 418350 183774 435922
rect 183154 418294 183250 418350
rect 183306 418294 183374 418350
rect 183430 418294 183498 418350
rect 183554 418294 183622 418350
rect 183678 418294 183774 418350
rect 183154 418226 183774 418294
rect 183154 418170 183250 418226
rect 183306 418170 183374 418226
rect 183430 418170 183498 418226
rect 183554 418170 183622 418226
rect 183678 418170 183774 418226
rect 183154 418102 183774 418170
rect 183154 418046 183250 418102
rect 183306 418046 183374 418102
rect 183430 418046 183498 418102
rect 183554 418046 183622 418102
rect 183678 418046 183774 418102
rect 183154 417978 183774 418046
rect 183154 417922 183250 417978
rect 183306 417922 183374 417978
rect 183430 417922 183498 417978
rect 183554 417922 183622 417978
rect 183678 417922 183774 417978
rect 183154 400350 183774 417922
rect 183154 400294 183250 400350
rect 183306 400294 183374 400350
rect 183430 400294 183498 400350
rect 183554 400294 183622 400350
rect 183678 400294 183774 400350
rect 183154 400226 183774 400294
rect 183154 400170 183250 400226
rect 183306 400170 183374 400226
rect 183430 400170 183498 400226
rect 183554 400170 183622 400226
rect 183678 400170 183774 400226
rect 183154 400102 183774 400170
rect 183154 400046 183250 400102
rect 183306 400046 183374 400102
rect 183430 400046 183498 400102
rect 183554 400046 183622 400102
rect 183678 400046 183774 400102
rect 183154 399978 183774 400046
rect 183154 399922 183250 399978
rect 183306 399922 183374 399978
rect 183430 399922 183498 399978
rect 183554 399922 183622 399978
rect 183678 399922 183774 399978
rect 183154 382350 183774 399922
rect 183154 382294 183250 382350
rect 183306 382294 183374 382350
rect 183430 382294 183498 382350
rect 183554 382294 183622 382350
rect 183678 382294 183774 382350
rect 183154 382226 183774 382294
rect 183154 382170 183250 382226
rect 183306 382170 183374 382226
rect 183430 382170 183498 382226
rect 183554 382170 183622 382226
rect 183678 382170 183774 382226
rect 183154 382102 183774 382170
rect 183154 382046 183250 382102
rect 183306 382046 183374 382102
rect 183430 382046 183498 382102
rect 183554 382046 183622 382102
rect 183678 382046 183774 382102
rect 183154 381978 183774 382046
rect 183154 381922 183250 381978
rect 183306 381922 183374 381978
rect 183430 381922 183498 381978
rect 183554 381922 183622 381978
rect 183678 381922 183774 381978
rect 183154 364350 183774 381922
rect 183154 364294 183250 364350
rect 183306 364294 183374 364350
rect 183430 364294 183498 364350
rect 183554 364294 183622 364350
rect 183678 364294 183774 364350
rect 183154 364226 183774 364294
rect 183154 364170 183250 364226
rect 183306 364170 183374 364226
rect 183430 364170 183498 364226
rect 183554 364170 183622 364226
rect 183678 364170 183774 364226
rect 183154 364102 183774 364170
rect 183154 364046 183250 364102
rect 183306 364046 183374 364102
rect 183430 364046 183498 364102
rect 183554 364046 183622 364102
rect 183678 364046 183774 364102
rect 183154 363978 183774 364046
rect 183154 363922 183250 363978
rect 183306 363922 183374 363978
rect 183430 363922 183498 363978
rect 183554 363922 183622 363978
rect 183678 363922 183774 363978
rect 183154 346350 183774 363922
rect 183154 346294 183250 346350
rect 183306 346294 183374 346350
rect 183430 346294 183498 346350
rect 183554 346294 183622 346350
rect 183678 346294 183774 346350
rect 183154 346226 183774 346294
rect 183154 346170 183250 346226
rect 183306 346170 183374 346226
rect 183430 346170 183498 346226
rect 183554 346170 183622 346226
rect 183678 346170 183774 346226
rect 183154 346102 183774 346170
rect 183154 346046 183250 346102
rect 183306 346046 183374 346102
rect 183430 346046 183498 346102
rect 183554 346046 183622 346102
rect 183678 346046 183774 346102
rect 183154 345978 183774 346046
rect 183154 345922 183250 345978
rect 183306 345922 183374 345978
rect 183430 345922 183498 345978
rect 183554 345922 183622 345978
rect 183678 345922 183774 345978
rect 183154 328350 183774 345922
rect 183154 328294 183250 328350
rect 183306 328294 183374 328350
rect 183430 328294 183498 328350
rect 183554 328294 183622 328350
rect 183678 328294 183774 328350
rect 183154 328226 183774 328294
rect 183154 328170 183250 328226
rect 183306 328170 183374 328226
rect 183430 328170 183498 328226
rect 183554 328170 183622 328226
rect 183678 328170 183774 328226
rect 183154 328102 183774 328170
rect 183154 328046 183250 328102
rect 183306 328046 183374 328102
rect 183430 328046 183498 328102
rect 183554 328046 183622 328102
rect 183678 328046 183774 328102
rect 183154 327978 183774 328046
rect 183154 327922 183250 327978
rect 183306 327922 183374 327978
rect 183430 327922 183498 327978
rect 183554 327922 183622 327978
rect 183678 327922 183774 327978
rect 183154 310350 183774 327922
rect 183154 310294 183250 310350
rect 183306 310294 183374 310350
rect 183430 310294 183498 310350
rect 183554 310294 183622 310350
rect 183678 310294 183774 310350
rect 183154 310226 183774 310294
rect 183154 310170 183250 310226
rect 183306 310170 183374 310226
rect 183430 310170 183498 310226
rect 183554 310170 183622 310226
rect 183678 310170 183774 310226
rect 183154 310102 183774 310170
rect 183154 310046 183250 310102
rect 183306 310046 183374 310102
rect 183430 310046 183498 310102
rect 183554 310046 183622 310102
rect 183678 310046 183774 310102
rect 183154 309978 183774 310046
rect 183154 309922 183250 309978
rect 183306 309922 183374 309978
rect 183430 309922 183498 309978
rect 183554 309922 183622 309978
rect 183678 309922 183774 309978
rect 183154 292350 183774 309922
rect 183154 292294 183250 292350
rect 183306 292294 183374 292350
rect 183430 292294 183498 292350
rect 183554 292294 183622 292350
rect 183678 292294 183774 292350
rect 183154 292226 183774 292294
rect 183154 292170 183250 292226
rect 183306 292170 183374 292226
rect 183430 292170 183498 292226
rect 183554 292170 183622 292226
rect 183678 292170 183774 292226
rect 183154 292102 183774 292170
rect 183154 292046 183250 292102
rect 183306 292046 183374 292102
rect 183430 292046 183498 292102
rect 183554 292046 183622 292102
rect 183678 292046 183774 292102
rect 183154 291978 183774 292046
rect 183154 291922 183250 291978
rect 183306 291922 183374 291978
rect 183430 291922 183498 291978
rect 183554 291922 183622 291978
rect 183678 291922 183774 291978
rect 183154 274350 183774 291922
rect 183154 274294 183250 274350
rect 183306 274294 183374 274350
rect 183430 274294 183498 274350
rect 183554 274294 183622 274350
rect 183678 274294 183774 274350
rect 183154 274226 183774 274294
rect 183154 274170 183250 274226
rect 183306 274170 183374 274226
rect 183430 274170 183498 274226
rect 183554 274170 183622 274226
rect 183678 274170 183774 274226
rect 183154 274102 183774 274170
rect 183154 274046 183250 274102
rect 183306 274046 183374 274102
rect 183430 274046 183498 274102
rect 183554 274046 183622 274102
rect 183678 274046 183774 274102
rect 183154 273978 183774 274046
rect 183154 273922 183250 273978
rect 183306 273922 183374 273978
rect 183430 273922 183498 273978
rect 183554 273922 183622 273978
rect 183678 273922 183774 273978
rect 183154 256350 183774 273922
rect 183154 256294 183250 256350
rect 183306 256294 183374 256350
rect 183430 256294 183498 256350
rect 183554 256294 183622 256350
rect 183678 256294 183774 256350
rect 183154 256226 183774 256294
rect 183154 256170 183250 256226
rect 183306 256170 183374 256226
rect 183430 256170 183498 256226
rect 183554 256170 183622 256226
rect 183678 256170 183774 256226
rect 183154 256102 183774 256170
rect 183154 256046 183250 256102
rect 183306 256046 183374 256102
rect 183430 256046 183498 256102
rect 183554 256046 183622 256102
rect 183678 256046 183774 256102
rect 183154 255978 183774 256046
rect 183154 255922 183250 255978
rect 183306 255922 183374 255978
rect 183430 255922 183498 255978
rect 183554 255922 183622 255978
rect 183678 255922 183774 255978
rect 183154 238350 183774 255922
rect 183154 238294 183250 238350
rect 183306 238294 183374 238350
rect 183430 238294 183498 238350
rect 183554 238294 183622 238350
rect 183678 238294 183774 238350
rect 183154 238226 183774 238294
rect 183154 238170 183250 238226
rect 183306 238170 183374 238226
rect 183430 238170 183498 238226
rect 183554 238170 183622 238226
rect 183678 238170 183774 238226
rect 183154 238102 183774 238170
rect 183154 238046 183250 238102
rect 183306 238046 183374 238102
rect 183430 238046 183498 238102
rect 183554 238046 183622 238102
rect 183678 238046 183774 238102
rect 183154 237978 183774 238046
rect 183154 237922 183250 237978
rect 183306 237922 183374 237978
rect 183430 237922 183498 237978
rect 183554 237922 183622 237978
rect 183678 237922 183774 237978
rect 183154 220350 183774 237922
rect 183154 220294 183250 220350
rect 183306 220294 183374 220350
rect 183430 220294 183498 220350
rect 183554 220294 183622 220350
rect 183678 220294 183774 220350
rect 183154 220226 183774 220294
rect 183154 220170 183250 220226
rect 183306 220170 183374 220226
rect 183430 220170 183498 220226
rect 183554 220170 183622 220226
rect 183678 220170 183774 220226
rect 183154 220102 183774 220170
rect 183154 220046 183250 220102
rect 183306 220046 183374 220102
rect 183430 220046 183498 220102
rect 183554 220046 183622 220102
rect 183678 220046 183774 220102
rect 183154 219978 183774 220046
rect 183154 219922 183250 219978
rect 183306 219922 183374 219978
rect 183430 219922 183498 219978
rect 183554 219922 183622 219978
rect 183678 219922 183774 219978
rect 183154 202350 183774 219922
rect 183154 202294 183250 202350
rect 183306 202294 183374 202350
rect 183430 202294 183498 202350
rect 183554 202294 183622 202350
rect 183678 202294 183774 202350
rect 183154 202226 183774 202294
rect 183154 202170 183250 202226
rect 183306 202170 183374 202226
rect 183430 202170 183498 202226
rect 183554 202170 183622 202226
rect 183678 202170 183774 202226
rect 183154 202102 183774 202170
rect 183154 202046 183250 202102
rect 183306 202046 183374 202102
rect 183430 202046 183498 202102
rect 183554 202046 183622 202102
rect 183678 202046 183774 202102
rect 183154 201978 183774 202046
rect 183154 201922 183250 201978
rect 183306 201922 183374 201978
rect 183430 201922 183498 201978
rect 183554 201922 183622 201978
rect 183678 201922 183774 201978
rect 183154 184350 183774 201922
rect 183154 184294 183250 184350
rect 183306 184294 183374 184350
rect 183430 184294 183498 184350
rect 183554 184294 183622 184350
rect 183678 184294 183774 184350
rect 183154 184226 183774 184294
rect 183154 184170 183250 184226
rect 183306 184170 183374 184226
rect 183430 184170 183498 184226
rect 183554 184170 183622 184226
rect 183678 184170 183774 184226
rect 183154 184102 183774 184170
rect 183154 184046 183250 184102
rect 183306 184046 183374 184102
rect 183430 184046 183498 184102
rect 183554 184046 183622 184102
rect 183678 184046 183774 184102
rect 183154 183978 183774 184046
rect 183154 183922 183250 183978
rect 183306 183922 183374 183978
rect 183430 183922 183498 183978
rect 183554 183922 183622 183978
rect 183678 183922 183774 183978
rect 183154 166350 183774 183922
rect 183154 166294 183250 166350
rect 183306 166294 183374 166350
rect 183430 166294 183498 166350
rect 183554 166294 183622 166350
rect 183678 166294 183774 166350
rect 183154 166226 183774 166294
rect 183154 166170 183250 166226
rect 183306 166170 183374 166226
rect 183430 166170 183498 166226
rect 183554 166170 183622 166226
rect 183678 166170 183774 166226
rect 183154 166102 183774 166170
rect 183154 166046 183250 166102
rect 183306 166046 183374 166102
rect 183430 166046 183498 166102
rect 183554 166046 183622 166102
rect 183678 166046 183774 166102
rect 183154 165978 183774 166046
rect 183154 165922 183250 165978
rect 183306 165922 183374 165978
rect 183430 165922 183498 165978
rect 183554 165922 183622 165978
rect 183678 165922 183774 165978
rect 183154 148350 183774 165922
rect 183154 148294 183250 148350
rect 183306 148294 183374 148350
rect 183430 148294 183498 148350
rect 183554 148294 183622 148350
rect 183678 148294 183774 148350
rect 183154 148226 183774 148294
rect 183154 148170 183250 148226
rect 183306 148170 183374 148226
rect 183430 148170 183498 148226
rect 183554 148170 183622 148226
rect 183678 148170 183774 148226
rect 183154 148102 183774 148170
rect 183154 148046 183250 148102
rect 183306 148046 183374 148102
rect 183430 148046 183498 148102
rect 183554 148046 183622 148102
rect 183678 148046 183774 148102
rect 183154 147978 183774 148046
rect 183154 147922 183250 147978
rect 183306 147922 183374 147978
rect 183430 147922 183498 147978
rect 183554 147922 183622 147978
rect 183678 147922 183774 147978
rect 183154 130350 183774 147922
rect 183154 130294 183250 130350
rect 183306 130294 183374 130350
rect 183430 130294 183498 130350
rect 183554 130294 183622 130350
rect 183678 130294 183774 130350
rect 183154 130226 183774 130294
rect 183154 130170 183250 130226
rect 183306 130170 183374 130226
rect 183430 130170 183498 130226
rect 183554 130170 183622 130226
rect 183678 130170 183774 130226
rect 183154 130102 183774 130170
rect 183154 130046 183250 130102
rect 183306 130046 183374 130102
rect 183430 130046 183498 130102
rect 183554 130046 183622 130102
rect 183678 130046 183774 130102
rect 183154 129978 183774 130046
rect 183154 129922 183250 129978
rect 183306 129922 183374 129978
rect 183430 129922 183498 129978
rect 183554 129922 183622 129978
rect 183678 129922 183774 129978
rect 183154 112350 183774 129922
rect 183154 112294 183250 112350
rect 183306 112294 183374 112350
rect 183430 112294 183498 112350
rect 183554 112294 183622 112350
rect 183678 112294 183774 112350
rect 183154 112226 183774 112294
rect 183154 112170 183250 112226
rect 183306 112170 183374 112226
rect 183430 112170 183498 112226
rect 183554 112170 183622 112226
rect 183678 112170 183774 112226
rect 183154 112102 183774 112170
rect 183154 112046 183250 112102
rect 183306 112046 183374 112102
rect 183430 112046 183498 112102
rect 183554 112046 183622 112102
rect 183678 112046 183774 112102
rect 183154 111978 183774 112046
rect 183154 111922 183250 111978
rect 183306 111922 183374 111978
rect 183430 111922 183498 111978
rect 183554 111922 183622 111978
rect 183678 111922 183774 111978
rect 183154 94350 183774 111922
rect 183154 94294 183250 94350
rect 183306 94294 183374 94350
rect 183430 94294 183498 94350
rect 183554 94294 183622 94350
rect 183678 94294 183774 94350
rect 183154 94226 183774 94294
rect 183154 94170 183250 94226
rect 183306 94170 183374 94226
rect 183430 94170 183498 94226
rect 183554 94170 183622 94226
rect 183678 94170 183774 94226
rect 183154 94102 183774 94170
rect 183154 94046 183250 94102
rect 183306 94046 183374 94102
rect 183430 94046 183498 94102
rect 183554 94046 183622 94102
rect 183678 94046 183774 94102
rect 183154 93978 183774 94046
rect 183154 93922 183250 93978
rect 183306 93922 183374 93978
rect 183430 93922 183498 93978
rect 183554 93922 183622 93978
rect 183678 93922 183774 93978
rect 183154 76350 183774 93922
rect 183154 76294 183250 76350
rect 183306 76294 183374 76350
rect 183430 76294 183498 76350
rect 183554 76294 183622 76350
rect 183678 76294 183774 76350
rect 183154 76226 183774 76294
rect 183154 76170 183250 76226
rect 183306 76170 183374 76226
rect 183430 76170 183498 76226
rect 183554 76170 183622 76226
rect 183678 76170 183774 76226
rect 183154 76102 183774 76170
rect 183154 76046 183250 76102
rect 183306 76046 183374 76102
rect 183430 76046 183498 76102
rect 183554 76046 183622 76102
rect 183678 76046 183774 76102
rect 183154 75978 183774 76046
rect 183154 75922 183250 75978
rect 183306 75922 183374 75978
rect 183430 75922 183498 75978
rect 183554 75922 183622 75978
rect 183678 75922 183774 75978
rect 183154 58350 183774 75922
rect 183154 58294 183250 58350
rect 183306 58294 183374 58350
rect 183430 58294 183498 58350
rect 183554 58294 183622 58350
rect 183678 58294 183774 58350
rect 183154 58226 183774 58294
rect 183154 58170 183250 58226
rect 183306 58170 183374 58226
rect 183430 58170 183498 58226
rect 183554 58170 183622 58226
rect 183678 58170 183774 58226
rect 183154 58102 183774 58170
rect 183154 58046 183250 58102
rect 183306 58046 183374 58102
rect 183430 58046 183498 58102
rect 183554 58046 183622 58102
rect 183678 58046 183774 58102
rect 183154 57978 183774 58046
rect 183154 57922 183250 57978
rect 183306 57922 183374 57978
rect 183430 57922 183498 57978
rect 183554 57922 183622 57978
rect 183678 57922 183774 57978
rect 183154 40350 183774 57922
rect 183154 40294 183250 40350
rect 183306 40294 183374 40350
rect 183430 40294 183498 40350
rect 183554 40294 183622 40350
rect 183678 40294 183774 40350
rect 183154 40226 183774 40294
rect 183154 40170 183250 40226
rect 183306 40170 183374 40226
rect 183430 40170 183498 40226
rect 183554 40170 183622 40226
rect 183678 40170 183774 40226
rect 183154 40102 183774 40170
rect 183154 40046 183250 40102
rect 183306 40046 183374 40102
rect 183430 40046 183498 40102
rect 183554 40046 183622 40102
rect 183678 40046 183774 40102
rect 183154 39978 183774 40046
rect 183154 39922 183250 39978
rect 183306 39922 183374 39978
rect 183430 39922 183498 39978
rect 183554 39922 183622 39978
rect 183678 39922 183774 39978
rect 183154 22350 183774 39922
rect 183154 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 183774 22350
rect 183154 22226 183774 22294
rect 183154 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 183774 22226
rect 183154 22102 183774 22170
rect 183154 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 183774 22102
rect 183154 21978 183774 22046
rect 183154 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 183774 21978
rect 183154 4350 183774 21922
rect 183154 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 183774 4350
rect 183154 4226 183774 4294
rect 183154 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 183774 4226
rect 183154 4102 183774 4170
rect 183154 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 183774 4102
rect 183154 3978 183774 4046
rect 183154 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 183774 3978
rect 183154 -160 183774 3922
rect 183154 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 183774 -160
rect 183154 -284 183774 -216
rect 183154 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 183774 -284
rect 183154 -408 183774 -340
rect 183154 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 183774 -408
rect 183154 -532 183774 -464
rect 183154 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 183774 -532
rect 183154 -1644 183774 -588
rect 186874 598172 187494 598268
rect 186874 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 187494 598172
rect 186874 598048 187494 598116
rect 186874 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 187494 598048
rect 186874 597924 187494 597992
rect 186874 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 187494 597924
rect 186874 597800 187494 597868
rect 186874 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 187494 597800
rect 186874 586350 187494 597744
rect 186874 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 187494 586350
rect 186874 586226 187494 586294
rect 186874 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 187494 586226
rect 186874 586102 187494 586170
rect 186874 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 187494 586102
rect 186874 585978 187494 586046
rect 186874 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 187494 585978
rect 186874 568350 187494 585922
rect 186874 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 187494 568350
rect 186874 568226 187494 568294
rect 186874 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 187494 568226
rect 186874 568102 187494 568170
rect 186874 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 187494 568102
rect 186874 567978 187494 568046
rect 186874 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 187494 567978
rect 186874 550350 187494 567922
rect 186874 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 187494 550350
rect 186874 550226 187494 550294
rect 186874 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 187494 550226
rect 186874 550102 187494 550170
rect 186874 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 187494 550102
rect 186874 549978 187494 550046
rect 186874 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 187494 549978
rect 186874 532350 187494 549922
rect 186874 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 187494 532350
rect 186874 532226 187494 532294
rect 186874 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 187494 532226
rect 186874 532102 187494 532170
rect 186874 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 187494 532102
rect 186874 531978 187494 532046
rect 186874 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 187494 531978
rect 186874 514350 187494 531922
rect 186874 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 187494 514350
rect 186874 514226 187494 514294
rect 186874 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 187494 514226
rect 186874 514102 187494 514170
rect 186874 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 187494 514102
rect 186874 513978 187494 514046
rect 186874 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 187494 513978
rect 186874 496350 187494 513922
rect 186874 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496294 187494 496350
rect 186874 496226 187494 496294
rect 186874 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496170 187494 496226
rect 186874 496102 187494 496170
rect 186874 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496046 187494 496102
rect 186874 495978 187494 496046
rect 186874 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495922 187494 495978
rect 186874 478350 187494 495922
rect 186874 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 187494 478350
rect 186874 478226 187494 478294
rect 186874 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 187494 478226
rect 186874 478102 187494 478170
rect 186874 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 187494 478102
rect 186874 477978 187494 478046
rect 186874 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 187494 477978
rect 186874 460350 187494 477922
rect 186874 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 187494 460350
rect 186874 460226 187494 460294
rect 186874 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 187494 460226
rect 186874 460102 187494 460170
rect 186874 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 187494 460102
rect 186874 459978 187494 460046
rect 186874 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 187494 459978
rect 186874 442350 187494 459922
rect 186874 442294 186970 442350
rect 187026 442294 187094 442350
rect 187150 442294 187218 442350
rect 187274 442294 187342 442350
rect 187398 442294 187494 442350
rect 186874 442226 187494 442294
rect 186874 442170 186970 442226
rect 187026 442170 187094 442226
rect 187150 442170 187218 442226
rect 187274 442170 187342 442226
rect 187398 442170 187494 442226
rect 186874 442102 187494 442170
rect 186874 442046 186970 442102
rect 187026 442046 187094 442102
rect 187150 442046 187218 442102
rect 187274 442046 187342 442102
rect 187398 442046 187494 442102
rect 186874 441978 187494 442046
rect 186874 441922 186970 441978
rect 187026 441922 187094 441978
rect 187150 441922 187218 441978
rect 187274 441922 187342 441978
rect 187398 441922 187494 441978
rect 186874 424350 187494 441922
rect 186874 424294 186970 424350
rect 187026 424294 187094 424350
rect 187150 424294 187218 424350
rect 187274 424294 187342 424350
rect 187398 424294 187494 424350
rect 186874 424226 187494 424294
rect 186874 424170 186970 424226
rect 187026 424170 187094 424226
rect 187150 424170 187218 424226
rect 187274 424170 187342 424226
rect 187398 424170 187494 424226
rect 186874 424102 187494 424170
rect 186874 424046 186970 424102
rect 187026 424046 187094 424102
rect 187150 424046 187218 424102
rect 187274 424046 187342 424102
rect 187398 424046 187494 424102
rect 186874 423978 187494 424046
rect 186874 423922 186970 423978
rect 187026 423922 187094 423978
rect 187150 423922 187218 423978
rect 187274 423922 187342 423978
rect 187398 423922 187494 423978
rect 186874 406350 187494 423922
rect 186874 406294 186970 406350
rect 187026 406294 187094 406350
rect 187150 406294 187218 406350
rect 187274 406294 187342 406350
rect 187398 406294 187494 406350
rect 186874 406226 187494 406294
rect 186874 406170 186970 406226
rect 187026 406170 187094 406226
rect 187150 406170 187218 406226
rect 187274 406170 187342 406226
rect 187398 406170 187494 406226
rect 186874 406102 187494 406170
rect 186874 406046 186970 406102
rect 187026 406046 187094 406102
rect 187150 406046 187218 406102
rect 187274 406046 187342 406102
rect 187398 406046 187494 406102
rect 186874 405978 187494 406046
rect 186874 405922 186970 405978
rect 187026 405922 187094 405978
rect 187150 405922 187218 405978
rect 187274 405922 187342 405978
rect 187398 405922 187494 405978
rect 186874 388350 187494 405922
rect 186874 388294 186970 388350
rect 187026 388294 187094 388350
rect 187150 388294 187218 388350
rect 187274 388294 187342 388350
rect 187398 388294 187494 388350
rect 186874 388226 187494 388294
rect 186874 388170 186970 388226
rect 187026 388170 187094 388226
rect 187150 388170 187218 388226
rect 187274 388170 187342 388226
rect 187398 388170 187494 388226
rect 186874 388102 187494 388170
rect 186874 388046 186970 388102
rect 187026 388046 187094 388102
rect 187150 388046 187218 388102
rect 187274 388046 187342 388102
rect 187398 388046 187494 388102
rect 186874 387978 187494 388046
rect 186874 387922 186970 387978
rect 187026 387922 187094 387978
rect 187150 387922 187218 387978
rect 187274 387922 187342 387978
rect 187398 387922 187494 387978
rect 186874 370350 187494 387922
rect 186874 370294 186970 370350
rect 187026 370294 187094 370350
rect 187150 370294 187218 370350
rect 187274 370294 187342 370350
rect 187398 370294 187494 370350
rect 186874 370226 187494 370294
rect 186874 370170 186970 370226
rect 187026 370170 187094 370226
rect 187150 370170 187218 370226
rect 187274 370170 187342 370226
rect 187398 370170 187494 370226
rect 186874 370102 187494 370170
rect 186874 370046 186970 370102
rect 187026 370046 187094 370102
rect 187150 370046 187218 370102
rect 187274 370046 187342 370102
rect 187398 370046 187494 370102
rect 186874 369978 187494 370046
rect 186874 369922 186970 369978
rect 187026 369922 187094 369978
rect 187150 369922 187218 369978
rect 187274 369922 187342 369978
rect 187398 369922 187494 369978
rect 186874 352350 187494 369922
rect 186874 352294 186970 352350
rect 187026 352294 187094 352350
rect 187150 352294 187218 352350
rect 187274 352294 187342 352350
rect 187398 352294 187494 352350
rect 186874 352226 187494 352294
rect 186874 352170 186970 352226
rect 187026 352170 187094 352226
rect 187150 352170 187218 352226
rect 187274 352170 187342 352226
rect 187398 352170 187494 352226
rect 186874 352102 187494 352170
rect 186874 352046 186970 352102
rect 187026 352046 187094 352102
rect 187150 352046 187218 352102
rect 187274 352046 187342 352102
rect 187398 352046 187494 352102
rect 186874 351978 187494 352046
rect 186874 351922 186970 351978
rect 187026 351922 187094 351978
rect 187150 351922 187218 351978
rect 187274 351922 187342 351978
rect 187398 351922 187494 351978
rect 186874 334350 187494 351922
rect 186874 334294 186970 334350
rect 187026 334294 187094 334350
rect 187150 334294 187218 334350
rect 187274 334294 187342 334350
rect 187398 334294 187494 334350
rect 186874 334226 187494 334294
rect 186874 334170 186970 334226
rect 187026 334170 187094 334226
rect 187150 334170 187218 334226
rect 187274 334170 187342 334226
rect 187398 334170 187494 334226
rect 186874 334102 187494 334170
rect 186874 334046 186970 334102
rect 187026 334046 187094 334102
rect 187150 334046 187218 334102
rect 187274 334046 187342 334102
rect 187398 334046 187494 334102
rect 186874 333978 187494 334046
rect 186874 333922 186970 333978
rect 187026 333922 187094 333978
rect 187150 333922 187218 333978
rect 187274 333922 187342 333978
rect 187398 333922 187494 333978
rect 186874 316350 187494 333922
rect 186874 316294 186970 316350
rect 187026 316294 187094 316350
rect 187150 316294 187218 316350
rect 187274 316294 187342 316350
rect 187398 316294 187494 316350
rect 186874 316226 187494 316294
rect 186874 316170 186970 316226
rect 187026 316170 187094 316226
rect 187150 316170 187218 316226
rect 187274 316170 187342 316226
rect 187398 316170 187494 316226
rect 186874 316102 187494 316170
rect 186874 316046 186970 316102
rect 187026 316046 187094 316102
rect 187150 316046 187218 316102
rect 187274 316046 187342 316102
rect 187398 316046 187494 316102
rect 186874 315978 187494 316046
rect 186874 315922 186970 315978
rect 187026 315922 187094 315978
rect 187150 315922 187218 315978
rect 187274 315922 187342 315978
rect 187398 315922 187494 315978
rect 186874 298350 187494 315922
rect 186874 298294 186970 298350
rect 187026 298294 187094 298350
rect 187150 298294 187218 298350
rect 187274 298294 187342 298350
rect 187398 298294 187494 298350
rect 186874 298226 187494 298294
rect 186874 298170 186970 298226
rect 187026 298170 187094 298226
rect 187150 298170 187218 298226
rect 187274 298170 187342 298226
rect 187398 298170 187494 298226
rect 186874 298102 187494 298170
rect 186874 298046 186970 298102
rect 187026 298046 187094 298102
rect 187150 298046 187218 298102
rect 187274 298046 187342 298102
rect 187398 298046 187494 298102
rect 186874 297978 187494 298046
rect 186874 297922 186970 297978
rect 187026 297922 187094 297978
rect 187150 297922 187218 297978
rect 187274 297922 187342 297978
rect 187398 297922 187494 297978
rect 186874 280350 187494 297922
rect 186874 280294 186970 280350
rect 187026 280294 187094 280350
rect 187150 280294 187218 280350
rect 187274 280294 187342 280350
rect 187398 280294 187494 280350
rect 186874 280226 187494 280294
rect 186874 280170 186970 280226
rect 187026 280170 187094 280226
rect 187150 280170 187218 280226
rect 187274 280170 187342 280226
rect 187398 280170 187494 280226
rect 186874 280102 187494 280170
rect 186874 280046 186970 280102
rect 187026 280046 187094 280102
rect 187150 280046 187218 280102
rect 187274 280046 187342 280102
rect 187398 280046 187494 280102
rect 186874 279978 187494 280046
rect 186874 279922 186970 279978
rect 187026 279922 187094 279978
rect 187150 279922 187218 279978
rect 187274 279922 187342 279978
rect 187398 279922 187494 279978
rect 186874 262350 187494 279922
rect 186874 262294 186970 262350
rect 187026 262294 187094 262350
rect 187150 262294 187218 262350
rect 187274 262294 187342 262350
rect 187398 262294 187494 262350
rect 186874 262226 187494 262294
rect 186874 262170 186970 262226
rect 187026 262170 187094 262226
rect 187150 262170 187218 262226
rect 187274 262170 187342 262226
rect 187398 262170 187494 262226
rect 186874 262102 187494 262170
rect 186874 262046 186970 262102
rect 187026 262046 187094 262102
rect 187150 262046 187218 262102
rect 187274 262046 187342 262102
rect 187398 262046 187494 262102
rect 186874 261978 187494 262046
rect 186874 261922 186970 261978
rect 187026 261922 187094 261978
rect 187150 261922 187218 261978
rect 187274 261922 187342 261978
rect 187398 261922 187494 261978
rect 186874 244350 187494 261922
rect 186874 244294 186970 244350
rect 187026 244294 187094 244350
rect 187150 244294 187218 244350
rect 187274 244294 187342 244350
rect 187398 244294 187494 244350
rect 186874 244226 187494 244294
rect 186874 244170 186970 244226
rect 187026 244170 187094 244226
rect 187150 244170 187218 244226
rect 187274 244170 187342 244226
rect 187398 244170 187494 244226
rect 186874 244102 187494 244170
rect 186874 244046 186970 244102
rect 187026 244046 187094 244102
rect 187150 244046 187218 244102
rect 187274 244046 187342 244102
rect 187398 244046 187494 244102
rect 186874 243978 187494 244046
rect 186874 243922 186970 243978
rect 187026 243922 187094 243978
rect 187150 243922 187218 243978
rect 187274 243922 187342 243978
rect 187398 243922 187494 243978
rect 186874 226350 187494 243922
rect 186874 226294 186970 226350
rect 187026 226294 187094 226350
rect 187150 226294 187218 226350
rect 187274 226294 187342 226350
rect 187398 226294 187494 226350
rect 186874 226226 187494 226294
rect 186874 226170 186970 226226
rect 187026 226170 187094 226226
rect 187150 226170 187218 226226
rect 187274 226170 187342 226226
rect 187398 226170 187494 226226
rect 186874 226102 187494 226170
rect 186874 226046 186970 226102
rect 187026 226046 187094 226102
rect 187150 226046 187218 226102
rect 187274 226046 187342 226102
rect 187398 226046 187494 226102
rect 186874 225978 187494 226046
rect 186874 225922 186970 225978
rect 187026 225922 187094 225978
rect 187150 225922 187218 225978
rect 187274 225922 187342 225978
rect 187398 225922 187494 225978
rect 186874 208350 187494 225922
rect 186874 208294 186970 208350
rect 187026 208294 187094 208350
rect 187150 208294 187218 208350
rect 187274 208294 187342 208350
rect 187398 208294 187494 208350
rect 186874 208226 187494 208294
rect 186874 208170 186970 208226
rect 187026 208170 187094 208226
rect 187150 208170 187218 208226
rect 187274 208170 187342 208226
rect 187398 208170 187494 208226
rect 186874 208102 187494 208170
rect 186874 208046 186970 208102
rect 187026 208046 187094 208102
rect 187150 208046 187218 208102
rect 187274 208046 187342 208102
rect 187398 208046 187494 208102
rect 186874 207978 187494 208046
rect 186874 207922 186970 207978
rect 187026 207922 187094 207978
rect 187150 207922 187218 207978
rect 187274 207922 187342 207978
rect 187398 207922 187494 207978
rect 186874 190350 187494 207922
rect 186874 190294 186970 190350
rect 187026 190294 187094 190350
rect 187150 190294 187218 190350
rect 187274 190294 187342 190350
rect 187398 190294 187494 190350
rect 186874 190226 187494 190294
rect 186874 190170 186970 190226
rect 187026 190170 187094 190226
rect 187150 190170 187218 190226
rect 187274 190170 187342 190226
rect 187398 190170 187494 190226
rect 186874 190102 187494 190170
rect 186874 190046 186970 190102
rect 187026 190046 187094 190102
rect 187150 190046 187218 190102
rect 187274 190046 187342 190102
rect 187398 190046 187494 190102
rect 186874 189978 187494 190046
rect 186874 189922 186970 189978
rect 187026 189922 187094 189978
rect 187150 189922 187218 189978
rect 187274 189922 187342 189978
rect 187398 189922 187494 189978
rect 186874 172350 187494 189922
rect 186874 172294 186970 172350
rect 187026 172294 187094 172350
rect 187150 172294 187218 172350
rect 187274 172294 187342 172350
rect 187398 172294 187494 172350
rect 186874 172226 187494 172294
rect 186874 172170 186970 172226
rect 187026 172170 187094 172226
rect 187150 172170 187218 172226
rect 187274 172170 187342 172226
rect 187398 172170 187494 172226
rect 186874 172102 187494 172170
rect 186874 172046 186970 172102
rect 187026 172046 187094 172102
rect 187150 172046 187218 172102
rect 187274 172046 187342 172102
rect 187398 172046 187494 172102
rect 186874 171978 187494 172046
rect 186874 171922 186970 171978
rect 187026 171922 187094 171978
rect 187150 171922 187218 171978
rect 187274 171922 187342 171978
rect 187398 171922 187494 171978
rect 186874 154350 187494 171922
rect 186874 154294 186970 154350
rect 187026 154294 187094 154350
rect 187150 154294 187218 154350
rect 187274 154294 187342 154350
rect 187398 154294 187494 154350
rect 186874 154226 187494 154294
rect 186874 154170 186970 154226
rect 187026 154170 187094 154226
rect 187150 154170 187218 154226
rect 187274 154170 187342 154226
rect 187398 154170 187494 154226
rect 186874 154102 187494 154170
rect 186874 154046 186970 154102
rect 187026 154046 187094 154102
rect 187150 154046 187218 154102
rect 187274 154046 187342 154102
rect 187398 154046 187494 154102
rect 186874 153978 187494 154046
rect 186874 153922 186970 153978
rect 187026 153922 187094 153978
rect 187150 153922 187218 153978
rect 187274 153922 187342 153978
rect 187398 153922 187494 153978
rect 186874 136350 187494 153922
rect 186874 136294 186970 136350
rect 187026 136294 187094 136350
rect 187150 136294 187218 136350
rect 187274 136294 187342 136350
rect 187398 136294 187494 136350
rect 186874 136226 187494 136294
rect 186874 136170 186970 136226
rect 187026 136170 187094 136226
rect 187150 136170 187218 136226
rect 187274 136170 187342 136226
rect 187398 136170 187494 136226
rect 186874 136102 187494 136170
rect 186874 136046 186970 136102
rect 187026 136046 187094 136102
rect 187150 136046 187218 136102
rect 187274 136046 187342 136102
rect 187398 136046 187494 136102
rect 186874 135978 187494 136046
rect 186874 135922 186970 135978
rect 187026 135922 187094 135978
rect 187150 135922 187218 135978
rect 187274 135922 187342 135978
rect 187398 135922 187494 135978
rect 186874 118350 187494 135922
rect 186874 118294 186970 118350
rect 187026 118294 187094 118350
rect 187150 118294 187218 118350
rect 187274 118294 187342 118350
rect 187398 118294 187494 118350
rect 186874 118226 187494 118294
rect 186874 118170 186970 118226
rect 187026 118170 187094 118226
rect 187150 118170 187218 118226
rect 187274 118170 187342 118226
rect 187398 118170 187494 118226
rect 186874 118102 187494 118170
rect 186874 118046 186970 118102
rect 187026 118046 187094 118102
rect 187150 118046 187218 118102
rect 187274 118046 187342 118102
rect 187398 118046 187494 118102
rect 186874 117978 187494 118046
rect 186874 117922 186970 117978
rect 187026 117922 187094 117978
rect 187150 117922 187218 117978
rect 187274 117922 187342 117978
rect 187398 117922 187494 117978
rect 186874 100350 187494 117922
rect 186874 100294 186970 100350
rect 187026 100294 187094 100350
rect 187150 100294 187218 100350
rect 187274 100294 187342 100350
rect 187398 100294 187494 100350
rect 186874 100226 187494 100294
rect 186874 100170 186970 100226
rect 187026 100170 187094 100226
rect 187150 100170 187218 100226
rect 187274 100170 187342 100226
rect 187398 100170 187494 100226
rect 186874 100102 187494 100170
rect 186874 100046 186970 100102
rect 187026 100046 187094 100102
rect 187150 100046 187218 100102
rect 187274 100046 187342 100102
rect 187398 100046 187494 100102
rect 186874 99978 187494 100046
rect 186874 99922 186970 99978
rect 187026 99922 187094 99978
rect 187150 99922 187218 99978
rect 187274 99922 187342 99978
rect 187398 99922 187494 99978
rect 186874 82350 187494 99922
rect 186874 82294 186970 82350
rect 187026 82294 187094 82350
rect 187150 82294 187218 82350
rect 187274 82294 187342 82350
rect 187398 82294 187494 82350
rect 186874 82226 187494 82294
rect 186874 82170 186970 82226
rect 187026 82170 187094 82226
rect 187150 82170 187218 82226
rect 187274 82170 187342 82226
rect 187398 82170 187494 82226
rect 186874 82102 187494 82170
rect 186874 82046 186970 82102
rect 187026 82046 187094 82102
rect 187150 82046 187218 82102
rect 187274 82046 187342 82102
rect 187398 82046 187494 82102
rect 186874 81978 187494 82046
rect 186874 81922 186970 81978
rect 187026 81922 187094 81978
rect 187150 81922 187218 81978
rect 187274 81922 187342 81978
rect 187398 81922 187494 81978
rect 186874 64350 187494 81922
rect 186874 64294 186970 64350
rect 187026 64294 187094 64350
rect 187150 64294 187218 64350
rect 187274 64294 187342 64350
rect 187398 64294 187494 64350
rect 186874 64226 187494 64294
rect 186874 64170 186970 64226
rect 187026 64170 187094 64226
rect 187150 64170 187218 64226
rect 187274 64170 187342 64226
rect 187398 64170 187494 64226
rect 186874 64102 187494 64170
rect 186874 64046 186970 64102
rect 187026 64046 187094 64102
rect 187150 64046 187218 64102
rect 187274 64046 187342 64102
rect 187398 64046 187494 64102
rect 186874 63978 187494 64046
rect 186874 63922 186970 63978
rect 187026 63922 187094 63978
rect 187150 63922 187218 63978
rect 187274 63922 187342 63978
rect 187398 63922 187494 63978
rect 186874 46350 187494 63922
rect 186874 46294 186970 46350
rect 187026 46294 187094 46350
rect 187150 46294 187218 46350
rect 187274 46294 187342 46350
rect 187398 46294 187494 46350
rect 186874 46226 187494 46294
rect 186874 46170 186970 46226
rect 187026 46170 187094 46226
rect 187150 46170 187218 46226
rect 187274 46170 187342 46226
rect 187398 46170 187494 46226
rect 186874 46102 187494 46170
rect 186874 46046 186970 46102
rect 187026 46046 187094 46102
rect 187150 46046 187218 46102
rect 187274 46046 187342 46102
rect 187398 46046 187494 46102
rect 186874 45978 187494 46046
rect 186874 45922 186970 45978
rect 187026 45922 187094 45978
rect 187150 45922 187218 45978
rect 187274 45922 187342 45978
rect 187398 45922 187494 45978
rect 186874 28350 187494 45922
rect 186874 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 187494 28350
rect 186874 28226 187494 28294
rect 186874 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 187494 28226
rect 186874 28102 187494 28170
rect 186874 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 187494 28102
rect 186874 27978 187494 28046
rect 186874 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 187494 27978
rect 186874 10350 187494 27922
rect 186874 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 187494 10350
rect 186874 10226 187494 10294
rect 186874 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 187494 10226
rect 186874 10102 187494 10170
rect 186874 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 187494 10102
rect 186874 9978 187494 10046
rect 186874 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 187494 9978
rect 186874 -1120 187494 9922
rect 186874 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 187494 -1120
rect 186874 -1244 187494 -1176
rect 186874 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 187494 -1244
rect 186874 -1368 187494 -1300
rect 186874 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 187494 -1368
rect 186874 -1492 187494 -1424
rect 186874 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 187494 -1492
rect 186874 -1644 187494 -1548
rect 201154 597212 201774 598268
rect 201154 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 201774 597212
rect 201154 597088 201774 597156
rect 201154 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 201774 597088
rect 201154 596964 201774 597032
rect 201154 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 201774 596964
rect 201154 596840 201774 596908
rect 201154 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 201774 596840
rect 201154 580350 201774 596784
rect 201154 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 201774 580350
rect 201154 580226 201774 580294
rect 201154 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 201774 580226
rect 201154 580102 201774 580170
rect 201154 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 201774 580102
rect 201154 579978 201774 580046
rect 201154 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 201774 579978
rect 201154 562350 201774 579922
rect 201154 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 201774 562350
rect 201154 562226 201774 562294
rect 201154 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 201774 562226
rect 201154 562102 201774 562170
rect 201154 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 201774 562102
rect 201154 561978 201774 562046
rect 201154 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 201774 561978
rect 201154 544350 201774 561922
rect 201154 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 201774 544350
rect 201154 544226 201774 544294
rect 201154 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 201774 544226
rect 201154 544102 201774 544170
rect 201154 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 201774 544102
rect 201154 543978 201774 544046
rect 201154 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 201774 543978
rect 201154 526350 201774 543922
rect 201154 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 201774 526350
rect 201154 526226 201774 526294
rect 201154 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 201774 526226
rect 201154 526102 201774 526170
rect 201154 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 201774 526102
rect 201154 525978 201774 526046
rect 201154 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 201774 525978
rect 201154 508350 201774 525922
rect 201154 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 201774 508350
rect 201154 508226 201774 508294
rect 201154 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 201774 508226
rect 201154 508102 201774 508170
rect 201154 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 201774 508102
rect 201154 507978 201774 508046
rect 201154 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 201774 507978
rect 201154 490350 201774 507922
rect 204874 598172 205494 598268
rect 204874 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 205494 598172
rect 204874 598048 205494 598116
rect 204874 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 205494 598048
rect 204874 597924 205494 597992
rect 204874 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 205494 597924
rect 204874 597800 205494 597868
rect 204874 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 205494 597800
rect 204874 586350 205494 597744
rect 204874 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 205494 586350
rect 204874 586226 205494 586294
rect 204874 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 205494 586226
rect 204874 586102 205494 586170
rect 204874 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 205494 586102
rect 204874 585978 205494 586046
rect 204874 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 205494 585978
rect 204874 568350 205494 585922
rect 204874 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 205494 568350
rect 204874 568226 205494 568294
rect 204874 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 205494 568226
rect 204874 568102 205494 568170
rect 204874 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 205494 568102
rect 204874 567978 205494 568046
rect 204874 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 205494 567978
rect 204874 550350 205494 567922
rect 204874 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 205494 550350
rect 204874 550226 205494 550294
rect 204874 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 205494 550226
rect 204874 550102 205494 550170
rect 204874 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 205494 550102
rect 204874 549978 205494 550046
rect 204874 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 205494 549978
rect 204874 532350 205494 549922
rect 204874 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 205494 532350
rect 204874 532226 205494 532294
rect 204874 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 205494 532226
rect 204874 532102 205494 532170
rect 204874 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 205494 532102
rect 204874 531978 205494 532046
rect 204874 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 205494 531978
rect 204874 514350 205494 531922
rect 204874 514294 204970 514350
rect 205026 514294 205094 514350
rect 205150 514294 205218 514350
rect 205274 514294 205342 514350
rect 205398 514294 205494 514350
rect 204874 514226 205494 514294
rect 204874 514170 204970 514226
rect 205026 514170 205094 514226
rect 205150 514170 205218 514226
rect 205274 514170 205342 514226
rect 205398 514170 205494 514226
rect 204874 514102 205494 514170
rect 204874 514046 204970 514102
rect 205026 514046 205094 514102
rect 205150 514046 205218 514102
rect 205274 514046 205342 514102
rect 205398 514046 205494 514102
rect 204874 513978 205494 514046
rect 204874 513922 204970 513978
rect 205026 513922 205094 513978
rect 205150 513922 205218 513978
rect 205274 513922 205342 513978
rect 205398 513922 205494 513978
rect 204874 499846 205494 513922
rect 219154 597212 219774 598268
rect 219154 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 219774 597212
rect 219154 597088 219774 597156
rect 219154 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 219774 597088
rect 219154 596964 219774 597032
rect 219154 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 219774 596964
rect 219154 596840 219774 596908
rect 219154 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 219774 596840
rect 219154 580350 219774 596784
rect 219154 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 219774 580350
rect 219154 580226 219774 580294
rect 219154 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 219774 580226
rect 219154 580102 219774 580170
rect 219154 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 219774 580102
rect 219154 579978 219774 580046
rect 219154 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 219774 579978
rect 219154 562350 219774 579922
rect 219154 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 219774 562350
rect 219154 562226 219774 562294
rect 219154 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 219774 562226
rect 219154 562102 219774 562170
rect 219154 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 219774 562102
rect 219154 561978 219774 562046
rect 219154 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 219774 561978
rect 219154 544350 219774 561922
rect 219154 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 219774 544350
rect 219154 544226 219774 544294
rect 219154 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 219774 544226
rect 219154 544102 219774 544170
rect 219154 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 219774 544102
rect 219154 543978 219774 544046
rect 219154 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 219774 543978
rect 219154 526350 219774 543922
rect 219154 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 219774 526350
rect 219154 526226 219774 526294
rect 219154 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 219774 526226
rect 219154 526102 219774 526170
rect 219154 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 219774 526102
rect 219154 525978 219774 526046
rect 219154 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 219774 525978
rect 219154 508350 219774 525922
rect 219154 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 219774 508350
rect 219154 508226 219774 508294
rect 219154 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 219774 508226
rect 219154 508102 219774 508170
rect 219154 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 219774 508102
rect 219154 507978 219774 508046
rect 219154 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 219774 507978
rect 219154 499846 219774 507922
rect 222874 598172 223494 598268
rect 222874 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 223494 598172
rect 222874 598048 223494 598116
rect 222874 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 223494 598048
rect 222874 597924 223494 597992
rect 222874 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 223494 597924
rect 222874 597800 223494 597868
rect 222874 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 223494 597800
rect 222874 586350 223494 597744
rect 222874 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 223494 586350
rect 222874 586226 223494 586294
rect 222874 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 223494 586226
rect 222874 586102 223494 586170
rect 222874 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 223494 586102
rect 222874 585978 223494 586046
rect 222874 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 223494 585978
rect 222874 568350 223494 585922
rect 222874 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 223494 568350
rect 222874 568226 223494 568294
rect 222874 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 223494 568226
rect 222874 568102 223494 568170
rect 222874 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 223494 568102
rect 222874 567978 223494 568046
rect 222874 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 223494 567978
rect 222874 550350 223494 567922
rect 222874 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 223494 550350
rect 222874 550226 223494 550294
rect 222874 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 223494 550226
rect 222874 550102 223494 550170
rect 222874 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 223494 550102
rect 222874 549978 223494 550046
rect 222874 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 223494 549978
rect 222874 532350 223494 549922
rect 222874 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 223494 532350
rect 222874 532226 223494 532294
rect 222874 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 223494 532226
rect 222874 532102 223494 532170
rect 222874 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 223494 532102
rect 222874 531978 223494 532046
rect 222874 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 223494 531978
rect 222874 514350 223494 531922
rect 222874 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 223494 514350
rect 222874 514226 223494 514294
rect 222874 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 223494 514226
rect 222874 514102 223494 514170
rect 222874 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 223494 514102
rect 222874 513978 223494 514046
rect 222874 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 223494 513978
rect 222874 499846 223494 513922
rect 237154 597212 237774 598268
rect 237154 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 237774 597212
rect 237154 597088 237774 597156
rect 237154 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 237774 597088
rect 237154 596964 237774 597032
rect 237154 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 237774 596964
rect 237154 596840 237774 596908
rect 237154 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 237774 596840
rect 237154 580350 237774 596784
rect 237154 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 237774 580350
rect 237154 580226 237774 580294
rect 237154 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 237774 580226
rect 237154 580102 237774 580170
rect 237154 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 237774 580102
rect 237154 579978 237774 580046
rect 237154 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 237774 579978
rect 237154 562350 237774 579922
rect 237154 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 237774 562350
rect 237154 562226 237774 562294
rect 237154 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 237774 562226
rect 237154 562102 237774 562170
rect 237154 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 237774 562102
rect 237154 561978 237774 562046
rect 237154 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 237774 561978
rect 237154 544350 237774 561922
rect 237154 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 237774 544350
rect 237154 544226 237774 544294
rect 237154 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 237774 544226
rect 237154 544102 237774 544170
rect 237154 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 237774 544102
rect 237154 543978 237774 544046
rect 237154 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 237774 543978
rect 237154 526350 237774 543922
rect 237154 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 237774 526350
rect 237154 526226 237774 526294
rect 237154 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 237774 526226
rect 237154 526102 237774 526170
rect 237154 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 237774 526102
rect 237154 525978 237774 526046
rect 237154 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 237774 525978
rect 237154 508350 237774 525922
rect 237154 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 237774 508350
rect 237154 508226 237774 508294
rect 237154 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 237774 508226
rect 237154 508102 237774 508170
rect 237154 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 237774 508102
rect 237154 507978 237774 508046
rect 237154 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 237774 507978
rect 237154 499846 237774 507922
rect 240874 598172 241494 598268
rect 240874 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 241494 598172
rect 240874 598048 241494 598116
rect 240874 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 241494 598048
rect 240874 597924 241494 597992
rect 240874 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 241494 597924
rect 240874 597800 241494 597868
rect 240874 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 241494 597800
rect 240874 586350 241494 597744
rect 240874 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 241494 586350
rect 240874 586226 241494 586294
rect 240874 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 241494 586226
rect 240874 586102 241494 586170
rect 240874 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 241494 586102
rect 240874 585978 241494 586046
rect 240874 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 241494 585978
rect 240874 568350 241494 585922
rect 240874 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 241494 568350
rect 240874 568226 241494 568294
rect 240874 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 241494 568226
rect 240874 568102 241494 568170
rect 240874 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 241494 568102
rect 240874 567978 241494 568046
rect 240874 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 241494 567978
rect 240874 550350 241494 567922
rect 240874 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 241494 550350
rect 240874 550226 241494 550294
rect 240874 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 241494 550226
rect 240874 550102 241494 550170
rect 240874 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 241494 550102
rect 240874 549978 241494 550046
rect 240874 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 241494 549978
rect 240874 532350 241494 549922
rect 240874 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 241494 532350
rect 240874 532226 241494 532294
rect 240874 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 241494 532226
rect 240874 532102 241494 532170
rect 240874 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 241494 532102
rect 240874 531978 241494 532046
rect 240874 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 241494 531978
rect 240874 514350 241494 531922
rect 240874 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 241494 514350
rect 240874 514226 241494 514294
rect 240874 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 241494 514226
rect 240874 514102 241494 514170
rect 240874 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 241494 514102
rect 240874 513978 241494 514046
rect 240874 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 241494 513978
rect 240874 499846 241494 513922
rect 255154 597212 255774 598268
rect 255154 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 255774 597212
rect 255154 597088 255774 597156
rect 255154 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 255774 597088
rect 255154 596964 255774 597032
rect 255154 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 255774 596964
rect 255154 596840 255774 596908
rect 255154 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 255774 596840
rect 255154 580350 255774 596784
rect 255154 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 255774 580350
rect 255154 580226 255774 580294
rect 255154 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 255774 580226
rect 255154 580102 255774 580170
rect 255154 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 255774 580102
rect 255154 579978 255774 580046
rect 255154 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 255774 579978
rect 255154 562350 255774 579922
rect 255154 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 255774 562350
rect 255154 562226 255774 562294
rect 255154 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 255774 562226
rect 255154 562102 255774 562170
rect 255154 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 255774 562102
rect 255154 561978 255774 562046
rect 255154 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 255774 561978
rect 255154 544350 255774 561922
rect 255154 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 255774 544350
rect 255154 544226 255774 544294
rect 255154 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 255774 544226
rect 255154 544102 255774 544170
rect 255154 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 255774 544102
rect 255154 543978 255774 544046
rect 255154 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 255774 543978
rect 255154 526350 255774 543922
rect 255154 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 255774 526350
rect 255154 526226 255774 526294
rect 255154 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 255774 526226
rect 255154 526102 255774 526170
rect 255154 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 255774 526102
rect 255154 525978 255774 526046
rect 255154 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 255774 525978
rect 255154 508350 255774 525922
rect 255154 508294 255250 508350
rect 255306 508294 255374 508350
rect 255430 508294 255498 508350
rect 255554 508294 255622 508350
rect 255678 508294 255774 508350
rect 255154 508226 255774 508294
rect 255154 508170 255250 508226
rect 255306 508170 255374 508226
rect 255430 508170 255498 508226
rect 255554 508170 255622 508226
rect 255678 508170 255774 508226
rect 255154 508102 255774 508170
rect 255154 508046 255250 508102
rect 255306 508046 255374 508102
rect 255430 508046 255498 508102
rect 255554 508046 255622 508102
rect 255678 508046 255774 508102
rect 255154 507978 255774 508046
rect 255154 507922 255250 507978
rect 255306 507922 255374 507978
rect 255430 507922 255498 507978
rect 255554 507922 255622 507978
rect 255678 507922 255774 507978
rect 255154 499846 255774 507922
rect 258874 598172 259494 598268
rect 258874 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 259494 598172
rect 258874 598048 259494 598116
rect 258874 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 259494 598048
rect 258874 597924 259494 597992
rect 258874 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 259494 597924
rect 258874 597800 259494 597868
rect 258874 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 259494 597800
rect 258874 586350 259494 597744
rect 258874 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 259494 586350
rect 258874 586226 259494 586294
rect 258874 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 259494 586226
rect 258874 586102 259494 586170
rect 258874 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 259494 586102
rect 258874 585978 259494 586046
rect 258874 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 259494 585978
rect 258874 568350 259494 585922
rect 258874 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 259494 568350
rect 258874 568226 259494 568294
rect 258874 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 259494 568226
rect 258874 568102 259494 568170
rect 258874 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 259494 568102
rect 258874 567978 259494 568046
rect 258874 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 259494 567978
rect 258874 550350 259494 567922
rect 258874 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 259494 550350
rect 258874 550226 259494 550294
rect 258874 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 259494 550226
rect 258874 550102 259494 550170
rect 258874 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 259494 550102
rect 258874 549978 259494 550046
rect 258874 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 259494 549978
rect 258874 532350 259494 549922
rect 258874 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 259494 532350
rect 258874 532226 259494 532294
rect 258874 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 259494 532226
rect 258874 532102 259494 532170
rect 258874 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 259494 532102
rect 258874 531978 259494 532046
rect 258874 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 259494 531978
rect 258874 514350 259494 531922
rect 258874 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 259494 514350
rect 258874 514226 259494 514294
rect 258874 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 259494 514226
rect 258874 514102 259494 514170
rect 258874 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 259494 514102
rect 258874 513978 259494 514046
rect 258874 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 259494 513978
rect 258874 499846 259494 513922
rect 273154 597212 273774 598268
rect 273154 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 273774 597212
rect 273154 597088 273774 597156
rect 273154 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 273774 597088
rect 273154 596964 273774 597032
rect 273154 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 273774 596964
rect 273154 596840 273774 596908
rect 273154 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 273774 596840
rect 273154 580350 273774 596784
rect 273154 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 273774 580350
rect 273154 580226 273774 580294
rect 273154 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 273774 580226
rect 273154 580102 273774 580170
rect 273154 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 273774 580102
rect 273154 579978 273774 580046
rect 273154 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 273774 579978
rect 273154 562350 273774 579922
rect 273154 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 273774 562350
rect 273154 562226 273774 562294
rect 273154 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 273774 562226
rect 273154 562102 273774 562170
rect 273154 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 273774 562102
rect 273154 561978 273774 562046
rect 273154 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 273774 561978
rect 273154 544350 273774 561922
rect 273154 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 273774 544350
rect 273154 544226 273774 544294
rect 273154 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 273774 544226
rect 273154 544102 273774 544170
rect 273154 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 273774 544102
rect 273154 543978 273774 544046
rect 273154 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 273774 543978
rect 273154 526350 273774 543922
rect 273154 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 273774 526350
rect 273154 526226 273774 526294
rect 273154 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 273774 526226
rect 273154 526102 273774 526170
rect 273154 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 273774 526102
rect 273154 525978 273774 526046
rect 273154 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 273774 525978
rect 273154 508350 273774 525922
rect 273154 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 273774 508350
rect 273154 508226 273774 508294
rect 273154 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 273774 508226
rect 273154 508102 273774 508170
rect 273154 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 273774 508102
rect 273154 507978 273774 508046
rect 273154 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 273774 507978
rect 273154 499846 273774 507922
rect 276874 598172 277494 598268
rect 276874 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 277494 598172
rect 276874 598048 277494 598116
rect 276874 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 277494 598048
rect 276874 597924 277494 597992
rect 276874 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 277494 597924
rect 276874 597800 277494 597868
rect 276874 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 277494 597800
rect 276874 586350 277494 597744
rect 276874 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 277494 586350
rect 276874 586226 277494 586294
rect 276874 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 277494 586226
rect 276874 586102 277494 586170
rect 276874 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 277494 586102
rect 276874 585978 277494 586046
rect 276874 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 277494 585978
rect 276874 568350 277494 585922
rect 276874 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 277494 568350
rect 276874 568226 277494 568294
rect 276874 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 277494 568226
rect 276874 568102 277494 568170
rect 276874 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 277494 568102
rect 276874 567978 277494 568046
rect 276874 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 277494 567978
rect 276874 550350 277494 567922
rect 276874 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 277494 550350
rect 276874 550226 277494 550294
rect 276874 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 277494 550226
rect 276874 550102 277494 550170
rect 276874 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 277494 550102
rect 276874 549978 277494 550046
rect 276874 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 277494 549978
rect 276874 532350 277494 549922
rect 276874 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 277494 532350
rect 276874 532226 277494 532294
rect 276874 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 277494 532226
rect 276874 532102 277494 532170
rect 276874 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 277494 532102
rect 276874 531978 277494 532046
rect 276874 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 277494 531978
rect 276874 514350 277494 531922
rect 276874 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 277494 514350
rect 276874 514226 277494 514294
rect 276874 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 277494 514226
rect 276874 514102 277494 514170
rect 276874 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 277494 514102
rect 276874 513978 277494 514046
rect 276874 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 277494 513978
rect 276874 499846 277494 513922
rect 291154 597212 291774 598268
rect 291154 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 291774 597212
rect 291154 597088 291774 597156
rect 291154 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 291774 597088
rect 291154 596964 291774 597032
rect 291154 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 291774 596964
rect 291154 596840 291774 596908
rect 291154 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 291774 596840
rect 291154 580350 291774 596784
rect 291154 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 291774 580350
rect 291154 580226 291774 580294
rect 291154 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 291774 580226
rect 291154 580102 291774 580170
rect 291154 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 291774 580102
rect 291154 579978 291774 580046
rect 291154 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 291774 579978
rect 291154 562350 291774 579922
rect 291154 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 291774 562350
rect 291154 562226 291774 562294
rect 291154 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 291774 562226
rect 291154 562102 291774 562170
rect 291154 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 291774 562102
rect 291154 561978 291774 562046
rect 291154 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 291774 561978
rect 291154 544350 291774 561922
rect 291154 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 291774 544350
rect 291154 544226 291774 544294
rect 291154 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 291774 544226
rect 291154 544102 291774 544170
rect 291154 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 291774 544102
rect 291154 543978 291774 544046
rect 291154 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 291774 543978
rect 291154 526350 291774 543922
rect 291154 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 291774 526350
rect 291154 526226 291774 526294
rect 291154 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 291774 526226
rect 291154 526102 291774 526170
rect 291154 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 291774 526102
rect 291154 525978 291774 526046
rect 291154 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 291774 525978
rect 291154 508350 291774 525922
rect 291154 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 291774 508350
rect 291154 508226 291774 508294
rect 291154 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 291774 508226
rect 291154 508102 291774 508170
rect 291154 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 291774 508102
rect 291154 507978 291774 508046
rect 291154 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 291774 507978
rect 291154 499846 291774 507922
rect 294874 598172 295494 598268
rect 294874 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 295494 598172
rect 294874 598048 295494 598116
rect 294874 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 295494 598048
rect 294874 597924 295494 597992
rect 294874 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 295494 597924
rect 294874 597800 295494 597868
rect 294874 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 295494 597800
rect 294874 586350 295494 597744
rect 294874 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 295494 586350
rect 294874 586226 295494 586294
rect 294874 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 295494 586226
rect 294874 586102 295494 586170
rect 294874 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 295494 586102
rect 294874 585978 295494 586046
rect 294874 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 295494 585978
rect 294874 568350 295494 585922
rect 294874 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 295494 568350
rect 294874 568226 295494 568294
rect 294874 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 295494 568226
rect 294874 568102 295494 568170
rect 294874 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 295494 568102
rect 294874 567978 295494 568046
rect 294874 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 295494 567978
rect 294874 550350 295494 567922
rect 294874 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 295494 550350
rect 294874 550226 295494 550294
rect 294874 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 295494 550226
rect 294874 550102 295494 550170
rect 294874 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 295494 550102
rect 294874 549978 295494 550046
rect 294874 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 295494 549978
rect 294874 532350 295494 549922
rect 294874 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 295494 532350
rect 294874 532226 295494 532294
rect 294874 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 295494 532226
rect 294874 532102 295494 532170
rect 294874 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 295494 532102
rect 294874 531978 295494 532046
rect 294874 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 295494 531978
rect 294874 514350 295494 531922
rect 294874 514294 294970 514350
rect 295026 514294 295094 514350
rect 295150 514294 295218 514350
rect 295274 514294 295342 514350
rect 295398 514294 295494 514350
rect 294874 514226 295494 514294
rect 294874 514170 294970 514226
rect 295026 514170 295094 514226
rect 295150 514170 295218 514226
rect 295274 514170 295342 514226
rect 295398 514170 295494 514226
rect 294874 514102 295494 514170
rect 294874 514046 294970 514102
rect 295026 514046 295094 514102
rect 295150 514046 295218 514102
rect 295274 514046 295342 514102
rect 295398 514046 295494 514102
rect 294874 513978 295494 514046
rect 294874 513922 294970 513978
rect 295026 513922 295094 513978
rect 295150 513922 295218 513978
rect 295274 513922 295342 513978
rect 295398 513922 295494 513978
rect 294874 499846 295494 513922
rect 309154 597212 309774 598268
rect 309154 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 309774 597212
rect 309154 597088 309774 597156
rect 309154 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 309774 597088
rect 309154 596964 309774 597032
rect 309154 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 309774 596964
rect 309154 596840 309774 596908
rect 309154 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 309774 596840
rect 309154 580350 309774 596784
rect 309154 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 309774 580350
rect 309154 580226 309774 580294
rect 309154 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 309774 580226
rect 309154 580102 309774 580170
rect 309154 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 309774 580102
rect 309154 579978 309774 580046
rect 309154 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 309774 579978
rect 309154 562350 309774 579922
rect 309154 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 309774 562350
rect 309154 562226 309774 562294
rect 309154 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 309774 562226
rect 309154 562102 309774 562170
rect 309154 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 309774 562102
rect 309154 561978 309774 562046
rect 309154 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 309774 561978
rect 309154 544350 309774 561922
rect 309154 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 309774 544350
rect 309154 544226 309774 544294
rect 309154 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 309774 544226
rect 309154 544102 309774 544170
rect 309154 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 309774 544102
rect 309154 543978 309774 544046
rect 309154 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 309774 543978
rect 309154 526350 309774 543922
rect 309154 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 309774 526350
rect 309154 526226 309774 526294
rect 309154 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 309774 526226
rect 309154 526102 309774 526170
rect 309154 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 309774 526102
rect 309154 525978 309774 526046
rect 309154 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 309774 525978
rect 309154 508350 309774 525922
rect 309154 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 309774 508350
rect 309154 508226 309774 508294
rect 309154 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 309774 508226
rect 309154 508102 309774 508170
rect 309154 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 309774 508102
rect 309154 507978 309774 508046
rect 309154 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 309774 507978
rect 309154 499846 309774 507922
rect 312874 598172 313494 598268
rect 312874 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 313494 598172
rect 312874 598048 313494 598116
rect 312874 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 313494 598048
rect 312874 597924 313494 597992
rect 312874 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 313494 597924
rect 312874 597800 313494 597868
rect 312874 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 313494 597800
rect 312874 586350 313494 597744
rect 312874 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 313494 586350
rect 312874 586226 313494 586294
rect 312874 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 313494 586226
rect 312874 586102 313494 586170
rect 312874 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 313494 586102
rect 312874 585978 313494 586046
rect 312874 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 313494 585978
rect 312874 568350 313494 585922
rect 312874 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 313494 568350
rect 312874 568226 313494 568294
rect 312874 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 313494 568226
rect 312874 568102 313494 568170
rect 312874 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 313494 568102
rect 312874 567978 313494 568046
rect 312874 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 313494 567978
rect 312874 550350 313494 567922
rect 312874 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 313494 550350
rect 312874 550226 313494 550294
rect 312874 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 313494 550226
rect 312874 550102 313494 550170
rect 312874 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 313494 550102
rect 312874 549978 313494 550046
rect 312874 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 313494 549978
rect 312874 532350 313494 549922
rect 312874 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 313494 532350
rect 312874 532226 313494 532294
rect 312874 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 313494 532226
rect 312874 532102 313494 532170
rect 312874 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 313494 532102
rect 312874 531978 313494 532046
rect 312874 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 313494 531978
rect 312874 514350 313494 531922
rect 312874 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 313494 514350
rect 312874 514226 313494 514294
rect 312874 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 313494 514226
rect 312874 514102 313494 514170
rect 312874 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 313494 514102
rect 312874 513978 313494 514046
rect 312874 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 313494 513978
rect 312874 499846 313494 513922
rect 327154 597212 327774 598268
rect 327154 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 327774 597212
rect 327154 597088 327774 597156
rect 327154 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 327774 597088
rect 327154 596964 327774 597032
rect 327154 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 327774 596964
rect 327154 596840 327774 596908
rect 327154 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 327774 596840
rect 327154 580350 327774 596784
rect 327154 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 327774 580350
rect 327154 580226 327774 580294
rect 327154 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 327774 580226
rect 327154 580102 327774 580170
rect 327154 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 327774 580102
rect 327154 579978 327774 580046
rect 327154 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 327774 579978
rect 327154 562350 327774 579922
rect 327154 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 327774 562350
rect 327154 562226 327774 562294
rect 327154 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 327774 562226
rect 327154 562102 327774 562170
rect 327154 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 327774 562102
rect 327154 561978 327774 562046
rect 327154 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 327774 561978
rect 327154 544350 327774 561922
rect 327154 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 327774 544350
rect 327154 544226 327774 544294
rect 327154 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 327774 544226
rect 327154 544102 327774 544170
rect 327154 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 327774 544102
rect 327154 543978 327774 544046
rect 327154 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 327774 543978
rect 327154 526350 327774 543922
rect 327154 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 327774 526350
rect 327154 526226 327774 526294
rect 327154 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 327774 526226
rect 327154 526102 327774 526170
rect 327154 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 327774 526102
rect 327154 525978 327774 526046
rect 327154 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 327774 525978
rect 327154 508350 327774 525922
rect 327154 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 327774 508350
rect 327154 508226 327774 508294
rect 327154 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 327774 508226
rect 327154 508102 327774 508170
rect 327154 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 327774 508102
rect 327154 507978 327774 508046
rect 327154 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 327774 507978
rect 327154 499846 327774 507922
rect 330874 598172 331494 598268
rect 330874 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 331494 598172
rect 330874 598048 331494 598116
rect 330874 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 331494 598048
rect 330874 597924 331494 597992
rect 330874 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 331494 597924
rect 330874 597800 331494 597868
rect 330874 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 331494 597800
rect 330874 586350 331494 597744
rect 330874 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 331494 586350
rect 330874 586226 331494 586294
rect 330874 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 331494 586226
rect 330874 586102 331494 586170
rect 330874 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 331494 586102
rect 330874 585978 331494 586046
rect 330874 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 331494 585978
rect 330874 568350 331494 585922
rect 330874 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 331494 568350
rect 330874 568226 331494 568294
rect 330874 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 331494 568226
rect 330874 568102 331494 568170
rect 330874 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 331494 568102
rect 330874 567978 331494 568046
rect 330874 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 331494 567978
rect 330874 550350 331494 567922
rect 330874 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 331494 550350
rect 330874 550226 331494 550294
rect 330874 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 331494 550226
rect 330874 550102 331494 550170
rect 330874 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 331494 550102
rect 330874 549978 331494 550046
rect 330874 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 331494 549978
rect 330874 532350 331494 549922
rect 330874 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 331494 532350
rect 330874 532226 331494 532294
rect 330874 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 331494 532226
rect 330874 532102 331494 532170
rect 330874 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 331494 532102
rect 330874 531978 331494 532046
rect 330874 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 331494 531978
rect 330874 514350 331494 531922
rect 330874 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 331494 514350
rect 330874 514226 331494 514294
rect 330874 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 331494 514226
rect 330874 514102 331494 514170
rect 330874 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 331494 514102
rect 330874 513978 331494 514046
rect 330874 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 331494 513978
rect 330874 499846 331494 513922
rect 345154 597212 345774 598268
rect 345154 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 345774 597212
rect 345154 597088 345774 597156
rect 345154 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 345774 597088
rect 345154 596964 345774 597032
rect 345154 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 345774 596964
rect 345154 596840 345774 596908
rect 345154 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 345774 596840
rect 345154 580350 345774 596784
rect 345154 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 345774 580350
rect 345154 580226 345774 580294
rect 345154 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 345774 580226
rect 345154 580102 345774 580170
rect 345154 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 345774 580102
rect 345154 579978 345774 580046
rect 345154 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 345774 579978
rect 345154 562350 345774 579922
rect 345154 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 345774 562350
rect 345154 562226 345774 562294
rect 345154 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 345774 562226
rect 345154 562102 345774 562170
rect 345154 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 345774 562102
rect 345154 561978 345774 562046
rect 345154 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 345774 561978
rect 345154 544350 345774 561922
rect 345154 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 345774 544350
rect 345154 544226 345774 544294
rect 345154 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 345774 544226
rect 345154 544102 345774 544170
rect 345154 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 345774 544102
rect 345154 543978 345774 544046
rect 345154 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 345774 543978
rect 345154 526350 345774 543922
rect 345154 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 345774 526350
rect 345154 526226 345774 526294
rect 345154 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 345774 526226
rect 345154 526102 345774 526170
rect 345154 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 345774 526102
rect 345154 525978 345774 526046
rect 345154 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 345774 525978
rect 345154 508350 345774 525922
rect 345154 508294 345250 508350
rect 345306 508294 345374 508350
rect 345430 508294 345498 508350
rect 345554 508294 345622 508350
rect 345678 508294 345774 508350
rect 345154 508226 345774 508294
rect 345154 508170 345250 508226
rect 345306 508170 345374 508226
rect 345430 508170 345498 508226
rect 345554 508170 345622 508226
rect 345678 508170 345774 508226
rect 345154 508102 345774 508170
rect 345154 508046 345250 508102
rect 345306 508046 345374 508102
rect 345430 508046 345498 508102
rect 345554 508046 345622 508102
rect 345678 508046 345774 508102
rect 345154 507978 345774 508046
rect 345154 507922 345250 507978
rect 345306 507922 345374 507978
rect 345430 507922 345498 507978
rect 345554 507922 345622 507978
rect 345678 507922 345774 507978
rect 345154 499846 345774 507922
rect 348874 598172 349494 598268
rect 348874 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 349494 598172
rect 348874 598048 349494 598116
rect 348874 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 349494 598048
rect 348874 597924 349494 597992
rect 348874 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 349494 597924
rect 348874 597800 349494 597868
rect 348874 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 349494 597800
rect 348874 586350 349494 597744
rect 348874 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 349494 586350
rect 348874 586226 349494 586294
rect 348874 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 349494 586226
rect 348874 586102 349494 586170
rect 348874 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 349494 586102
rect 348874 585978 349494 586046
rect 348874 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 349494 585978
rect 348874 568350 349494 585922
rect 348874 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 349494 568350
rect 348874 568226 349494 568294
rect 348874 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 349494 568226
rect 348874 568102 349494 568170
rect 348874 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 349494 568102
rect 348874 567978 349494 568046
rect 348874 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 349494 567978
rect 348874 550350 349494 567922
rect 348874 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 349494 550350
rect 348874 550226 349494 550294
rect 348874 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 349494 550226
rect 348874 550102 349494 550170
rect 348874 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 349494 550102
rect 348874 549978 349494 550046
rect 348874 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 349494 549978
rect 348874 532350 349494 549922
rect 348874 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 349494 532350
rect 348874 532226 349494 532294
rect 348874 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 349494 532226
rect 348874 532102 349494 532170
rect 348874 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 349494 532102
rect 348874 531978 349494 532046
rect 348874 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 349494 531978
rect 348874 514350 349494 531922
rect 348874 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 349494 514350
rect 348874 514226 349494 514294
rect 348874 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 349494 514226
rect 348874 514102 349494 514170
rect 348874 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 349494 514102
rect 348874 513978 349494 514046
rect 348874 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 349494 513978
rect 348874 499846 349494 513922
rect 363154 597212 363774 598268
rect 363154 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 363774 597212
rect 363154 597088 363774 597156
rect 363154 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 363774 597088
rect 363154 596964 363774 597032
rect 363154 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 363774 596964
rect 363154 596840 363774 596908
rect 363154 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 363774 596840
rect 363154 580350 363774 596784
rect 363154 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 363774 580350
rect 363154 580226 363774 580294
rect 363154 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 363774 580226
rect 363154 580102 363774 580170
rect 363154 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 363774 580102
rect 363154 579978 363774 580046
rect 363154 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 363774 579978
rect 363154 562350 363774 579922
rect 363154 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 363774 562350
rect 363154 562226 363774 562294
rect 363154 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 363774 562226
rect 363154 562102 363774 562170
rect 363154 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 363774 562102
rect 363154 561978 363774 562046
rect 363154 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 363774 561978
rect 363154 544350 363774 561922
rect 363154 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 363774 544350
rect 363154 544226 363774 544294
rect 363154 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 363774 544226
rect 363154 544102 363774 544170
rect 363154 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 363774 544102
rect 363154 543978 363774 544046
rect 363154 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 363774 543978
rect 363154 526350 363774 543922
rect 363154 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 363774 526350
rect 363154 526226 363774 526294
rect 363154 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 363774 526226
rect 363154 526102 363774 526170
rect 363154 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 363774 526102
rect 363154 525978 363774 526046
rect 363154 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 363774 525978
rect 363154 508350 363774 525922
rect 363154 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 363774 508350
rect 363154 508226 363774 508294
rect 363154 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 363774 508226
rect 363154 508102 363774 508170
rect 363154 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 363774 508102
rect 363154 507978 363774 508046
rect 363154 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 363774 507978
rect 363154 499846 363774 507922
rect 366874 598172 367494 598268
rect 366874 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 367494 598172
rect 366874 598048 367494 598116
rect 366874 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 367494 598048
rect 366874 597924 367494 597992
rect 366874 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 367494 597924
rect 366874 597800 367494 597868
rect 366874 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 367494 597800
rect 366874 586350 367494 597744
rect 366874 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 367494 586350
rect 366874 586226 367494 586294
rect 366874 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 367494 586226
rect 366874 586102 367494 586170
rect 366874 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 367494 586102
rect 366874 585978 367494 586046
rect 366874 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 367494 585978
rect 366874 568350 367494 585922
rect 366874 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 367494 568350
rect 366874 568226 367494 568294
rect 366874 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 367494 568226
rect 366874 568102 367494 568170
rect 366874 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 367494 568102
rect 366874 567978 367494 568046
rect 366874 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 367494 567978
rect 366874 550350 367494 567922
rect 366874 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 367494 550350
rect 366874 550226 367494 550294
rect 366874 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 367494 550226
rect 366874 550102 367494 550170
rect 366874 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 367494 550102
rect 366874 549978 367494 550046
rect 366874 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 367494 549978
rect 366874 532350 367494 549922
rect 366874 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 367494 532350
rect 366874 532226 367494 532294
rect 366874 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 367494 532226
rect 366874 532102 367494 532170
rect 366874 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 367494 532102
rect 366874 531978 367494 532046
rect 366874 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 367494 531978
rect 366874 514350 367494 531922
rect 366874 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 367494 514350
rect 366874 514226 367494 514294
rect 366874 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 367494 514226
rect 366874 514102 367494 514170
rect 366874 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 367494 514102
rect 366874 513978 367494 514046
rect 366874 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 367494 513978
rect 366874 499846 367494 513922
rect 381154 597212 381774 598268
rect 381154 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 381774 597212
rect 381154 597088 381774 597156
rect 381154 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 381774 597088
rect 381154 596964 381774 597032
rect 381154 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 381774 596964
rect 381154 596840 381774 596908
rect 381154 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 381774 596840
rect 381154 580350 381774 596784
rect 381154 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 381774 580350
rect 381154 580226 381774 580294
rect 381154 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 381774 580226
rect 381154 580102 381774 580170
rect 381154 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 381774 580102
rect 381154 579978 381774 580046
rect 381154 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 381774 579978
rect 381154 562350 381774 579922
rect 381154 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 381774 562350
rect 381154 562226 381774 562294
rect 381154 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 381774 562226
rect 381154 562102 381774 562170
rect 381154 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 381774 562102
rect 381154 561978 381774 562046
rect 381154 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 381774 561978
rect 381154 544350 381774 561922
rect 381154 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 381774 544350
rect 381154 544226 381774 544294
rect 381154 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 381774 544226
rect 381154 544102 381774 544170
rect 381154 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 381774 544102
rect 381154 543978 381774 544046
rect 381154 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 381774 543978
rect 381154 526350 381774 543922
rect 381154 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 381774 526350
rect 381154 526226 381774 526294
rect 381154 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 381774 526226
rect 381154 526102 381774 526170
rect 381154 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 381774 526102
rect 381154 525978 381774 526046
rect 381154 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 381774 525978
rect 381154 508350 381774 525922
rect 381154 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 381774 508350
rect 381154 508226 381774 508294
rect 381154 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 381774 508226
rect 381154 508102 381774 508170
rect 381154 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 381774 508102
rect 381154 507978 381774 508046
rect 381154 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 381774 507978
rect 381154 499846 381774 507922
rect 384874 598172 385494 598268
rect 384874 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 385494 598172
rect 384874 598048 385494 598116
rect 384874 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 385494 598048
rect 384874 597924 385494 597992
rect 384874 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 385494 597924
rect 384874 597800 385494 597868
rect 384874 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 385494 597800
rect 384874 586350 385494 597744
rect 384874 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 385494 586350
rect 384874 586226 385494 586294
rect 384874 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 385494 586226
rect 384874 586102 385494 586170
rect 384874 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 385494 586102
rect 384874 585978 385494 586046
rect 384874 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 385494 585978
rect 384874 568350 385494 585922
rect 384874 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 385494 568350
rect 384874 568226 385494 568294
rect 384874 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 385494 568226
rect 384874 568102 385494 568170
rect 384874 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 385494 568102
rect 384874 567978 385494 568046
rect 384874 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 385494 567978
rect 384874 550350 385494 567922
rect 384874 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 385494 550350
rect 384874 550226 385494 550294
rect 384874 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 385494 550226
rect 384874 550102 385494 550170
rect 384874 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 385494 550102
rect 384874 549978 385494 550046
rect 384874 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 385494 549978
rect 384874 532350 385494 549922
rect 384874 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 385494 532350
rect 384874 532226 385494 532294
rect 384874 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 385494 532226
rect 384874 532102 385494 532170
rect 384874 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 385494 532102
rect 384874 531978 385494 532046
rect 384874 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 385494 531978
rect 384874 514350 385494 531922
rect 384874 514294 384970 514350
rect 385026 514294 385094 514350
rect 385150 514294 385218 514350
rect 385274 514294 385342 514350
rect 385398 514294 385494 514350
rect 384874 514226 385494 514294
rect 384874 514170 384970 514226
rect 385026 514170 385094 514226
rect 385150 514170 385218 514226
rect 385274 514170 385342 514226
rect 385398 514170 385494 514226
rect 384874 514102 385494 514170
rect 384874 514046 384970 514102
rect 385026 514046 385094 514102
rect 385150 514046 385218 514102
rect 385274 514046 385342 514102
rect 385398 514046 385494 514102
rect 384874 513978 385494 514046
rect 384874 513922 384970 513978
rect 385026 513922 385094 513978
rect 385150 513922 385218 513978
rect 385274 513922 385342 513978
rect 385398 513922 385494 513978
rect 384874 499846 385494 513922
rect 399154 597212 399774 598268
rect 399154 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 399774 597212
rect 399154 597088 399774 597156
rect 399154 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 399774 597088
rect 399154 596964 399774 597032
rect 399154 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 399774 596964
rect 399154 596840 399774 596908
rect 399154 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 399774 596840
rect 399154 580350 399774 596784
rect 399154 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 399774 580350
rect 399154 580226 399774 580294
rect 399154 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 399774 580226
rect 399154 580102 399774 580170
rect 399154 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 399774 580102
rect 399154 579978 399774 580046
rect 399154 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 399774 579978
rect 399154 562350 399774 579922
rect 399154 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 399774 562350
rect 399154 562226 399774 562294
rect 399154 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 399774 562226
rect 399154 562102 399774 562170
rect 399154 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 399774 562102
rect 399154 561978 399774 562046
rect 399154 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 399774 561978
rect 399154 544350 399774 561922
rect 399154 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 399774 544350
rect 399154 544226 399774 544294
rect 399154 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 399774 544226
rect 399154 544102 399774 544170
rect 399154 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 399774 544102
rect 399154 543978 399774 544046
rect 399154 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 399774 543978
rect 399154 526350 399774 543922
rect 399154 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 399774 526350
rect 399154 526226 399774 526294
rect 399154 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 399774 526226
rect 399154 526102 399774 526170
rect 399154 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 399774 526102
rect 399154 525978 399774 526046
rect 399154 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 399774 525978
rect 399154 508350 399774 525922
rect 399154 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 399774 508350
rect 399154 508226 399774 508294
rect 399154 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 399774 508226
rect 399154 508102 399774 508170
rect 399154 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 399774 508102
rect 399154 507978 399774 508046
rect 399154 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 399774 507978
rect 399154 499846 399774 507922
rect 402874 598172 403494 598268
rect 402874 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 403494 598172
rect 402874 598048 403494 598116
rect 402874 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 403494 598048
rect 402874 597924 403494 597992
rect 402874 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 403494 597924
rect 402874 597800 403494 597868
rect 402874 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 403494 597800
rect 402874 586350 403494 597744
rect 402874 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 403494 586350
rect 402874 586226 403494 586294
rect 402874 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 403494 586226
rect 402874 586102 403494 586170
rect 402874 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 403494 586102
rect 402874 585978 403494 586046
rect 402874 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 403494 585978
rect 402874 568350 403494 585922
rect 402874 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 403494 568350
rect 402874 568226 403494 568294
rect 402874 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 403494 568226
rect 402874 568102 403494 568170
rect 402874 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 403494 568102
rect 402874 567978 403494 568046
rect 402874 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 403494 567978
rect 402874 550350 403494 567922
rect 402874 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 403494 550350
rect 402874 550226 403494 550294
rect 402874 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 403494 550226
rect 402874 550102 403494 550170
rect 402874 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 403494 550102
rect 402874 549978 403494 550046
rect 402874 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 403494 549978
rect 402874 532350 403494 549922
rect 402874 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 403494 532350
rect 402874 532226 403494 532294
rect 402874 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 403494 532226
rect 402874 532102 403494 532170
rect 402874 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 403494 532102
rect 402874 531978 403494 532046
rect 402874 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 403494 531978
rect 402874 514350 403494 531922
rect 402874 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 403494 514350
rect 402874 514226 403494 514294
rect 402874 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 403494 514226
rect 402874 514102 403494 514170
rect 402874 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 403494 514102
rect 402874 513978 403494 514046
rect 402874 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 403494 513978
rect 402874 499846 403494 513922
rect 417154 597212 417774 598268
rect 417154 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 417774 597212
rect 417154 597088 417774 597156
rect 417154 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 417774 597088
rect 417154 596964 417774 597032
rect 417154 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 417774 596964
rect 417154 596840 417774 596908
rect 417154 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 417774 596840
rect 417154 580350 417774 596784
rect 417154 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 417774 580350
rect 417154 580226 417774 580294
rect 417154 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 417774 580226
rect 417154 580102 417774 580170
rect 417154 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 417774 580102
rect 417154 579978 417774 580046
rect 417154 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 417774 579978
rect 417154 562350 417774 579922
rect 417154 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 417774 562350
rect 417154 562226 417774 562294
rect 417154 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 417774 562226
rect 417154 562102 417774 562170
rect 417154 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 417774 562102
rect 417154 561978 417774 562046
rect 417154 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 417774 561978
rect 417154 544350 417774 561922
rect 417154 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 417774 544350
rect 417154 544226 417774 544294
rect 417154 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 417774 544226
rect 417154 544102 417774 544170
rect 417154 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 417774 544102
rect 417154 543978 417774 544046
rect 417154 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 417774 543978
rect 417154 526350 417774 543922
rect 417154 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 417774 526350
rect 417154 526226 417774 526294
rect 417154 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 417774 526226
rect 417154 526102 417774 526170
rect 417154 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 417774 526102
rect 417154 525978 417774 526046
rect 417154 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 417774 525978
rect 417154 508350 417774 525922
rect 417154 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 417774 508350
rect 417154 508226 417774 508294
rect 417154 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 417774 508226
rect 417154 508102 417774 508170
rect 417154 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 417774 508102
rect 417154 507978 417774 508046
rect 417154 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 417774 507978
rect 417154 499846 417774 507922
rect 420874 598172 421494 598268
rect 420874 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 421494 598172
rect 420874 598048 421494 598116
rect 420874 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 421494 598048
rect 420874 597924 421494 597992
rect 420874 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 421494 597924
rect 420874 597800 421494 597868
rect 420874 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 421494 597800
rect 420874 586350 421494 597744
rect 420874 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 421494 586350
rect 420874 586226 421494 586294
rect 420874 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 421494 586226
rect 420874 586102 421494 586170
rect 420874 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 421494 586102
rect 420874 585978 421494 586046
rect 420874 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 421494 585978
rect 420874 568350 421494 585922
rect 420874 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 421494 568350
rect 420874 568226 421494 568294
rect 420874 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 421494 568226
rect 420874 568102 421494 568170
rect 420874 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 421494 568102
rect 420874 567978 421494 568046
rect 420874 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 421494 567978
rect 420874 550350 421494 567922
rect 420874 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 421494 550350
rect 420874 550226 421494 550294
rect 420874 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 421494 550226
rect 420874 550102 421494 550170
rect 420874 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 421494 550102
rect 420874 549978 421494 550046
rect 420874 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 421494 549978
rect 420874 532350 421494 549922
rect 420874 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 421494 532350
rect 420874 532226 421494 532294
rect 420874 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 421494 532226
rect 420874 532102 421494 532170
rect 420874 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 421494 532102
rect 420874 531978 421494 532046
rect 420874 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 421494 531978
rect 420874 514350 421494 531922
rect 420874 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 421494 514350
rect 420874 514226 421494 514294
rect 420874 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 421494 514226
rect 420874 514102 421494 514170
rect 420874 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 421494 514102
rect 420874 513978 421494 514046
rect 420874 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 421494 513978
rect 420874 499846 421494 513922
rect 435154 597212 435774 598268
rect 435154 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 435774 597212
rect 435154 597088 435774 597156
rect 435154 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 435774 597088
rect 435154 596964 435774 597032
rect 435154 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 435774 596964
rect 435154 596840 435774 596908
rect 435154 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 435774 596840
rect 435154 580350 435774 596784
rect 435154 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 435774 580350
rect 435154 580226 435774 580294
rect 435154 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 435774 580226
rect 435154 580102 435774 580170
rect 435154 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 435774 580102
rect 435154 579978 435774 580046
rect 435154 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 435774 579978
rect 435154 562350 435774 579922
rect 435154 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 435774 562350
rect 435154 562226 435774 562294
rect 435154 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 435774 562226
rect 435154 562102 435774 562170
rect 435154 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 435774 562102
rect 435154 561978 435774 562046
rect 435154 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 435774 561978
rect 435154 544350 435774 561922
rect 435154 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 435774 544350
rect 435154 544226 435774 544294
rect 435154 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 435774 544226
rect 435154 544102 435774 544170
rect 435154 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 435774 544102
rect 435154 543978 435774 544046
rect 435154 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 435774 543978
rect 435154 526350 435774 543922
rect 435154 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 435774 526350
rect 435154 526226 435774 526294
rect 435154 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 435774 526226
rect 435154 526102 435774 526170
rect 435154 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 435774 526102
rect 435154 525978 435774 526046
rect 435154 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 435774 525978
rect 435154 508350 435774 525922
rect 435154 508294 435250 508350
rect 435306 508294 435374 508350
rect 435430 508294 435498 508350
rect 435554 508294 435622 508350
rect 435678 508294 435774 508350
rect 435154 508226 435774 508294
rect 435154 508170 435250 508226
rect 435306 508170 435374 508226
rect 435430 508170 435498 508226
rect 435554 508170 435622 508226
rect 435678 508170 435774 508226
rect 435154 508102 435774 508170
rect 435154 508046 435250 508102
rect 435306 508046 435374 508102
rect 435430 508046 435498 508102
rect 435554 508046 435622 508102
rect 435678 508046 435774 508102
rect 435154 507978 435774 508046
rect 435154 507922 435250 507978
rect 435306 507922 435374 507978
rect 435430 507922 435498 507978
rect 435554 507922 435622 507978
rect 435678 507922 435774 507978
rect 435154 499846 435774 507922
rect 438874 598172 439494 598268
rect 438874 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 439494 598172
rect 438874 598048 439494 598116
rect 438874 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 439494 598048
rect 438874 597924 439494 597992
rect 438874 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 439494 597924
rect 438874 597800 439494 597868
rect 438874 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 439494 597800
rect 438874 586350 439494 597744
rect 438874 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 439494 586350
rect 438874 586226 439494 586294
rect 438874 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 439494 586226
rect 438874 586102 439494 586170
rect 438874 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 439494 586102
rect 438874 585978 439494 586046
rect 438874 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 439494 585978
rect 438874 568350 439494 585922
rect 438874 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 439494 568350
rect 438874 568226 439494 568294
rect 438874 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 439494 568226
rect 438874 568102 439494 568170
rect 438874 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 439494 568102
rect 438874 567978 439494 568046
rect 438874 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 439494 567978
rect 438874 550350 439494 567922
rect 438874 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 439494 550350
rect 438874 550226 439494 550294
rect 438874 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 439494 550226
rect 438874 550102 439494 550170
rect 438874 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 439494 550102
rect 438874 549978 439494 550046
rect 438874 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 439494 549978
rect 438874 532350 439494 549922
rect 438874 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 439494 532350
rect 438874 532226 439494 532294
rect 438874 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 439494 532226
rect 438874 532102 439494 532170
rect 438874 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 439494 532102
rect 438874 531978 439494 532046
rect 438874 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 439494 531978
rect 438874 514350 439494 531922
rect 438874 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 439494 514350
rect 438874 514226 439494 514294
rect 438874 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 439494 514226
rect 438874 514102 439494 514170
rect 438874 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 439494 514102
rect 438874 513978 439494 514046
rect 438874 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 439494 513978
rect 438874 499846 439494 513922
rect 453154 597212 453774 598268
rect 453154 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 453774 597212
rect 453154 597088 453774 597156
rect 453154 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 453774 597088
rect 453154 596964 453774 597032
rect 453154 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 453774 596964
rect 453154 596840 453774 596908
rect 453154 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 453774 596840
rect 453154 580350 453774 596784
rect 453154 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 453774 580350
rect 453154 580226 453774 580294
rect 453154 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 453774 580226
rect 453154 580102 453774 580170
rect 453154 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 453774 580102
rect 453154 579978 453774 580046
rect 453154 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 453774 579978
rect 453154 562350 453774 579922
rect 453154 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 453774 562350
rect 453154 562226 453774 562294
rect 453154 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 453774 562226
rect 453154 562102 453774 562170
rect 453154 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 453774 562102
rect 453154 561978 453774 562046
rect 453154 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 453774 561978
rect 453154 544350 453774 561922
rect 453154 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 453774 544350
rect 453154 544226 453774 544294
rect 453154 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 453774 544226
rect 453154 544102 453774 544170
rect 453154 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 453774 544102
rect 453154 543978 453774 544046
rect 453154 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 453774 543978
rect 453154 526350 453774 543922
rect 453154 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 453774 526350
rect 453154 526226 453774 526294
rect 453154 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 453774 526226
rect 453154 526102 453774 526170
rect 453154 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 453774 526102
rect 453154 525978 453774 526046
rect 453154 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 453774 525978
rect 453154 508350 453774 525922
rect 453154 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 453774 508350
rect 453154 508226 453774 508294
rect 453154 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 453774 508226
rect 453154 508102 453774 508170
rect 453154 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 453774 508102
rect 453154 507978 453774 508046
rect 453154 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 453774 507978
rect 453154 499846 453774 507922
rect 456874 598172 457494 598268
rect 456874 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 457494 598172
rect 456874 598048 457494 598116
rect 456874 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 457494 598048
rect 456874 597924 457494 597992
rect 456874 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 457494 597924
rect 456874 597800 457494 597868
rect 456874 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 457494 597800
rect 456874 586350 457494 597744
rect 456874 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 457494 586350
rect 456874 586226 457494 586294
rect 456874 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 457494 586226
rect 456874 586102 457494 586170
rect 456874 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 457494 586102
rect 456874 585978 457494 586046
rect 456874 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 457494 585978
rect 456874 568350 457494 585922
rect 456874 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 457494 568350
rect 456874 568226 457494 568294
rect 456874 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 457494 568226
rect 456874 568102 457494 568170
rect 456874 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 457494 568102
rect 456874 567978 457494 568046
rect 456874 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 457494 567978
rect 456874 550350 457494 567922
rect 456874 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 457494 550350
rect 456874 550226 457494 550294
rect 456874 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 457494 550226
rect 456874 550102 457494 550170
rect 456874 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 457494 550102
rect 456874 549978 457494 550046
rect 456874 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 457494 549978
rect 456874 532350 457494 549922
rect 456874 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 457494 532350
rect 456874 532226 457494 532294
rect 456874 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 457494 532226
rect 456874 532102 457494 532170
rect 456874 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 457494 532102
rect 456874 531978 457494 532046
rect 456874 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 457494 531978
rect 456874 514350 457494 531922
rect 456874 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 457494 514350
rect 456874 514226 457494 514294
rect 456874 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 457494 514226
rect 456874 514102 457494 514170
rect 456874 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 457494 514102
rect 456874 513978 457494 514046
rect 456874 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 457494 513978
rect 456874 499846 457494 513922
rect 471154 597212 471774 598268
rect 471154 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 471774 597212
rect 471154 597088 471774 597156
rect 471154 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 471774 597088
rect 471154 596964 471774 597032
rect 471154 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 471774 596964
rect 471154 596840 471774 596908
rect 471154 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 471774 596840
rect 471154 580350 471774 596784
rect 471154 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 471774 580350
rect 471154 580226 471774 580294
rect 471154 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 471774 580226
rect 471154 580102 471774 580170
rect 471154 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 471774 580102
rect 471154 579978 471774 580046
rect 471154 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 471774 579978
rect 471154 562350 471774 579922
rect 471154 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 471774 562350
rect 471154 562226 471774 562294
rect 471154 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 471774 562226
rect 471154 562102 471774 562170
rect 471154 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 471774 562102
rect 471154 561978 471774 562046
rect 471154 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 471774 561978
rect 471154 544350 471774 561922
rect 471154 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 471774 544350
rect 471154 544226 471774 544294
rect 471154 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 471774 544226
rect 471154 544102 471774 544170
rect 471154 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 471774 544102
rect 471154 543978 471774 544046
rect 471154 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 471774 543978
rect 471154 526350 471774 543922
rect 471154 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 471774 526350
rect 471154 526226 471774 526294
rect 471154 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 471774 526226
rect 471154 526102 471774 526170
rect 471154 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 471774 526102
rect 471154 525978 471774 526046
rect 471154 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 471774 525978
rect 471154 508350 471774 525922
rect 471154 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 471774 508350
rect 471154 508226 471774 508294
rect 471154 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 471774 508226
rect 471154 508102 471774 508170
rect 471154 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 471774 508102
rect 471154 507978 471774 508046
rect 471154 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 471774 507978
rect 471154 499846 471774 507922
rect 474874 598172 475494 598268
rect 474874 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 475494 598172
rect 474874 598048 475494 598116
rect 474874 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 475494 598048
rect 474874 597924 475494 597992
rect 474874 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 475494 597924
rect 474874 597800 475494 597868
rect 474874 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 475494 597800
rect 474874 586350 475494 597744
rect 474874 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 475494 586350
rect 474874 586226 475494 586294
rect 474874 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 475494 586226
rect 474874 586102 475494 586170
rect 474874 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 475494 586102
rect 474874 585978 475494 586046
rect 474874 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 475494 585978
rect 474874 568350 475494 585922
rect 474874 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 475494 568350
rect 474874 568226 475494 568294
rect 474874 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 475494 568226
rect 474874 568102 475494 568170
rect 474874 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 475494 568102
rect 474874 567978 475494 568046
rect 474874 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 475494 567978
rect 474874 550350 475494 567922
rect 474874 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 475494 550350
rect 474874 550226 475494 550294
rect 474874 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 475494 550226
rect 474874 550102 475494 550170
rect 474874 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 475494 550102
rect 474874 549978 475494 550046
rect 474874 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 475494 549978
rect 474874 532350 475494 549922
rect 474874 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 475494 532350
rect 474874 532226 475494 532294
rect 474874 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 475494 532226
rect 474874 532102 475494 532170
rect 474874 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 475494 532102
rect 474874 531978 475494 532046
rect 474874 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 475494 531978
rect 474874 514350 475494 531922
rect 474874 514294 474970 514350
rect 475026 514294 475094 514350
rect 475150 514294 475218 514350
rect 475274 514294 475342 514350
rect 475398 514294 475494 514350
rect 474874 514226 475494 514294
rect 474874 514170 474970 514226
rect 475026 514170 475094 514226
rect 475150 514170 475218 514226
rect 475274 514170 475342 514226
rect 475398 514170 475494 514226
rect 474874 514102 475494 514170
rect 474874 514046 474970 514102
rect 475026 514046 475094 514102
rect 475150 514046 475218 514102
rect 475274 514046 475342 514102
rect 475398 514046 475494 514102
rect 474874 513978 475494 514046
rect 474874 513922 474970 513978
rect 475026 513922 475094 513978
rect 475150 513922 475218 513978
rect 475274 513922 475342 513978
rect 475398 513922 475494 513978
rect 474874 499846 475494 513922
rect 489154 597212 489774 598268
rect 489154 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 489774 597212
rect 489154 597088 489774 597156
rect 489154 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 489774 597088
rect 489154 596964 489774 597032
rect 489154 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 489774 596964
rect 489154 596840 489774 596908
rect 489154 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 489774 596840
rect 489154 580350 489774 596784
rect 489154 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 489774 580350
rect 489154 580226 489774 580294
rect 489154 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 489774 580226
rect 489154 580102 489774 580170
rect 489154 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 489774 580102
rect 489154 579978 489774 580046
rect 489154 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 489774 579978
rect 489154 562350 489774 579922
rect 489154 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 489774 562350
rect 489154 562226 489774 562294
rect 489154 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 489774 562226
rect 489154 562102 489774 562170
rect 489154 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 489774 562102
rect 489154 561978 489774 562046
rect 489154 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 489774 561978
rect 489154 544350 489774 561922
rect 489154 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 489774 544350
rect 489154 544226 489774 544294
rect 489154 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 489774 544226
rect 489154 544102 489774 544170
rect 489154 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 489774 544102
rect 489154 543978 489774 544046
rect 489154 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 489774 543978
rect 489154 526350 489774 543922
rect 489154 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 489774 526350
rect 489154 526226 489774 526294
rect 489154 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 489774 526226
rect 489154 526102 489774 526170
rect 489154 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 489774 526102
rect 489154 525978 489774 526046
rect 489154 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 489774 525978
rect 489154 508350 489774 525922
rect 489154 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 489774 508350
rect 489154 508226 489774 508294
rect 489154 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 489774 508226
rect 489154 508102 489774 508170
rect 489154 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 489774 508102
rect 489154 507978 489774 508046
rect 489154 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 489774 507978
rect 489154 499846 489774 507922
rect 492874 598172 493494 598268
rect 492874 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 493494 598172
rect 492874 598048 493494 598116
rect 492874 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 493494 598048
rect 492874 597924 493494 597992
rect 492874 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 493494 597924
rect 492874 597800 493494 597868
rect 492874 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 493494 597800
rect 492874 586350 493494 597744
rect 492874 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 493494 586350
rect 492874 586226 493494 586294
rect 492874 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 493494 586226
rect 492874 586102 493494 586170
rect 492874 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 493494 586102
rect 492874 585978 493494 586046
rect 492874 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 493494 585978
rect 492874 568350 493494 585922
rect 492874 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 493494 568350
rect 492874 568226 493494 568294
rect 492874 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 493494 568226
rect 492874 568102 493494 568170
rect 492874 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 493494 568102
rect 492874 567978 493494 568046
rect 492874 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 493494 567978
rect 492874 550350 493494 567922
rect 492874 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 493494 550350
rect 492874 550226 493494 550294
rect 492874 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 493494 550226
rect 492874 550102 493494 550170
rect 492874 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 493494 550102
rect 492874 549978 493494 550046
rect 492874 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 493494 549978
rect 492874 532350 493494 549922
rect 492874 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 493494 532350
rect 492874 532226 493494 532294
rect 492874 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 493494 532226
rect 492874 532102 493494 532170
rect 492874 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 493494 532102
rect 492874 531978 493494 532046
rect 492874 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 493494 531978
rect 492874 514350 493494 531922
rect 492874 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 493494 514350
rect 492874 514226 493494 514294
rect 492874 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 493494 514226
rect 492874 514102 493494 514170
rect 492874 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 493494 514102
rect 492874 513978 493494 514046
rect 492874 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 493494 513978
rect 492874 499846 493494 513922
rect 507154 597212 507774 598268
rect 507154 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 507774 597212
rect 507154 597088 507774 597156
rect 507154 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 507774 597088
rect 507154 596964 507774 597032
rect 507154 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 507774 596964
rect 507154 596840 507774 596908
rect 507154 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 507774 596840
rect 507154 580350 507774 596784
rect 507154 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 507774 580350
rect 507154 580226 507774 580294
rect 507154 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 507774 580226
rect 507154 580102 507774 580170
rect 507154 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 507774 580102
rect 507154 579978 507774 580046
rect 507154 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 507774 579978
rect 507154 562350 507774 579922
rect 507154 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 507774 562350
rect 507154 562226 507774 562294
rect 507154 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 507774 562226
rect 507154 562102 507774 562170
rect 507154 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 507774 562102
rect 507154 561978 507774 562046
rect 507154 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 507774 561978
rect 507154 544350 507774 561922
rect 507154 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 507774 544350
rect 507154 544226 507774 544294
rect 507154 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 507774 544226
rect 507154 544102 507774 544170
rect 507154 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 507774 544102
rect 507154 543978 507774 544046
rect 507154 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 507774 543978
rect 507154 526350 507774 543922
rect 507154 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 507774 526350
rect 507154 526226 507774 526294
rect 507154 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 507774 526226
rect 507154 526102 507774 526170
rect 507154 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 507774 526102
rect 507154 525978 507774 526046
rect 507154 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 507774 525978
rect 507154 508350 507774 525922
rect 507154 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 507774 508350
rect 507154 508226 507774 508294
rect 507154 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 507774 508226
rect 507154 508102 507774 508170
rect 507154 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 507774 508102
rect 507154 507978 507774 508046
rect 507154 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 507774 507978
rect 467180 499380 467236 499390
rect 412860 499156 412916 499166
rect 413308 499156 413364 499166
rect 412916 499100 413308 499156
rect 412860 499090 412916 499100
rect 413308 499090 413364 499100
rect 467180 499044 467236 499324
rect 467180 498978 467236 498988
rect 219808 496333 220128 496350
rect 219808 496277 219878 496333
rect 219934 496277 220002 496333
rect 220058 496277 220128 496333
rect 219808 496209 220128 496277
rect 219808 496153 219878 496209
rect 219934 496153 220002 496209
rect 220058 496153 220128 496209
rect 219808 496085 220128 496153
rect 219808 496029 219878 496085
rect 219934 496029 220002 496085
rect 220058 496029 220128 496085
rect 219808 495961 220128 496029
rect 219808 495905 219878 495961
rect 219934 495905 220002 495961
rect 220058 495905 220128 495961
rect 219808 495888 220128 495905
rect 250528 496333 250848 496350
rect 250528 496277 250598 496333
rect 250654 496277 250722 496333
rect 250778 496277 250848 496333
rect 250528 496209 250848 496277
rect 250528 496153 250598 496209
rect 250654 496153 250722 496209
rect 250778 496153 250848 496209
rect 250528 496085 250848 496153
rect 250528 496029 250598 496085
rect 250654 496029 250722 496085
rect 250778 496029 250848 496085
rect 250528 495961 250848 496029
rect 250528 495905 250598 495961
rect 250654 495905 250722 495961
rect 250778 495905 250848 495961
rect 250528 495888 250848 495905
rect 281248 496333 281568 496350
rect 281248 496277 281318 496333
rect 281374 496277 281442 496333
rect 281498 496277 281568 496333
rect 281248 496209 281568 496277
rect 281248 496153 281318 496209
rect 281374 496153 281442 496209
rect 281498 496153 281568 496209
rect 281248 496085 281568 496153
rect 281248 496029 281318 496085
rect 281374 496029 281442 496085
rect 281498 496029 281568 496085
rect 281248 495961 281568 496029
rect 281248 495905 281318 495961
rect 281374 495905 281442 495961
rect 281498 495905 281568 495961
rect 281248 495888 281568 495905
rect 311968 496333 312288 496350
rect 311968 496277 312038 496333
rect 312094 496277 312162 496333
rect 312218 496277 312288 496333
rect 311968 496209 312288 496277
rect 311968 496153 312038 496209
rect 312094 496153 312162 496209
rect 312218 496153 312288 496209
rect 311968 496085 312288 496153
rect 311968 496029 312038 496085
rect 312094 496029 312162 496085
rect 312218 496029 312288 496085
rect 311968 495961 312288 496029
rect 311968 495905 312038 495961
rect 312094 495905 312162 495961
rect 312218 495905 312288 495961
rect 311968 495888 312288 495905
rect 342688 496333 343008 496350
rect 342688 496277 342758 496333
rect 342814 496277 342882 496333
rect 342938 496277 343008 496333
rect 342688 496209 343008 496277
rect 342688 496153 342758 496209
rect 342814 496153 342882 496209
rect 342938 496153 343008 496209
rect 342688 496085 343008 496153
rect 342688 496029 342758 496085
rect 342814 496029 342882 496085
rect 342938 496029 343008 496085
rect 342688 495961 343008 496029
rect 342688 495905 342758 495961
rect 342814 495905 342882 495961
rect 342938 495905 343008 495961
rect 342688 495888 343008 495905
rect 373408 496333 373728 496350
rect 373408 496277 373478 496333
rect 373534 496277 373602 496333
rect 373658 496277 373728 496333
rect 373408 496209 373728 496277
rect 373408 496153 373478 496209
rect 373534 496153 373602 496209
rect 373658 496153 373728 496209
rect 373408 496085 373728 496153
rect 373408 496029 373478 496085
rect 373534 496029 373602 496085
rect 373658 496029 373728 496085
rect 373408 495961 373728 496029
rect 373408 495905 373478 495961
rect 373534 495905 373602 495961
rect 373658 495905 373728 495961
rect 373408 495888 373728 495905
rect 404128 496333 404448 496350
rect 404128 496277 404198 496333
rect 404254 496277 404322 496333
rect 404378 496277 404448 496333
rect 404128 496209 404448 496277
rect 404128 496153 404198 496209
rect 404254 496153 404322 496209
rect 404378 496153 404448 496209
rect 404128 496085 404448 496153
rect 404128 496029 404198 496085
rect 404254 496029 404322 496085
rect 404378 496029 404448 496085
rect 404128 495961 404448 496029
rect 404128 495905 404198 495961
rect 404254 495905 404322 495961
rect 404378 495905 404448 495961
rect 404128 495888 404448 495905
rect 434848 496333 435168 496350
rect 434848 496277 434918 496333
rect 434974 496277 435042 496333
rect 435098 496277 435168 496333
rect 434848 496209 435168 496277
rect 434848 496153 434918 496209
rect 434974 496153 435042 496209
rect 435098 496153 435168 496209
rect 434848 496085 435168 496153
rect 434848 496029 434918 496085
rect 434974 496029 435042 496085
rect 435098 496029 435168 496085
rect 434848 495961 435168 496029
rect 434848 495905 434918 495961
rect 434974 495905 435042 495961
rect 435098 495905 435168 495961
rect 434848 495888 435168 495905
rect 465568 496333 465888 496350
rect 465568 496277 465638 496333
rect 465694 496277 465762 496333
rect 465818 496277 465888 496333
rect 465568 496209 465888 496277
rect 465568 496153 465638 496209
rect 465694 496153 465762 496209
rect 465818 496153 465888 496209
rect 465568 496085 465888 496153
rect 465568 496029 465638 496085
rect 465694 496029 465762 496085
rect 465818 496029 465888 496085
rect 465568 495961 465888 496029
rect 465568 495905 465638 495961
rect 465694 495905 465762 495961
rect 465818 495905 465888 495961
rect 465568 495888 465888 495905
rect 496288 496333 496608 496350
rect 496288 496277 496358 496333
rect 496414 496277 496482 496333
rect 496538 496277 496608 496333
rect 496288 496209 496608 496277
rect 496288 496153 496358 496209
rect 496414 496153 496482 496209
rect 496538 496153 496608 496209
rect 496288 496085 496608 496153
rect 496288 496029 496358 496085
rect 496414 496029 496482 496085
rect 496538 496029 496608 496085
rect 496288 495961 496608 496029
rect 496288 495905 496358 495961
rect 496414 495905 496482 495961
rect 496538 495905 496608 495961
rect 496288 495888 496608 495905
rect 201154 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 201774 490350
rect 201154 490226 201774 490294
rect 201154 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 201774 490226
rect 201154 490102 201774 490170
rect 201154 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 201774 490102
rect 201154 489978 201774 490046
rect 201154 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 201774 489978
rect 201154 472350 201774 489922
rect 204448 490350 204768 490384
rect 204448 490294 204518 490350
rect 204574 490294 204642 490350
rect 204698 490294 204768 490350
rect 204448 490226 204768 490294
rect 204448 490170 204518 490226
rect 204574 490170 204642 490226
rect 204698 490170 204768 490226
rect 204448 490102 204768 490170
rect 204448 490046 204518 490102
rect 204574 490046 204642 490102
rect 204698 490046 204768 490102
rect 204448 489978 204768 490046
rect 204448 489922 204518 489978
rect 204574 489922 204642 489978
rect 204698 489922 204768 489978
rect 204448 489888 204768 489922
rect 235168 490350 235488 490384
rect 235168 490294 235238 490350
rect 235294 490294 235362 490350
rect 235418 490294 235488 490350
rect 235168 490226 235488 490294
rect 235168 490170 235238 490226
rect 235294 490170 235362 490226
rect 235418 490170 235488 490226
rect 235168 490102 235488 490170
rect 235168 490046 235238 490102
rect 235294 490046 235362 490102
rect 235418 490046 235488 490102
rect 235168 489978 235488 490046
rect 235168 489922 235238 489978
rect 235294 489922 235362 489978
rect 235418 489922 235488 489978
rect 235168 489888 235488 489922
rect 265888 490350 266208 490384
rect 265888 490294 265958 490350
rect 266014 490294 266082 490350
rect 266138 490294 266208 490350
rect 265888 490226 266208 490294
rect 265888 490170 265958 490226
rect 266014 490170 266082 490226
rect 266138 490170 266208 490226
rect 265888 490102 266208 490170
rect 265888 490046 265958 490102
rect 266014 490046 266082 490102
rect 266138 490046 266208 490102
rect 265888 489978 266208 490046
rect 265888 489922 265958 489978
rect 266014 489922 266082 489978
rect 266138 489922 266208 489978
rect 265888 489888 266208 489922
rect 296608 490350 296928 490384
rect 296608 490294 296678 490350
rect 296734 490294 296802 490350
rect 296858 490294 296928 490350
rect 296608 490226 296928 490294
rect 296608 490170 296678 490226
rect 296734 490170 296802 490226
rect 296858 490170 296928 490226
rect 296608 490102 296928 490170
rect 296608 490046 296678 490102
rect 296734 490046 296802 490102
rect 296858 490046 296928 490102
rect 296608 489978 296928 490046
rect 296608 489922 296678 489978
rect 296734 489922 296802 489978
rect 296858 489922 296928 489978
rect 296608 489888 296928 489922
rect 327328 490350 327648 490384
rect 327328 490294 327398 490350
rect 327454 490294 327522 490350
rect 327578 490294 327648 490350
rect 327328 490226 327648 490294
rect 327328 490170 327398 490226
rect 327454 490170 327522 490226
rect 327578 490170 327648 490226
rect 327328 490102 327648 490170
rect 327328 490046 327398 490102
rect 327454 490046 327522 490102
rect 327578 490046 327648 490102
rect 327328 489978 327648 490046
rect 327328 489922 327398 489978
rect 327454 489922 327522 489978
rect 327578 489922 327648 489978
rect 327328 489888 327648 489922
rect 358048 490350 358368 490384
rect 358048 490294 358118 490350
rect 358174 490294 358242 490350
rect 358298 490294 358368 490350
rect 358048 490226 358368 490294
rect 358048 490170 358118 490226
rect 358174 490170 358242 490226
rect 358298 490170 358368 490226
rect 358048 490102 358368 490170
rect 358048 490046 358118 490102
rect 358174 490046 358242 490102
rect 358298 490046 358368 490102
rect 358048 489978 358368 490046
rect 358048 489922 358118 489978
rect 358174 489922 358242 489978
rect 358298 489922 358368 489978
rect 358048 489888 358368 489922
rect 388768 490350 389088 490384
rect 388768 490294 388838 490350
rect 388894 490294 388962 490350
rect 389018 490294 389088 490350
rect 388768 490226 389088 490294
rect 388768 490170 388838 490226
rect 388894 490170 388962 490226
rect 389018 490170 389088 490226
rect 388768 490102 389088 490170
rect 388768 490046 388838 490102
rect 388894 490046 388962 490102
rect 389018 490046 389088 490102
rect 388768 489978 389088 490046
rect 388768 489922 388838 489978
rect 388894 489922 388962 489978
rect 389018 489922 389088 489978
rect 388768 489888 389088 489922
rect 419488 490350 419808 490384
rect 419488 490294 419558 490350
rect 419614 490294 419682 490350
rect 419738 490294 419808 490350
rect 419488 490226 419808 490294
rect 419488 490170 419558 490226
rect 419614 490170 419682 490226
rect 419738 490170 419808 490226
rect 419488 490102 419808 490170
rect 419488 490046 419558 490102
rect 419614 490046 419682 490102
rect 419738 490046 419808 490102
rect 419488 489978 419808 490046
rect 419488 489922 419558 489978
rect 419614 489922 419682 489978
rect 419738 489922 419808 489978
rect 419488 489888 419808 489922
rect 450208 490350 450528 490384
rect 450208 490294 450278 490350
rect 450334 490294 450402 490350
rect 450458 490294 450528 490350
rect 450208 490226 450528 490294
rect 450208 490170 450278 490226
rect 450334 490170 450402 490226
rect 450458 490170 450528 490226
rect 450208 490102 450528 490170
rect 450208 490046 450278 490102
rect 450334 490046 450402 490102
rect 450458 490046 450528 490102
rect 450208 489978 450528 490046
rect 450208 489922 450278 489978
rect 450334 489922 450402 489978
rect 450458 489922 450528 489978
rect 450208 489888 450528 489922
rect 480928 490350 481248 490384
rect 480928 490294 480998 490350
rect 481054 490294 481122 490350
rect 481178 490294 481248 490350
rect 480928 490226 481248 490294
rect 480928 490170 480998 490226
rect 481054 490170 481122 490226
rect 481178 490170 481248 490226
rect 480928 490102 481248 490170
rect 480928 490046 480998 490102
rect 481054 490046 481122 490102
rect 481178 490046 481248 490102
rect 480928 489978 481248 490046
rect 480928 489922 480998 489978
rect 481054 489922 481122 489978
rect 481178 489922 481248 489978
rect 480928 489888 481248 489922
rect 507154 490350 507774 507922
rect 507154 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 507774 490350
rect 507154 490226 507774 490294
rect 507154 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 507774 490226
rect 507154 490102 507774 490170
rect 507154 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 507774 490102
rect 507154 489978 507774 490046
rect 507154 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 507774 489978
rect 219808 478350 220128 478384
rect 219808 478294 219878 478350
rect 219934 478294 220002 478350
rect 220058 478294 220128 478350
rect 219808 478226 220128 478294
rect 219808 478170 219878 478226
rect 219934 478170 220002 478226
rect 220058 478170 220128 478226
rect 219808 478102 220128 478170
rect 219808 478046 219878 478102
rect 219934 478046 220002 478102
rect 220058 478046 220128 478102
rect 219808 477978 220128 478046
rect 219808 477922 219878 477978
rect 219934 477922 220002 477978
rect 220058 477922 220128 477978
rect 219808 477888 220128 477922
rect 250528 478350 250848 478384
rect 250528 478294 250598 478350
rect 250654 478294 250722 478350
rect 250778 478294 250848 478350
rect 250528 478226 250848 478294
rect 250528 478170 250598 478226
rect 250654 478170 250722 478226
rect 250778 478170 250848 478226
rect 250528 478102 250848 478170
rect 250528 478046 250598 478102
rect 250654 478046 250722 478102
rect 250778 478046 250848 478102
rect 250528 477978 250848 478046
rect 250528 477922 250598 477978
rect 250654 477922 250722 477978
rect 250778 477922 250848 477978
rect 250528 477888 250848 477922
rect 281248 478350 281568 478384
rect 281248 478294 281318 478350
rect 281374 478294 281442 478350
rect 281498 478294 281568 478350
rect 281248 478226 281568 478294
rect 281248 478170 281318 478226
rect 281374 478170 281442 478226
rect 281498 478170 281568 478226
rect 281248 478102 281568 478170
rect 281248 478046 281318 478102
rect 281374 478046 281442 478102
rect 281498 478046 281568 478102
rect 281248 477978 281568 478046
rect 281248 477922 281318 477978
rect 281374 477922 281442 477978
rect 281498 477922 281568 477978
rect 281248 477888 281568 477922
rect 311968 478350 312288 478384
rect 311968 478294 312038 478350
rect 312094 478294 312162 478350
rect 312218 478294 312288 478350
rect 311968 478226 312288 478294
rect 311968 478170 312038 478226
rect 312094 478170 312162 478226
rect 312218 478170 312288 478226
rect 311968 478102 312288 478170
rect 311968 478046 312038 478102
rect 312094 478046 312162 478102
rect 312218 478046 312288 478102
rect 311968 477978 312288 478046
rect 311968 477922 312038 477978
rect 312094 477922 312162 477978
rect 312218 477922 312288 477978
rect 311968 477888 312288 477922
rect 342688 478350 343008 478384
rect 342688 478294 342758 478350
rect 342814 478294 342882 478350
rect 342938 478294 343008 478350
rect 342688 478226 343008 478294
rect 342688 478170 342758 478226
rect 342814 478170 342882 478226
rect 342938 478170 343008 478226
rect 342688 478102 343008 478170
rect 342688 478046 342758 478102
rect 342814 478046 342882 478102
rect 342938 478046 343008 478102
rect 342688 477978 343008 478046
rect 342688 477922 342758 477978
rect 342814 477922 342882 477978
rect 342938 477922 343008 477978
rect 342688 477888 343008 477922
rect 373408 478350 373728 478384
rect 373408 478294 373478 478350
rect 373534 478294 373602 478350
rect 373658 478294 373728 478350
rect 373408 478226 373728 478294
rect 373408 478170 373478 478226
rect 373534 478170 373602 478226
rect 373658 478170 373728 478226
rect 373408 478102 373728 478170
rect 373408 478046 373478 478102
rect 373534 478046 373602 478102
rect 373658 478046 373728 478102
rect 373408 477978 373728 478046
rect 373408 477922 373478 477978
rect 373534 477922 373602 477978
rect 373658 477922 373728 477978
rect 373408 477888 373728 477922
rect 404128 478350 404448 478384
rect 404128 478294 404198 478350
rect 404254 478294 404322 478350
rect 404378 478294 404448 478350
rect 404128 478226 404448 478294
rect 404128 478170 404198 478226
rect 404254 478170 404322 478226
rect 404378 478170 404448 478226
rect 404128 478102 404448 478170
rect 404128 478046 404198 478102
rect 404254 478046 404322 478102
rect 404378 478046 404448 478102
rect 404128 477978 404448 478046
rect 404128 477922 404198 477978
rect 404254 477922 404322 477978
rect 404378 477922 404448 477978
rect 404128 477888 404448 477922
rect 434848 478350 435168 478384
rect 434848 478294 434918 478350
rect 434974 478294 435042 478350
rect 435098 478294 435168 478350
rect 434848 478226 435168 478294
rect 434848 478170 434918 478226
rect 434974 478170 435042 478226
rect 435098 478170 435168 478226
rect 434848 478102 435168 478170
rect 434848 478046 434918 478102
rect 434974 478046 435042 478102
rect 435098 478046 435168 478102
rect 434848 477978 435168 478046
rect 434848 477922 434918 477978
rect 434974 477922 435042 477978
rect 435098 477922 435168 477978
rect 434848 477888 435168 477922
rect 465568 478350 465888 478384
rect 465568 478294 465638 478350
rect 465694 478294 465762 478350
rect 465818 478294 465888 478350
rect 465568 478226 465888 478294
rect 465568 478170 465638 478226
rect 465694 478170 465762 478226
rect 465818 478170 465888 478226
rect 465568 478102 465888 478170
rect 465568 478046 465638 478102
rect 465694 478046 465762 478102
rect 465818 478046 465888 478102
rect 465568 477978 465888 478046
rect 465568 477922 465638 477978
rect 465694 477922 465762 477978
rect 465818 477922 465888 477978
rect 465568 477888 465888 477922
rect 496288 478350 496608 478384
rect 496288 478294 496358 478350
rect 496414 478294 496482 478350
rect 496538 478294 496608 478350
rect 496288 478226 496608 478294
rect 496288 478170 496358 478226
rect 496414 478170 496482 478226
rect 496538 478170 496608 478226
rect 496288 478102 496608 478170
rect 496288 478046 496358 478102
rect 496414 478046 496482 478102
rect 496538 478046 496608 478102
rect 496288 477978 496608 478046
rect 496288 477922 496358 477978
rect 496414 477922 496482 477978
rect 496538 477922 496608 477978
rect 496288 477888 496608 477922
rect 201154 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 201774 472350
rect 201154 472226 201774 472294
rect 201154 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 201774 472226
rect 201154 472102 201774 472170
rect 201154 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 201774 472102
rect 201154 471978 201774 472046
rect 201154 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 201774 471978
rect 201154 454350 201774 471922
rect 204448 472350 204768 472384
rect 204448 472294 204518 472350
rect 204574 472294 204642 472350
rect 204698 472294 204768 472350
rect 204448 472226 204768 472294
rect 204448 472170 204518 472226
rect 204574 472170 204642 472226
rect 204698 472170 204768 472226
rect 204448 472102 204768 472170
rect 204448 472046 204518 472102
rect 204574 472046 204642 472102
rect 204698 472046 204768 472102
rect 204448 471978 204768 472046
rect 204448 471922 204518 471978
rect 204574 471922 204642 471978
rect 204698 471922 204768 471978
rect 204448 471888 204768 471922
rect 235168 472350 235488 472384
rect 235168 472294 235238 472350
rect 235294 472294 235362 472350
rect 235418 472294 235488 472350
rect 235168 472226 235488 472294
rect 235168 472170 235238 472226
rect 235294 472170 235362 472226
rect 235418 472170 235488 472226
rect 235168 472102 235488 472170
rect 235168 472046 235238 472102
rect 235294 472046 235362 472102
rect 235418 472046 235488 472102
rect 235168 471978 235488 472046
rect 235168 471922 235238 471978
rect 235294 471922 235362 471978
rect 235418 471922 235488 471978
rect 235168 471888 235488 471922
rect 265888 472350 266208 472384
rect 265888 472294 265958 472350
rect 266014 472294 266082 472350
rect 266138 472294 266208 472350
rect 265888 472226 266208 472294
rect 265888 472170 265958 472226
rect 266014 472170 266082 472226
rect 266138 472170 266208 472226
rect 265888 472102 266208 472170
rect 265888 472046 265958 472102
rect 266014 472046 266082 472102
rect 266138 472046 266208 472102
rect 265888 471978 266208 472046
rect 265888 471922 265958 471978
rect 266014 471922 266082 471978
rect 266138 471922 266208 471978
rect 265888 471888 266208 471922
rect 296608 472350 296928 472384
rect 296608 472294 296678 472350
rect 296734 472294 296802 472350
rect 296858 472294 296928 472350
rect 296608 472226 296928 472294
rect 296608 472170 296678 472226
rect 296734 472170 296802 472226
rect 296858 472170 296928 472226
rect 296608 472102 296928 472170
rect 296608 472046 296678 472102
rect 296734 472046 296802 472102
rect 296858 472046 296928 472102
rect 296608 471978 296928 472046
rect 296608 471922 296678 471978
rect 296734 471922 296802 471978
rect 296858 471922 296928 471978
rect 296608 471888 296928 471922
rect 327328 472350 327648 472384
rect 327328 472294 327398 472350
rect 327454 472294 327522 472350
rect 327578 472294 327648 472350
rect 327328 472226 327648 472294
rect 327328 472170 327398 472226
rect 327454 472170 327522 472226
rect 327578 472170 327648 472226
rect 327328 472102 327648 472170
rect 327328 472046 327398 472102
rect 327454 472046 327522 472102
rect 327578 472046 327648 472102
rect 327328 471978 327648 472046
rect 327328 471922 327398 471978
rect 327454 471922 327522 471978
rect 327578 471922 327648 471978
rect 327328 471888 327648 471922
rect 358048 472350 358368 472384
rect 358048 472294 358118 472350
rect 358174 472294 358242 472350
rect 358298 472294 358368 472350
rect 358048 472226 358368 472294
rect 358048 472170 358118 472226
rect 358174 472170 358242 472226
rect 358298 472170 358368 472226
rect 358048 472102 358368 472170
rect 358048 472046 358118 472102
rect 358174 472046 358242 472102
rect 358298 472046 358368 472102
rect 358048 471978 358368 472046
rect 358048 471922 358118 471978
rect 358174 471922 358242 471978
rect 358298 471922 358368 471978
rect 358048 471888 358368 471922
rect 388768 472350 389088 472384
rect 388768 472294 388838 472350
rect 388894 472294 388962 472350
rect 389018 472294 389088 472350
rect 388768 472226 389088 472294
rect 388768 472170 388838 472226
rect 388894 472170 388962 472226
rect 389018 472170 389088 472226
rect 388768 472102 389088 472170
rect 388768 472046 388838 472102
rect 388894 472046 388962 472102
rect 389018 472046 389088 472102
rect 388768 471978 389088 472046
rect 388768 471922 388838 471978
rect 388894 471922 388962 471978
rect 389018 471922 389088 471978
rect 388768 471888 389088 471922
rect 419488 472350 419808 472384
rect 419488 472294 419558 472350
rect 419614 472294 419682 472350
rect 419738 472294 419808 472350
rect 419488 472226 419808 472294
rect 419488 472170 419558 472226
rect 419614 472170 419682 472226
rect 419738 472170 419808 472226
rect 419488 472102 419808 472170
rect 419488 472046 419558 472102
rect 419614 472046 419682 472102
rect 419738 472046 419808 472102
rect 419488 471978 419808 472046
rect 419488 471922 419558 471978
rect 419614 471922 419682 471978
rect 419738 471922 419808 471978
rect 419488 471888 419808 471922
rect 450208 472350 450528 472384
rect 450208 472294 450278 472350
rect 450334 472294 450402 472350
rect 450458 472294 450528 472350
rect 450208 472226 450528 472294
rect 450208 472170 450278 472226
rect 450334 472170 450402 472226
rect 450458 472170 450528 472226
rect 450208 472102 450528 472170
rect 450208 472046 450278 472102
rect 450334 472046 450402 472102
rect 450458 472046 450528 472102
rect 450208 471978 450528 472046
rect 450208 471922 450278 471978
rect 450334 471922 450402 471978
rect 450458 471922 450528 471978
rect 450208 471888 450528 471922
rect 480928 472350 481248 472384
rect 480928 472294 480998 472350
rect 481054 472294 481122 472350
rect 481178 472294 481248 472350
rect 480928 472226 481248 472294
rect 480928 472170 480998 472226
rect 481054 472170 481122 472226
rect 481178 472170 481248 472226
rect 480928 472102 481248 472170
rect 480928 472046 480998 472102
rect 481054 472046 481122 472102
rect 481178 472046 481248 472102
rect 480928 471978 481248 472046
rect 480928 471922 480998 471978
rect 481054 471922 481122 471978
rect 481178 471922 481248 471978
rect 480928 471888 481248 471922
rect 507154 472350 507774 489922
rect 507154 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 507774 472350
rect 507154 472226 507774 472294
rect 507154 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 507774 472226
rect 507154 472102 507774 472170
rect 507154 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 507774 472102
rect 507154 471978 507774 472046
rect 507154 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 507774 471978
rect 219808 460350 220128 460384
rect 219808 460294 219878 460350
rect 219934 460294 220002 460350
rect 220058 460294 220128 460350
rect 219808 460226 220128 460294
rect 219808 460170 219878 460226
rect 219934 460170 220002 460226
rect 220058 460170 220128 460226
rect 219808 460102 220128 460170
rect 219808 460046 219878 460102
rect 219934 460046 220002 460102
rect 220058 460046 220128 460102
rect 219808 459978 220128 460046
rect 219808 459922 219878 459978
rect 219934 459922 220002 459978
rect 220058 459922 220128 459978
rect 219808 459888 220128 459922
rect 250528 460350 250848 460384
rect 250528 460294 250598 460350
rect 250654 460294 250722 460350
rect 250778 460294 250848 460350
rect 250528 460226 250848 460294
rect 250528 460170 250598 460226
rect 250654 460170 250722 460226
rect 250778 460170 250848 460226
rect 250528 460102 250848 460170
rect 250528 460046 250598 460102
rect 250654 460046 250722 460102
rect 250778 460046 250848 460102
rect 250528 459978 250848 460046
rect 250528 459922 250598 459978
rect 250654 459922 250722 459978
rect 250778 459922 250848 459978
rect 250528 459888 250848 459922
rect 281248 460350 281568 460384
rect 281248 460294 281318 460350
rect 281374 460294 281442 460350
rect 281498 460294 281568 460350
rect 281248 460226 281568 460294
rect 281248 460170 281318 460226
rect 281374 460170 281442 460226
rect 281498 460170 281568 460226
rect 281248 460102 281568 460170
rect 281248 460046 281318 460102
rect 281374 460046 281442 460102
rect 281498 460046 281568 460102
rect 281248 459978 281568 460046
rect 281248 459922 281318 459978
rect 281374 459922 281442 459978
rect 281498 459922 281568 459978
rect 281248 459888 281568 459922
rect 311968 460350 312288 460384
rect 311968 460294 312038 460350
rect 312094 460294 312162 460350
rect 312218 460294 312288 460350
rect 311968 460226 312288 460294
rect 311968 460170 312038 460226
rect 312094 460170 312162 460226
rect 312218 460170 312288 460226
rect 311968 460102 312288 460170
rect 311968 460046 312038 460102
rect 312094 460046 312162 460102
rect 312218 460046 312288 460102
rect 311968 459978 312288 460046
rect 311968 459922 312038 459978
rect 312094 459922 312162 459978
rect 312218 459922 312288 459978
rect 311968 459888 312288 459922
rect 342688 460350 343008 460384
rect 342688 460294 342758 460350
rect 342814 460294 342882 460350
rect 342938 460294 343008 460350
rect 342688 460226 343008 460294
rect 342688 460170 342758 460226
rect 342814 460170 342882 460226
rect 342938 460170 343008 460226
rect 342688 460102 343008 460170
rect 342688 460046 342758 460102
rect 342814 460046 342882 460102
rect 342938 460046 343008 460102
rect 342688 459978 343008 460046
rect 342688 459922 342758 459978
rect 342814 459922 342882 459978
rect 342938 459922 343008 459978
rect 342688 459888 343008 459922
rect 373408 460350 373728 460384
rect 373408 460294 373478 460350
rect 373534 460294 373602 460350
rect 373658 460294 373728 460350
rect 373408 460226 373728 460294
rect 373408 460170 373478 460226
rect 373534 460170 373602 460226
rect 373658 460170 373728 460226
rect 373408 460102 373728 460170
rect 373408 460046 373478 460102
rect 373534 460046 373602 460102
rect 373658 460046 373728 460102
rect 373408 459978 373728 460046
rect 373408 459922 373478 459978
rect 373534 459922 373602 459978
rect 373658 459922 373728 459978
rect 373408 459888 373728 459922
rect 404128 460350 404448 460384
rect 404128 460294 404198 460350
rect 404254 460294 404322 460350
rect 404378 460294 404448 460350
rect 404128 460226 404448 460294
rect 404128 460170 404198 460226
rect 404254 460170 404322 460226
rect 404378 460170 404448 460226
rect 404128 460102 404448 460170
rect 404128 460046 404198 460102
rect 404254 460046 404322 460102
rect 404378 460046 404448 460102
rect 404128 459978 404448 460046
rect 404128 459922 404198 459978
rect 404254 459922 404322 459978
rect 404378 459922 404448 459978
rect 404128 459888 404448 459922
rect 434848 460350 435168 460384
rect 434848 460294 434918 460350
rect 434974 460294 435042 460350
rect 435098 460294 435168 460350
rect 434848 460226 435168 460294
rect 434848 460170 434918 460226
rect 434974 460170 435042 460226
rect 435098 460170 435168 460226
rect 434848 460102 435168 460170
rect 434848 460046 434918 460102
rect 434974 460046 435042 460102
rect 435098 460046 435168 460102
rect 434848 459978 435168 460046
rect 434848 459922 434918 459978
rect 434974 459922 435042 459978
rect 435098 459922 435168 459978
rect 434848 459888 435168 459922
rect 465568 460350 465888 460384
rect 465568 460294 465638 460350
rect 465694 460294 465762 460350
rect 465818 460294 465888 460350
rect 465568 460226 465888 460294
rect 465568 460170 465638 460226
rect 465694 460170 465762 460226
rect 465818 460170 465888 460226
rect 465568 460102 465888 460170
rect 465568 460046 465638 460102
rect 465694 460046 465762 460102
rect 465818 460046 465888 460102
rect 465568 459978 465888 460046
rect 465568 459922 465638 459978
rect 465694 459922 465762 459978
rect 465818 459922 465888 459978
rect 465568 459888 465888 459922
rect 496288 460350 496608 460384
rect 496288 460294 496358 460350
rect 496414 460294 496482 460350
rect 496538 460294 496608 460350
rect 496288 460226 496608 460294
rect 496288 460170 496358 460226
rect 496414 460170 496482 460226
rect 496538 460170 496608 460226
rect 496288 460102 496608 460170
rect 496288 460046 496358 460102
rect 496414 460046 496482 460102
rect 496538 460046 496608 460102
rect 496288 459978 496608 460046
rect 496288 459922 496358 459978
rect 496414 459922 496482 459978
rect 496538 459922 496608 459978
rect 496288 459888 496608 459922
rect 201154 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 201774 454350
rect 201154 454226 201774 454294
rect 201154 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 201774 454226
rect 201154 454102 201774 454170
rect 201154 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 201774 454102
rect 201154 453978 201774 454046
rect 201154 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 201774 453978
rect 201154 436350 201774 453922
rect 204448 454350 204768 454384
rect 204448 454294 204518 454350
rect 204574 454294 204642 454350
rect 204698 454294 204768 454350
rect 204448 454226 204768 454294
rect 204448 454170 204518 454226
rect 204574 454170 204642 454226
rect 204698 454170 204768 454226
rect 204448 454102 204768 454170
rect 204448 454046 204518 454102
rect 204574 454046 204642 454102
rect 204698 454046 204768 454102
rect 204448 453978 204768 454046
rect 204448 453922 204518 453978
rect 204574 453922 204642 453978
rect 204698 453922 204768 453978
rect 204448 453888 204768 453922
rect 235168 454350 235488 454384
rect 235168 454294 235238 454350
rect 235294 454294 235362 454350
rect 235418 454294 235488 454350
rect 235168 454226 235488 454294
rect 235168 454170 235238 454226
rect 235294 454170 235362 454226
rect 235418 454170 235488 454226
rect 235168 454102 235488 454170
rect 235168 454046 235238 454102
rect 235294 454046 235362 454102
rect 235418 454046 235488 454102
rect 235168 453978 235488 454046
rect 235168 453922 235238 453978
rect 235294 453922 235362 453978
rect 235418 453922 235488 453978
rect 235168 453888 235488 453922
rect 265888 454350 266208 454384
rect 265888 454294 265958 454350
rect 266014 454294 266082 454350
rect 266138 454294 266208 454350
rect 265888 454226 266208 454294
rect 265888 454170 265958 454226
rect 266014 454170 266082 454226
rect 266138 454170 266208 454226
rect 265888 454102 266208 454170
rect 265888 454046 265958 454102
rect 266014 454046 266082 454102
rect 266138 454046 266208 454102
rect 265888 453978 266208 454046
rect 265888 453922 265958 453978
rect 266014 453922 266082 453978
rect 266138 453922 266208 453978
rect 265888 453888 266208 453922
rect 296608 454350 296928 454384
rect 296608 454294 296678 454350
rect 296734 454294 296802 454350
rect 296858 454294 296928 454350
rect 296608 454226 296928 454294
rect 296608 454170 296678 454226
rect 296734 454170 296802 454226
rect 296858 454170 296928 454226
rect 296608 454102 296928 454170
rect 296608 454046 296678 454102
rect 296734 454046 296802 454102
rect 296858 454046 296928 454102
rect 296608 453978 296928 454046
rect 296608 453922 296678 453978
rect 296734 453922 296802 453978
rect 296858 453922 296928 453978
rect 296608 453888 296928 453922
rect 327328 454350 327648 454384
rect 327328 454294 327398 454350
rect 327454 454294 327522 454350
rect 327578 454294 327648 454350
rect 327328 454226 327648 454294
rect 327328 454170 327398 454226
rect 327454 454170 327522 454226
rect 327578 454170 327648 454226
rect 327328 454102 327648 454170
rect 327328 454046 327398 454102
rect 327454 454046 327522 454102
rect 327578 454046 327648 454102
rect 327328 453978 327648 454046
rect 327328 453922 327398 453978
rect 327454 453922 327522 453978
rect 327578 453922 327648 453978
rect 327328 453888 327648 453922
rect 358048 454350 358368 454384
rect 358048 454294 358118 454350
rect 358174 454294 358242 454350
rect 358298 454294 358368 454350
rect 358048 454226 358368 454294
rect 358048 454170 358118 454226
rect 358174 454170 358242 454226
rect 358298 454170 358368 454226
rect 358048 454102 358368 454170
rect 358048 454046 358118 454102
rect 358174 454046 358242 454102
rect 358298 454046 358368 454102
rect 358048 453978 358368 454046
rect 358048 453922 358118 453978
rect 358174 453922 358242 453978
rect 358298 453922 358368 453978
rect 358048 453888 358368 453922
rect 388768 454350 389088 454384
rect 388768 454294 388838 454350
rect 388894 454294 388962 454350
rect 389018 454294 389088 454350
rect 388768 454226 389088 454294
rect 388768 454170 388838 454226
rect 388894 454170 388962 454226
rect 389018 454170 389088 454226
rect 388768 454102 389088 454170
rect 388768 454046 388838 454102
rect 388894 454046 388962 454102
rect 389018 454046 389088 454102
rect 388768 453978 389088 454046
rect 388768 453922 388838 453978
rect 388894 453922 388962 453978
rect 389018 453922 389088 453978
rect 388768 453888 389088 453922
rect 419488 454350 419808 454384
rect 419488 454294 419558 454350
rect 419614 454294 419682 454350
rect 419738 454294 419808 454350
rect 419488 454226 419808 454294
rect 419488 454170 419558 454226
rect 419614 454170 419682 454226
rect 419738 454170 419808 454226
rect 419488 454102 419808 454170
rect 419488 454046 419558 454102
rect 419614 454046 419682 454102
rect 419738 454046 419808 454102
rect 419488 453978 419808 454046
rect 419488 453922 419558 453978
rect 419614 453922 419682 453978
rect 419738 453922 419808 453978
rect 419488 453888 419808 453922
rect 450208 454350 450528 454384
rect 450208 454294 450278 454350
rect 450334 454294 450402 454350
rect 450458 454294 450528 454350
rect 450208 454226 450528 454294
rect 450208 454170 450278 454226
rect 450334 454170 450402 454226
rect 450458 454170 450528 454226
rect 450208 454102 450528 454170
rect 450208 454046 450278 454102
rect 450334 454046 450402 454102
rect 450458 454046 450528 454102
rect 450208 453978 450528 454046
rect 450208 453922 450278 453978
rect 450334 453922 450402 453978
rect 450458 453922 450528 453978
rect 450208 453888 450528 453922
rect 480928 454350 481248 454384
rect 480928 454294 480998 454350
rect 481054 454294 481122 454350
rect 481178 454294 481248 454350
rect 480928 454226 481248 454294
rect 480928 454170 480998 454226
rect 481054 454170 481122 454226
rect 481178 454170 481248 454226
rect 480928 454102 481248 454170
rect 480928 454046 480998 454102
rect 481054 454046 481122 454102
rect 481178 454046 481248 454102
rect 480928 453978 481248 454046
rect 480928 453922 480998 453978
rect 481054 453922 481122 453978
rect 481178 453922 481248 453978
rect 480928 453888 481248 453922
rect 507154 454350 507774 471922
rect 507154 454294 507250 454350
rect 507306 454294 507374 454350
rect 507430 454294 507498 454350
rect 507554 454294 507622 454350
rect 507678 454294 507774 454350
rect 507154 454226 507774 454294
rect 507154 454170 507250 454226
rect 507306 454170 507374 454226
rect 507430 454170 507498 454226
rect 507554 454170 507622 454226
rect 507678 454170 507774 454226
rect 507154 454102 507774 454170
rect 507154 454046 507250 454102
rect 507306 454046 507374 454102
rect 507430 454046 507498 454102
rect 507554 454046 507622 454102
rect 507678 454046 507774 454102
rect 507154 453978 507774 454046
rect 507154 453922 507250 453978
rect 507306 453922 507374 453978
rect 507430 453922 507498 453978
rect 507554 453922 507622 453978
rect 507678 453922 507774 453978
rect 219808 442350 220128 442384
rect 219808 442294 219878 442350
rect 219934 442294 220002 442350
rect 220058 442294 220128 442350
rect 219808 442226 220128 442294
rect 219808 442170 219878 442226
rect 219934 442170 220002 442226
rect 220058 442170 220128 442226
rect 219808 442102 220128 442170
rect 219808 442046 219878 442102
rect 219934 442046 220002 442102
rect 220058 442046 220128 442102
rect 219808 441978 220128 442046
rect 219808 441922 219878 441978
rect 219934 441922 220002 441978
rect 220058 441922 220128 441978
rect 219808 441888 220128 441922
rect 250528 442350 250848 442384
rect 250528 442294 250598 442350
rect 250654 442294 250722 442350
rect 250778 442294 250848 442350
rect 250528 442226 250848 442294
rect 250528 442170 250598 442226
rect 250654 442170 250722 442226
rect 250778 442170 250848 442226
rect 250528 442102 250848 442170
rect 250528 442046 250598 442102
rect 250654 442046 250722 442102
rect 250778 442046 250848 442102
rect 250528 441978 250848 442046
rect 250528 441922 250598 441978
rect 250654 441922 250722 441978
rect 250778 441922 250848 441978
rect 250528 441888 250848 441922
rect 281248 442350 281568 442384
rect 281248 442294 281318 442350
rect 281374 442294 281442 442350
rect 281498 442294 281568 442350
rect 281248 442226 281568 442294
rect 281248 442170 281318 442226
rect 281374 442170 281442 442226
rect 281498 442170 281568 442226
rect 281248 442102 281568 442170
rect 281248 442046 281318 442102
rect 281374 442046 281442 442102
rect 281498 442046 281568 442102
rect 281248 441978 281568 442046
rect 281248 441922 281318 441978
rect 281374 441922 281442 441978
rect 281498 441922 281568 441978
rect 281248 441888 281568 441922
rect 311968 442350 312288 442384
rect 311968 442294 312038 442350
rect 312094 442294 312162 442350
rect 312218 442294 312288 442350
rect 311968 442226 312288 442294
rect 311968 442170 312038 442226
rect 312094 442170 312162 442226
rect 312218 442170 312288 442226
rect 311968 442102 312288 442170
rect 311968 442046 312038 442102
rect 312094 442046 312162 442102
rect 312218 442046 312288 442102
rect 311968 441978 312288 442046
rect 311968 441922 312038 441978
rect 312094 441922 312162 441978
rect 312218 441922 312288 441978
rect 311968 441888 312288 441922
rect 342688 442350 343008 442384
rect 342688 442294 342758 442350
rect 342814 442294 342882 442350
rect 342938 442294 343008 442350
rect 342688 442226 343008 442294
rect 342688 442170 342758 442226
rect 342814 442170 342882 442226
rect 342938 442170 343008 442226
rect 342688 442102 343008 442170
rect 342688 442046 342758 442102
rect 342814 442046 342882 442102
rect 342938 442046 343008 442102
rect 342688 441978 343008 442046
rect 342688 441922 342758 441978
rect 342814 441922 342882 441978
rect 342938 441922 343008 441978
rect 342688 441888 343008 441922
rect 373408 442350 373728 442384
rect 373408 442294 373478 442350
rect 373534 442294 373602 442350
rect 373658 442294 373728 442350
rect 373408 442226 373728 442294
rect 373408 442170 373478 442226
rect 373534 442170 373602 442226
rect 373658 442170 373728 442226
rect 373408 442102 373728 442170
rect 373408 442046 373478 442102
rect 373534 442046 373602 442102
rect 373658 442046 373728 442102
rect 373408 441978 373728 442046
rect 373408 441922 373478 441978
rect 373534 441922 373602 441978
rect 373658 441922 373728 441978
rect 373408 441888 373728 441922
rect 404128 442350 404448 442384
rect 404128 442294 404198 442350
rect 404254 442294 404322 442350
rect 404378 442294 404448 442350
rect 404128 442226 404448 442294
rect 404128 442170 404198 442226
rect 404254 442170 404322 442226
rect 404378 442170 404448 442226
rect 404128 442102 404448 442170
rect 404128 442046 404198 442102
rect 404254 442046 404322 442102
rect 404378 442046 404448 442102
rect 404128 441978 404448 442046
rect 404128 441922 404198 441978
rect 404254 441922 404322 441978
rect 404378 441922 404448 441978
rect 404128 441888 404448 441922
rect 434848 442350 435168 442384
rect 434848 442294 434918 442350
rect 434974 442294 435042 442350
rect 435098 442294 435168 442350
rect 434848 442226 435168 442294
rect 434848 442170 434918 442226
rect 434974 442170 435042 442226
rect 435098 442170 435168 442226
rect 434848 442102 435168 442170
rect 434848 442046 434918 442102
rect 434974 442046 435042 442102
rect 435098 442046 435168 442102
rect 434848 441978 435168 442046
rect 434848 441922 434918 441978
rect 434974 441922 435042 441978
rect 435098 441922 435168 441978
rect 434848 441888 435168 441922
rect 465568 442350 465888 442384
rect 465568 442294 465638 442350
rect 465694 442294 465762 442350
rect 465818 442294 465888 442350
rect 465568 442226 465888 442294
rect 465568 442170 465638 442226
rect 465694 442170 465762 442226
rect 465818 442170 465888 442226
rect 465568 442102 465888 442170
rect 465568 442046 465638 442102
rect 465694 442046 465762 442102
rect 465818 442046 465888 442102
rect 465568 441978 465888 442046
rect 465568 441922 465638 441978
rect 465694 441922 465762 441978
rect 465818 441922 465888 441978
rect 465568 441888 465888 441922
rect 496288 442350 496608 442384
rect 496288 442294 496358 442350
rect 496414 442294 496482 442350
rect 496538 442294 496608 442350
rect 496288 442226 496608 442294
rect 496288 442170 496358 442226
rect 496414 442170 496482 442226
rect 496538 442170 496608 442226
rect 496288 442102 496608 442170
rect 496288 442046 496358 442102
rect 496414 442046 496482 442102
rect 496538 442046 496608 442102
rect 496288 441978 496608 442046
rect 496288 441922 496358 441978
rect 496414 441922 496482 441978
rect 496538 441922 496608 441978
rect 496288 441888 496608 441922
rect 201154 436294 201250 436350
rect 201306 436294 201374 436350
rect 201430 436294 201498 436350
rect 201554 436294 201622 436350
rect 201678 436294 201774 436350
rect 201154 436226 201774 436294
rect 201154 436170 201250 436226
rect 201306 436170 201374 436226
rect 201430 436170 201498 436226
rect 201554 436170 201622 436226
rect 201678 436170 201774 436226
rect 201154 436102 201774 436170
rect 201154 436046 201250 436102
rect 201306 436046 201374 436102
rect 201430 436046 201498 436102
rect 201554 436046 201622 436102
rect 201678 436046 201774 436102
rect 201154 435978 201774 436046
rect 201154 435922 201250 435978
rect 201306 435922 201374 435978
rect 201430 435922 201498 435978
rect 201554 435922 201622 435978
rect 201678 435922 201774 435978
rect 201154 418350 201774 435922
rect 204448 436350 204768 436384
rect 204448 436294 204518 436350
rect 204574 436294 204642 436350
rect 204698 436294 204768 436350
rect 204448 436226 204768 436294
rect 204448 436170 204518 436226
rect 204574 436170 204642 436226
rect 204698 436170 204768 436226
rect 204448 436102 204768 436170
rect 204448 436046 204518 436102
rect 204574 436046 204642 436102
rect 204698 436046 204768 436102
rect 204448 435978 204768 436046
rect 204448 435922 204518 435978
rect 204574 435922 204642 435978
rect 204698 435922 204768 435978
rect 204448 435888 204768 435922
rect 235168 436350 235488 436384
rect 235168 436294 235238 436350
rect 235294 436294 235362 436350
rect 235418 436294 235488 436350
rect 235168 436226 235488 436294
rect 235168 436170 235238 436226
rect 235294 436170 235362 436226
rect 235418 436170 235488 436226
rect 235168 436102 235488 436170
rect 235168 436046 235238 436102
rect 235294 436046 235362 436102
rect 235418 436046 235488 436102
rect 235168 435978 235488 436046
rect 235168 435922 235238 435978
rect 235294 435922 235362 435978
rect 235418 435922 235488 435978
rect 235168 435888 235488 435922
rect 265888 436350 266208 436384
rect 265888 436294 265958 436350
rect 266014 436294 266082 436350
rect 266138 436294 266208 436350
rect 265888 436226 266208 436294
rect 265888 436170 265958 436226
rect 266014 436170 266082 436226
rect 266138 436170 266208 436226
rect 265888 436102 266208 436170
rect 265888 436046 265958 436102
rect 266014 436046 266082 436102
rect 266138 436046 266208 436102
rect 265888 435978 266208 436046
rect 265888 435922 265958 435978
rect 266014 435922 266082 435978
rect 266138 435922 266208 435978
rect 265888 435888 266208 435922
rect 296608 436350 296928 436384
rect 296608 436294 296678 436350
rect 296734 436294 296802 436350
rect 296858 436294 296928 436350
rect 296608 436226 296928 436294
rect 296608 436170 296678 436226
rect 296734 436170 296802 436226
rect 296858 436170 296928 436226
rect 296608 436102 296928 436170
rect 296608 436046 296678 436102
rect 296734 436046 296802 436102
rect 296858 436046 296928 436102
rect 296608 435978 296928 436046
rect 296608 435922 296678 435978
rect 296734 435922 296802 435978
rect 296858 435922 296928 435978
rect 296608 435888 296928 435922
rect 327328 436350 327648 436384
rect 327328 436294 327398 436350
rect 327454 436294 327522 436350
rect 327578 436294 327648 436350
rect 327328 436226 327648 436294
rect 327328 436170 327398 436226
rect 327454 436170 327522 436226
rect 327578 436170 327648 436226
rect 327328 436102 327648 436170
rect 327328 436046 327398 436102
rect 327454 436046 327522 436102
rect 327578 436046 327648 436102
rect 327328 435978 327648 436046
rect 327328 435922 327398 435978
rect 327454 435922 327522 435978
rect 327578 435922 327648 435978
rect 327328 435888 327648 435922
rect 358048 436350 358368 436384
rect 358048 436294 358118 436350
rect 358174 436294 358242 436350
rect 358298 436294 358368 436350
rect 358048 436226 358368 436294
rect 358048 436170 358118 436226
rect 358174 436170 358242 436226
rect 358298 436170 358368 436226
rect 358048 436102 358368 436170
rect 358048 436046 358118 436102
rect 358174 436046 358242 436102
rect 358298 436046 358368 436102
rect 358048 435978 358368 436046
rect 358048 435922 358118 435978
rect 358174 435922 358242 435978
rect 358298 435922 358368 435978
rect 358048 435888 358368 435922
rect 388768 436350 389088 436384
rect 388768 436294 388838 436350
rect 388894 436294 388962 436350
rect 389018 436294 389088 436350
rect 388768 436226 389088 436294
rect 388768 436170 388838 436226
rect 388894 436170 388962 436226
rect 389018 436170 389088 436226
rect 388768 436102 389088 436170
rect 388768 436046 388838 436102
rect 388894 436046 388962 436102
rect 389018 436046 389088 436102
rect 388768 435978 389088 436046
rect 388768 435922 388838 435978
rect 388894 435922 388962 435978
rect 389018 435922 389088 435978
rect 388768 435888 389088 435922
rect 419488 436350 419808 436384
rect 419488 436294 419558 436350
rect 419614 436294 419682 436350
rect 419738 436294 419808 436350
rect 419488 436226 419808 436294
rect 419488 436170 419558 436226
rect 419614 436170 419682 436226
rect 419738 436170 419808 436226
rect 419488 436102 419808 436170
rect 419488 436046 419558 436102
rect 419614 436046 419682 436102
rect 419738 436046 419808 436102
rect 419488 435978 419808 436046
rect 419488 435922 419558 435978
rect 419614 435922 419682 435978
rect 419738 435922 419808 435978
rect 419488 435888 419808 435922
rect 450208 436350 450528 436384
rect 450208 436294 450278 436350
rect 450334 436294 450402 436350
rect 450458 436294 450528 436350
rect 450208 436226 450528 436294
rect 450208 436170 450278 436226
rect 450334 436170 450402 436226
rect 450458 436170 450528 436226
rect 450208 436102 450528 436170
rect 450208 436046 450278 436102
rect 450334 436046 450402 436102
rect 450458 436046 450528 436102
rect 450208 435978 450528 436046
rect 450208 435922 450278 435978
rect 450334 435922 450402 435978
rect 450458 435922 450528 435978
rect 450208 435888 450528 435922
rect 480928 436350 481248 436384
rect 480928 436294 480998 436350
rect 481054 436294 481122 436350
rect 481178 436294 481248 436350
rect 480928 436226 481248 436294
rect 480928 436170 480998 436226
rect 481054 436170 481122 436226
rect 481178 436170 481248 436226
rect 480928 436102 481248 436170
rect 480928 436046 480998 436102
rect 481054 436046 481122 436102
rect 481178 436046 481248 436102
rect 480928 435978 481248 436046
rect 480928 435922 480998 435978
rect 481054 435922 481122 435978
rect 481178 435922 481248 435978
rect 480928 435888 481248 435922
rect 507154 436350 507774 453922
rect 507154 436294 507250 436350
rect 507306 436294 507374 436350
rect 507430 436294 507498 436350
rect 507554 436294 507622 436350
rect 507678 436294 507774 436350
rect 507154 436226 507774 436294
rect 507154 436170 507250 436226
rect 507306 436170 507374 436226
rect 507430 436170 507498 436226
rect 507554 436170 507622 436226
rect 507678 436170 507774 436226
rect 507154 436102 507774 436170
rect 507154 436046 507250 436102
rect 507306 436046 507374 436102
rect 507430 436046 507498 436102
rect 507554 436046 507622 436102
rect 507678 436046 507774 436102
rect 507154 435978 507774 436046
rect 507154 435922 507250 435978
rect 507306 435922 507374 435978
rect 507430 435922 507498 435978
rect 507554 435922 507622 435978
rect 507678 435922 507774 435978
rect 219808 424350 220128 424384
rect 219808 424294 219878 424350
rect 219934 424294 220002 424350
rect 220058 424294 220128 424350
rect 219808 424226 220128 424294
rect 219808 424170 219878 424226
rect 219934 424170 220002 424226
rect 220058 424170 220128 424226
rect 219808 424102 220128 424170
rect 219808 424046 219878 424102
rect 219934 424046 220002 424102
rect 220058 424046 220128 424102
rect 219808 423978 220128 424046
rect 219808 423922 219878 423978
rect 219934 423922 220002 423978
rect 220058 423922 220128 423978
rect 219808 423888 220128 423922
rect 250528 424350 250848 424384
rect 250528 424294 250598 424350
rect 250654 424294 250722 424350
rect 250778 424294 250848 424350
rect 250528 424226 250848 424294
rect 250528 424170 250598 424226
rect 250654 424170 250722 424226
rect 250778 424170 250848 424226
rect 250528 424102 250848 424170
rect 250528 424046 250598 424102
rect 250654 424046 250722 424102
rect 250778 424046 250848 424102
rect 250528 423978 250848 424046
rect 250528 423922 250598 423978
rect 250654 423922 250722 423978
rect 250778 423922 250848 423978
rect 250528 423888 250848 423922
rect 281248 424350 281568 424384
rect 281248 424294 281318 424350
rect 281374 424294 281442 424350
rect 281498 424294 281568 424350
rect 281248 424226 281568 424294
rect 281248 424170 281318 424226
rect 281374 424170 281442 424226
rect 281498 424170 281568 424226
rect 281248 424102 281568 424170
rect 281248 424046 281318 424102
rect 281374 424046 281442 424102
rect 281498 424046 281568 424102
rect 281248 423978 281568 424046
rect 281248 423922 281318 423978
rect 281374 423922 281442 423978
rect 281498 423922 281568 423978
rect 281248 423888 281568 423922
rect 311968 424350 312288 424384
rect 311968 424294 312038 424350
rect 312094 424294 312162 424350
rect 312218 424294 312288 424350
rect 311968 424226 312288 424294
rect 311968 424170 312038 424226
rect 312094 424170 312162 424226
rect 312218 424170 312288 424226
rect 311968 424102 312288 424170
rect 311968 424046 312038 424102
rect 312094 424046 312162 424102
rect 312218 424046 312288 424102
rect 311968 423978 312288 424046
rect 311968 423922 312038 423978
rect 312094 423922 312162 423978
rect 312218 423922 312288 423978
rect 311968 423888 312288 423922
rect 342688 424350 343008 424384
rect 342688 424294 342758 424350
rect 342814 424294 342882 424350
rect 342938 424294 343008 424350
rect 342688 424226 343008 424294
rect 342688 424170 342758 424226
rect 342814 424170 342882 424226
rect 342938 424170 343008 424226
rect 342688 424102 343008 424170
rect 342688 424046 342758 424102
rect 342814 424046 342882 424102
rect 342938 424046 343008 424102
rect 342688 423978 343008 424046
rect 342688 423922 342758 423978
rect 342814 423922 342882 423978
rect 342938 423922 343008 423978
rect 342688 423888 343008 423922
rect 373408 424350 373728 424384
rect 373408 424294 373478 424350
rect 373534 424294 373602 424350
rect 373658 424294 373728 424350
rect 373408 424226 373728 424294
rect 373408 424170 373478 424226
rect 373534 424170 373602 424226
rect 373658 424170 373728 424226
rect 373408 424102 373728 424170
rect 373408 424046 373478 424102
rect 373534 424046 373602 424102
rect 373658 424046 373728 424102
rect 373408 423978 373728 424046
rect 373408 423922 373478 423978
rect 373534 423922 373602 423978
rect 373658 423922 373728 423978
rect 373408 423888 373728 423922
rect 404128 424350 404448 424384
rect 404128 424294 404198 424350
rect 404254 424294 404322 424350
rect 404378 424294 404448 424350
rect 404128 424226 404448 424294
rect 404128 424170 404198 424226
rect 404254 424170 404322 424226
rect 404378 424170 404448 424226
rect 404128 424102 404448 424170
rect 404128 424046 404198 424102
rect 404254 424046 404322 424102
rect 404378 424046 404448 424102
rect 404128 423978 404448 424046
rect 404128 423922 404198 423978
rect 404254 423922 404322 423978
rect 404378 423922 404448 423978
rect 404128 423888 404448 423922
rect 434848 424350 435168 424384
rect 434848 424294 434918 424350
rect 434974 424294 435042 424350
rect 435098 424294 435168 424350
rect 434848 424226 435168 424294
rect 434848 424170 434918 424226
rect 434974 424170 435042 424226
rect 435098 424170 435168 424226
rect 434848 424102 435168 424170
rect 434848 424046 434918 424102
rect 434974 424046 435042 424102
rect 435098 424046 435168 424102
rect 434848 423978 435168 424046
rect 434848 423922 434918 423978
rect 434974 423922 435042 423978
rect 435098 423922 435168 423978
rect 434848 423888 435168 423922
rect 465568 424350 465888 424384
rect 465568 424294 465638 424350
rect 465694 424294 465762 424350
rect 465818 424294 465888 424350
rect 465568 424226 465888 424294
rect 465568 424170 465638 424226
rect 465694 424170 465762 424226
rect 465818 424170 465888 424226
rect 465568 424102 465888 424170
rect 465568 424046 465638 424102
rect 465694 424046 465762 424102
rect 465818 424046 465888 424102
rect 465568 423978 465888 424046
rect 465568 423922 465638 423978
rect 465694 423922 465762 423978
rect 465818 423922 465888 423978
rect 465568 423888 465888 423922
rect 496288 424350 496608 424384
rect 496288 424294 496358 424350
rect 496414 424294 496482 424350
rect 496538 424294 496608 424350
rect 496288 424226 496608 424294
rect 496288 424170 496358 424226
rect 496414 424170 496482 424226
rect 496538 424170 496608 424226
rect 496288 424102 496608 424170
rect 496288 424046 496358 424102
rect 496414 424046 496482 424102
rect 496538 424046 496608 424102
rect 496288 423978 496608 424046
rect 496288 423922 496358 423978
rect 496414 423922 496482 423978
rect 496538 423922 496608 423978
rect 496288 423888 496608 423922
rect 201154 418294 201250 418350
rect 201306 418294 201374 418350
rect 201430 418294 201498 418350
rect 201554 418294 201622 418350
rect 201678 418294 201774 418350
rect 201154 418226 201774 418294
rect 201154 418170 201250 418226
rect 201306 418170 201374 418226
rect 201430 418170 201498 418226
rect 201554 418170 201622 418226
rect 201678 418170 201774 418226
rect 201154 418102 201774 418170
rect 201154 418046 201250 418102
rect 201306 418046 201374 418102
rect 201430 418046 201498 418102
rect 201554 418046 201622 418102
rect 201678 418046 201774 418102
rect 201154 417978 201774 418046
rect 201154 417922 201250 417978
rect 201306 417922 201374 417978
rect 201430 417922 201498 417978
rect 201554 417922 201622 417978
rect 201678 417922 201774 417978
rect 201154 400350 201774 417922
rect 204448 418350 204768 418384
rect 204448 418294 204518 418350
rect 204574 418294 204642 418350
rect 204698 418294 204768 418350
rect 204448 418226 204768 418294
rect 204448 418170 204518 418226
rect 204574 418170 204642 418226
rect 204698 418170 204768 418226
rect 204448 418102 204768 418170
rect 204448 418046 204518 418102
rect 204574 418046 204642 418102
rect 204698 418046 204768 418102
rect 204448 417978 204768 418046
rect 204448 417922 204518 417978
rect 204574 417922 204642 417978
rect 204698 417922 204768 417978
rect 204448 417888 204768 417922
rect 235168 418350 235488 418384
rect 235168 418294 235238 418350
rect 235294 418294 235362 418350
rect 235418 418294 235488 418350
rect 235168 418226 235488 418294
rect 235168 418170 235238 418226
rect 235294 418170 235362 418226
rect 235418 418170 235488 418226
rect 235168 418102 235488 418170
rect 235168 418046 235238 418102
rect 235294 418046 235362 418102
rect 235418 418046 235488 418102
rect 235168 417978 235488 418046
rect 235168 417922 235238 417978
rect 235294 417922 235362 417978
rect 235418 417922 235488 417978
rect 235168 417888 235488 417922
rect 265888 418350 266208 418384
rect 265888 418294 265958 418350
rect 266014 418294 266082 418350
rect 266138 418294 266208 418350
rect 265888 418226 266208 418294
rect 265888 418170 265958 418226
rect 266014 418170 266082 418226
rect 266138 418170 266208 418226
rect 265888 418102 266208 418170
rect 265888 418046 265958 418102
rect 266014 418046 266082 418102
rect 266138 418046 266208 418102
rect 265888 417978 266208 418046
rect 265888 417922 265958 417978
rect 266014 417922 266082 417978
rect 266138 417922 266208 417978
rect 265888 417888 266208 417922
rect 296608 418350 296928 418384
rect 296608 418294 296678 418350
rect 296734 418294 296802 418350
rect 296858 418294 296928 418350
rect 296608 418226 296928 418294
rect 296608 418170 296678 418226
rect 296734 418170 296802 418226
rect 296858 418170 296928 418226
rect 296608 418102 296928 418170
rect 296608 418046 296678 418102
rect 296734 418046 296802 418102
rect 296858 418046 296928 418102
rect 296608 417978 296928 418046
rect 296608 417922 296678 417978
rect 296734 417922 296802 417978
rect 296858 417922 296928 417978
rect 296608 417888 296928 417922
rect 327328 418350 327648 418384
rect 327328 418294 327398 418350
rect 327454 418294 327522 418350
rect 327578 418294 327648 418350
rect 327328 418226 327648 418294
rect 327328 418170 327398 418226
rect 327454 418170 327522 418226
rect 327578 418170 327648 418226
rect 327328 418102 327648 418170
rect 327328 418046 327398 418102
rect 327454 418046 327522 418102
rect 327578 418046 327648 418102
rect 327328 417978 327648 418046
rect 327328 417922 327398 417978
rect 327454 417922 327522 417978
rect 327578 417922 327648 417978
rect 327328 417888 327648 417922
rect 358048 418350 358368 418384
rect 358048 418294 358118 418350
rect 358174 418294 358242 418350
rect 358298 418294 358368 418350
rect 358048 418226 358368 418294
rect 358048 418170 358118 418226
rect 358174 418170 358242 418226
rect 358298 418170 358368 418226
rect 358048 418102 358368 418170
rect 358048 418046 358118 418102
rect 358174 418046 358242 418102
rect 358298 418046 358368 418102
rect 358048 417978 358368 418046
rect 358048 417922 358118 417978
rect 358174 417922 358242 417978
rect 358298 417922 358368 417978
rect 358048 417888 358368 417922
rect 388768 418350 389088 418384
rect 388768 418294 388838 418350
rect 388894 418294 388962 418350
rect 389018 418294 389088 418350
rect 388768 418226 389088 418294
rect 388768 418170 388838 418226
rect 388894 418170 388962 418226
rect 389018 418170 389088 418226
rect 388768 418102 389088 418170
rect 388768 418046 388838 418102
rect 388894 418046 388962 418102
rect 389018 418046 389088 418102
rect 388768 417978 389088 418046
rect 388768 417922 388838 417978
rect 388894 417922 388962 417978
rect 389018 417922 389088 417978
rect 388768 417888 389088 417922
rect 419488 418350 419808 418384
rect 419488 418294 419558 418350
rect 419614 418294 419682 418350
rect 419738 418294 419808 418350
rect 419488 418226 419808 418294
rect 419488 418170 419558 418226
rect 419614 418170 419682 418226
rect 419738 418170 419808 418226
rect 419488 418102 419808 418170
rect 419488 418046 419558 418102
rect 419614 418046 419682 418102
rect 419738 418046 419808 418102
rect 419488 417978 419808 418046
rect 419488 417922 419558 417978
rect 419614 417922 419682 417978
rect 419738 417922 419808 417978
rect 419488 417888 419808 417922
rect 450208 418350 450528 418384
rect 450208 418294 450278 418350
rect 450334 418294 450402 418350
rect 450458 418294 450528 418350
rect 450208 418226 450528 418294
rect 450208 418170 450278 418226
rect 450334 418170 450402 418226
rect 450458 418170 450528 418226
rect 450208 418102 450528 418170
rect 450208 418046 450278 418102
rect 450334 418046 450402 418102
rect 450458 418046 450528 418102
rect 450208 417978 450528 418046
rect 450208 417922 450278 417978
rect 450334 417922 450402 417978
rect 450458 417922 450528 417978
rect 450208 417888 450528 417922
rect 480928 418350 481248 418384
rect 480928 418294 480998 418350
rect 481054 418294 481122 418350
rect 481178 418294 481248 418350
rect 480928 418226 481248 418294
rect 480928 418170 480998 418226
rect 481054 418170 481122 418226
rect 481178 418170 481248 418226
rect 480928 418102 481248 418170
rect 480928 418046 480998 418102
rect 481054 418046 481122 418102
rect 481178 418046 481248 418102
rect 480928 417978 481248 418046
rect 480928 417922 480998 417978
rect 481054 417922 481122 417978
rect 481178 417922 481248 417978
rect 480928 417888 481248 417922
rect 507154 418350 507774 435922
rect 507154 418294 507250 418350
rect 507306 418294 507374 418350
rect 507430 418294 507498 418350
rect 507554 418294 507622 418350
rect 507678 418294 507774 418350
rect 507154 418226 507774 418294
rect 507154 418170 507250 418226
rect 507306 418170 507374 418226
rect 507430 418170 507498 418226
rect 507554 418170 507622 418226
rect 507678 418170 507774 418226
rect 507154 418102 507774 418170
rect 507154 418046 507250 418102
rect 507306 418046 507374 418102
rect 507430 418046 507498 418102
rect 507554 418046 507622 418102
rect 507678 418046 507774 418102
rect 507154 417978 507774 418046
rect 507154 417922 507250 417978
rect 507306 417922 507374 417978
rect 507430 417922 507498 417978
rect 507554 417922 507622 417978
rect 507678 417922 507774 417978
rect 219808 406350 220128 406384
rect 219808 406294 219878 406350
rect 219934 406294 220002 406350
rect 220058 406294 220128 406350
rect 219808 406226 220128 406294
rect 219808 406170 219878 406226
rect 219934 406170 220002 406226
rect 220058 406170 220128 406226
rect 219808 406102 220128 406170
rect 219808 406046 219878 406102
rect 219934 406046 220002 406102
rect 220058 406046 220128 406102
rect 219808 405978 220128 406046
rect 219808 405922 219878 405978
rect 219934 405922 220002 405978
rect 220058 405922 220128 405978
rect 219808 405888 220128 405922
rect 250528 406350 250848 406384
rect 250528 406294 250598 406350
rect 250654 406294 250722 406350
rect 250778 406294 250848 406350
rect 250528 406226 250848 406294
rect 250528 406170 250598 406226
rect 250654 406170 250722 406226
rect 250778 406170 250848 406226
rect 250528 406102 250848 406170
rect 250528 406046 250598 406102
rect 250654 406046 250722 406102
rect 250778 406046 250848 406102
rect 250528 405978 250848 406046
rect 250528 405922 250598 405978
rect 250654 405922 250722 405978
rect 250778 405922 250848 405978
rect 250528 405888 250848 405922
rect 281248 406350 281568 406384
rect 281248 406294 281318 406350
rect 281374 406294 281442 406350
rect 281498 406294 281568 406350
rect 281248 406226 281568 406294
rect 281248 406170 281318 406226
rect 281374 406170 281442 406226
rect 281498 406170 281568 406226
rect 281248 406102 281568 406170
rect 281248 406046 281318 406102
rect 281374 406046 281442 406102
rect 281498 406046 281568 406102
rect 281248 405978 281568 406046
rect 281248 405922 281318 405978
rect 281374 405922 281442 405978
rect 281498 405922 281568 405978
rect 281248 405888 281568 405922
rect 311968 406350 312288 406384
rect 311968 406294 312038 406350
rect 312094 406294 312162 406350
rect 312218 406294 312288 406350
rect 311968 406226 312288 406294
rect 311968 406170 312038 406226
rect 312094 406170 312162 406226
rect 312218 406170 312288 406226
rect 311968 406102 312288 406170
rect 311968 406046 312038 406102
rect 312094 406046 312162 406102
rect 312218 406046 312288 406102
rect 311968 405978 312288 406046
rect 311968 405922 312038 405978
rect 312094 405922 312162 405978
rect 312218 405922 312288 405978
rect 311968 405888 312288 405922
rect 342688 406350 343008 406384
rect 342688 406294 342758 406350
rect 342814 406294 342882 406350
rect 342938 406294 343008 406350
rect 342688 406226 343008 406294
rect 342688 406170 342758 406226
rect 342814 406170 342882 406226
rect 342938 406170 343008 406226
rect 342688 406102 343008 406170
rect 342688 406046 342758 406102
rect 342814 406046 342882 406102
rect 342938 406046 343008 406102
rect 342688 405978 343008 406046
rect 342688 405922 342758 405978
rect 342814 405922 342882 405978
rect 342938 405922 343008 405978
rect 342688 405888 343008 405922
rect 373408 406350 373728 406384
rect 373408 406294 373478 406350
rect 373534 406294 373602 406350
rect 373658 406294 373728 406350
rect 373408 406226 373728 406294
rect 373408 406170 373478 406226
rect 373534 406170 373602 406226
rect 373658 406170 373728 406226
rect 373408 406102 373728 406170
rect 373408 406046 373478 406102
rect 373534 406046 373602 406102
rect 373658 406046 373728 406102
rect 373408 405978 373728 406046
rect 373408 405922 373478 405978
rect 373534 405922 373602 405978
rect 373658 405922 373728 405978
rect 373408 405888 373728 405922
rect 404128 406350 404448 406384
rect 404128 406294 404198 406350
rect 404254 406294 404322 406350
rect 404378 406294 404448 406350
rect 404128 406226 404448 406294
rect 404128 406170 404198 406226
rect 404254 406170 404322 406226
rect 404378 406170 404448 406226
rect 404128 406102 404448 406170
rect 404128 406046 404198 406102
rect 404254 406046 404322 406102
rect 404378 406046 404448 406102
rect 404128 405978 404448 406046
rect 404128 405922 404198 405978
rect 404254 405922 404322 405978
rect 404378 405922 404448 405978
rect 404128 405888 404448 405922
rect 434848 406350 435168 406384
rect 434848 406294 434918 406350
rect 434974 406294 435042 406350
rect 435098 406294 435168 406350
rect 434848 406226 435168 406294
rect 434848 406170 434918 406226
rect 434974 406170 435042 406226
rect 435098 406170 435168 406226
rect 434848 406102 435168 406170
rect 434848 406046 434918 406102
rect 434974 406046 435042 406102
rect 435098 406046 435168 406102
rect 434848 405978 435168 406046
rect 434848 405922 434918 405978
rect 434974 405922 435042 405978
rect 435098 405922 435168 405978
rect 434848 405888 435168 405922
rect 465568 406350 465888 406384
rect 465568 406294 465638 406350
rect 465694 406294 465762 406350
rect 465818 406294 465888 406350
rect 465568 406226 465888 406294
rect 465568 406170 465638 406226
rect 465694 406170 465762 406226
rect 465818 406170 465888 406226
rect 465568 406102 465888 406170
rect 465568 406046 465638 406102
rect 465694 406046 465762 406102
rect 465818 406046 465888 406102
rect 465568 405978 465888 406046
rect 465568 405922 465638 405978
rect 465694 405922 465762 405978
rect 465818 405922 465888 405978
rect 465568 405888 465888 405922
rect 496288 406350 496608 406384
rect 496288 406294 496358 406350
rect 496414 406294 496482 406350
rect 496538 406294 496608 406350
rect 496288 406226 496608 406294
rect 496288 406170 496358 406226
rect 496414 406170 496482 406226
rect 496538 406170 496608 406226
rect 496288 406102 496608 406170
rect 496288 406046 496358 406102
rect 496414 406046 496482 406102
rect 496538 406046 496608 406102
rect 496288 405978 496608 406046
rect 496288 405922 496358 405978
rect 496414 405922 496482 405978
rect 496538 405922 496608 405978
rect 496288 405888 496608 405922
rect 201154 400294 201250 400350
rect 201306 400294 201374 400350
rect 201430 400294 201498 400350
rect 201554 400294 201622 400350
rect 201678 400294 201774 400350
rect 201154 400226 201774 400294
rect 201154 400170 201250 400226
rect 201306 400170 201374 400226
rect 201430 400170 201498 400226
rect 201554 400170 201622 400226
rect 201678 400170 201774 400226
rect 201154 400102 201774 400170
rect 201154 400046 201250 400102
rect 201306 400046 201374 400102
rect 201430 400046 201498 400102
rect 201554 400046 201622 400102
rect 201678 400046 201774 400102
rect 201154 399978 201774 400046
rect 201154 399922 201250 399978
rect 201306 399922 201374 399978
rect 201430 399922 201498 399978
rect 201554 399922 201622 399978
rect 201678 399922 201774 399978
rect 201154 382350 201774 399922
rect 204448 400350 204768 400384
rect 204448 400294 204518 400350
rect 204574 400294 204642 400350
rect 204698 400294 204768 400350
rect 204448 400226 204768 400294
rect 204448 400170 204518 400226
rect 204574 400170 204642 400226
rect 204698 400170 204768 400226
rect 204448 400102 204768 400170
rect 204448 400046 204518 400102
rect 204574 400046 204642 400102
rect 204698 400046 204768 400102
rect 204448 399978 204768 400046
rect 204448 399922 204518 399978
rect 204574 399922 204642 399978
rect 204698 399922 204768 399978
rect 204448 399888 204768 399922
rect 235168 400350 235488 400384
rect 235168 400294 235238 400350
rect 235294 400294 235362 400350
rect 235418 400294 235488 400350
rect 235168 400226 235488 400294
rect 235168 400170 235238 400226
rect 235294 400170 235362 400226
rect 235418 400170 235488 400226
rect 235168 400102 235488 400170
rect 235168 400046 235238 400102
rect 235294 400046 235362 400102
rect 235418 400046 235488 400102
rect 235168 399978 235488 400046
rect 235168 399922 235238 399978
rect 235294 399922 235362 399978
rect 235418 399922 235488 399978
rect 235168 399888 235488 399922
rect 265888 400350 266208 400384
rect 265888 400294 265958 400350
rect 266014 400294 266082 400350
rect 266138 400294 266208 400350
rect 265888 400226 266208 400294
rect 265888 400170 265958 400226
rect 266014 400170 266082 400226
rect 266138 400170 266208 400226
rect 265888 400102 266208 400170
rect 265888 400046 265958 400102
rect 266014 400046 266082 400102
rect 266138 400046 266208 400102
rect 265888 399978 266208 400046
rect 265888 399922 265958 399978
rect 266014 399922 266082 399978
rect 266138 399922 266208 399978
rect 265888 399888 266208 399922
rect 296608 400350 296928 400384
rect 296608 400294 296678 400350
rect 296734 400294 296802 400350
rect 296858 400294 296928 400350
rect 296608 400226 296928 400294
rect 296608 400170 296678 400226
rect 296734 400170 296802 400226
rect 296858 400170 296928 400226
rect 296608 400102 296928 400170
rect 296608 400046 296678 400102
rect 296734 400046 296802 400102
rect 296858 400046 296928 400102
rect 296608 399978 296928 400046
rect 296608 399922 296678 399978
rect 296734 399922 296802 399978
rect 296858 399922 296928 399978
rect 296608 399888 296928 399922
rect 327328 400350 327648 400384
rect 327328 400294 327398 400350
rect 327454 400294 327522 400350
rect 327578 400294 327648 400350
rect 327328 400226 327648 400294
rect 327328 400170 327398 400226
rect 327454 400170 327522 400226
rect 327578 400170 327648 400226
rect 327328 400102 327648 400170
rect 327328 400046 327398 400102
rect 327454 400046 327522 400102
rect 327578 400046 327648 400102
rect 327328 399978 327648 400046
rect 327328 399922 327398 399978
rect 327454 399922 327522 399978
rect 327578 399922 327648 399978
rect 327328 399888 327648 399922
rect 358048 400350 358368 400384
rect 358048 400294 358118 400350
rect 358174 400294 358242 400350
rect 358298 400294 358368 400350
rect 358048 400226 358368 400294
rect 358048 400170 358118 400226
rect 358174 400170 358242 400226
rect 358298 400170 358368 400226
rect 358048 400102 358368 400170
rect 358048 400046 358118 400102
rect 358174 400046 358242 400102
rect 358298 400046 358368 400102
rect 358048 399978 358368 400046
rect 358048 399922 358118 399978
rect 358174 399922 358242 399978
rect 358298 399922 358368 399978
rect 358048 399888 358368 399922
rect 388768 400350 389088 400384
rect 388768 400294 388838 400350
rect 388894 400294 388962 400350
rect 389018 400294 389088 400350
rect 388768 400226 389088 400294
rect 388768 400170 388838 400226
rect 388894 400170 388962 400226
rect 389018 400170 389088 400226
rect 388768 400102 389088 400170
rect 388768 400046 388838 400102
rect 388894 400046 388962 400102
rect 389018 400046 389088 400102
rect 388768 399978 389088 400046
rect 388768 399922 388838 399978
rect 388894 399922 388962 399978
rect 389018 399922 389088 399978
rect 388768 399888 389088 399922
rect 419488 400350 419808 400384
rect 419488 400294 419558 400350
rect 419614 400294 419682 400350
rect 419738 400294 419808 400350
rect 419488 400226 419808 400294
rect 419488 400170 419558 400226
rect 419614 400170 419682 400226
rect 419738 400170 419808 400226
rect 419488 400102 419808 400170
rect 419488 400046 419558 400102
rect 419614 400046 419682 400102
rect 419738 400046 419808 400102
rect 419488 399978 419808 400046
rect 419488 399922 419558 399978
rect 419614 399922 419682 399978
rect 419738 399922 419808 399978
rect 419488 399888 419808 399922
rect 450208 400350 450528 400384
rect 450208 400294 450278 400350
rect 450334 400294 450402 400350
rect 450458 400294 450528 400350
rect 450208 400226 450528 400294
rect 450208 400170 450278 400226
rect 450334 400170 450402 400226
rect 450458 400170 450528 400226
rect 450208 400102 450528 400170
rect 450208 400046 450278 400102
rect 450334 400046 450402 400102
rect 450458 400046 450528 400102
rect 450208 399978 450528 400046
rect 450208 399922 450278 399978
rect 450334 399922 450402 399978
rect 450458 399922 450528 399978
rect 450208 399888 450528 399922
rect 480928 400350 481248 400384
rect 480928 400294 480998 400350
rect 481054 400294 481122 400350
rect 481178 400294 481248 400350
rect 480928 400226 481248 400294
rect 480928 400170 480998 400226
rect 481054 400170 481122 400226
rect 481178 400170 481248 400226
rect 480928 400102 481248 400170
rect 480928 400046 480998 400102
rect 481054 400046 481122 400102
rect 481178 400046 481248 400102
rect 480928 399978 481248 400046
rect 480928 399922 480998 399978
rect 481054 399922 481122 399978
rect 481178 399922 481248 399978
rect 480928 399888 481248 399922
rect 507154 400350 507774 417922
rect 507154 400294 507250 400350
rect 507306 400294 507374 400350
rect 507430 400294 507498 400350
rect 507554 400294 507622 400350
rect 507678 400294 507774 400350
rect 507154 400226 507774 400294
rect 507154 400170 507250 400226
rect 507306 400170 507374 400226
rect 507430 400170 507498 400226
rect 507554 400170 507622 400226
rect 507678 400170 507774 400226
rect 507154 400102 507774 400170
rect 507154 400046 507250 400102
rect 507306 400046 507374 400102
rect 507430 400046 507498 400102
rect 507554 400046 507622 400102
rect 507678 400046 507774 400102
rect 507154 399978 507774 400046
rect 507154 399922 507250 399978
rect 507306 399922 507374 399978
rect 507430 399922 507498 399978
rect 507554 399922 507622 399978
rect 507678 399922 507774 399978
rect 219808 388350 220128 388384
rect 219808 388294 219878 388350
rect 219934 388294 220002 388350
rect 220058 388294 220128 388350
rect 219808 388226 220128 388294
rect 219808 388170 219878 388226
rect 219934 388170 220002 388226
rect 220058 388170 220128 388226
rect 219808 388102 220128 388170
rect 219808 388046 219878 388102
rect 219934 388046 220002 388102
rect 220058 388046 220128 388102
rect 219808 387978 220128 388046
rect 219808 387922 219878 387978
rect 219934 387922 220002 387978
rect 220058 387922 220128 387978
rect 219808 387888 220128 387922
rect 250528 388350 250848 388384
rect 250528 388294 250598 388350
rect 250654 388294 250722 388350
rect 250778 388294 250848 388350
rect 250528 388226 250848 388294
rect 250528 388170 250598 388226
rect 250654 388170 250722 388226
rect 250778 388170 250848 388226
rect 250528 388102 250848 388170
rect 250528 388046 250598 388102
rect 250654 388046 250722 388102
rect 250778 388046 250848 388102
rect 250528 387978 250848 388046
rect 250528 387922 250598 387978
rect 250654 387922 250722 387978
rect 250778 387922 250848 387978
rect 250528 387888 250848 387922
rect 281248 388350 281568 388384
rect 281248 388294 281318 388350
rect 281374 388294 281442 388350
rect 281498 388294 281568 388350
rect 281248 388226 281568 388294
rect 281248 388170 281318 388226
rect 281374 388170 281442 388226
rect 281498 388170 281568 388226
rect 281248 388102 281568 388170
rect 281248 388046 281318 388102
rect 281374 388046 281442 388102
rect 281498 388046 281568 388102
rect 281248 387978 281568 388046
rect 281248 387922 281318 387978
rect 281374 387922 281442 387978
rect 281498 387922 281568 387978
rect 281248 387888 281568 387922
rect 311968 388350 312288 388384
rect 311968 388294 312038 388350
rect 312094 388294 312162 388350
rect 312218 388294 312288 388350
rect 311968 388226 312288 388294
rect 311968 388170 312038 388226
rect 312094 388170 312162 388226
rect 312218 388170 312288 388226
rect 311968 388102 312288 388170
rect 311968 388046 312038 388102
rect 312094 388046 312162 388102
rect 312218 388046 312288 388102
rect 311968 387978 312288 388046
rect 311968 387922 312038 387978
rect 312094 387922 312162 387978
rect 312218 387922 312288 387978
rect 311968 387888 312288 387922
rect 342688 388350 343008 388384
rect 342688 388294 342758 388350
rect 342814 388294 342882 388350
rect 342938 388294 343008 388350
rect 342688 388226 343008 388294
rect 342688 388170 342758 388226
rect 342814 388170 342882 388226
rect 342938 388170 343008 388226
rect 342688 388102 343008 388170
rect 342688 388046 342758 388102
rect 342814 388046 342882 388102
rect 342938 388046 343008 388102
rect 342688 387978 343008 388046
rect 342688 387922 342758 387978
rect 342814 387922 342882 387978
rect 342938 387922 343008 387978
rect 342688 387888 343008 387922
rect 373408 388350 373728 388384
rect 373408 388294 373478 388350
rect 373534 388294 373602 388350
rect 373658 388294 373728 388350
rect 373408 388226 373728 388294
rect 373408 388170 373478 388226
rect 373534 388170 373602 388226
rect 373658 388170 373728 388226
rect 373408 388102 373728 388170
rect 373408 388046 373478 388102
rect 373534 388046 373602 388102
rect 373658 388046 373728 388102
rect 373408 387978 373728 388046
rect 373408 387922 373478 387978
rect 373534 387922 373602 387978
rect 373658 387922 373728 387978
rect 373408 387888 373728 387922
rect 404128 388350 404448 388384
rect 404128 388294 404198 388350
rect 404254 388294 404322 388350
rect 404378 388294 404448 388350
rect 404128 388226 404448 388294
rect 404128 388170 404198 388226
rect 404254 388170 404322 388226
rect 404378 388170 404448 388226
rect 404128 388102 404448 388170
rect 404128 388046 404198 388102
rect 404254 388046 404322 388102
rect 404378 388046 404448 388102
rect 404128 387978 404448 388046
rect 404128 387922 404198 387978
rect 404254 387922 404322 387978
rect 404378 387922 404448 387978
rect 404128 387888 404448 387922
rect 434848 388350 435168 388384
rect 434848 388294 434918 388350
rect 434974 388294 435042 388350
rect 435098 388294 435168 388350
rect 434848 388226 435168 388294
rect 434848 388170 434918 388226
rect 434974 388170 435042 388226
rect 435098 388170 435168 388226
rect 434848 388102 435168 388170
rect 434848 388046 434918 388102
rect 434974 388046 435042 388102
rect 435098 388046 435168 388102
rect 434848 387978 435168 388046
rect 434848 387922 434918 387978
rect 434974 387922 435042 387978
rect 435098 387922 435168 387978
rect 434848 387888 435168 387922
rect 465568 388350 465888 388384
rect 465568 388294 465638 388350
rect 465694 388294 465762 388350
rect 465818 388294 465888 388350
rect 465568 388226 465888 388294
rect 465568 388170 465638 388226
rect 465694 388170 465762 388226
rect 465818 388170 465888 388226
rect 465568 388102 465888 388170
rect 465568 388046 465638 388102
rect 465694 388046 465762 388102
rect 465818 388046 465888 388102
rect 465568 387978 465888 388046
rect 465568 387922 465638 387978
rect 465694 387922 465762 387978
rect 465818 387922 465888 387978
rect 465568 387888 465888 387922
rect 496288 388350 496608 388384
rect 496288 388294 496358 388350
rect 496414 388294 496482 388350
rect 496538 388294 496608 388350
rect 496288 388226 496608 388294
rect 496288 388170 496358 388226
rect 496414 388170 496482 388226
rect 496538 388170 496608 388226
rect 496288 388102 496608 388170
rect 496288 388046 496358 388102
rect 496414 388046 496482 388102
rect 496538 388046 496608 388102
rect 496288 387978 496608 388046
rect 496288 387922 496358 387978
rect 496414 387922 496482 387978
rect 496538 387922 496608 387978
rect 496288 387888 496608 387922
rect 201154 382294 201250 382350
rect 201306 382294 201374 382350
rect 201430 382294 201498 382350
rect 201554 382294 201622 382350
rect 201678 382294 201774 382350
rect 201154 382226 201774 382294
rect 201154 382170 201250 382226
rect 201306 382170 201374 382226
rect 201430 382170 201498 382226
rect 201554 382170 201622 382226
rect 201678 382170 201774 382226
rect 201154 382102 201774 382170
rect 201154 382046 201250 382102
rect 201306 382046 201374 382102
rect 201430 382046 201498 382102
rect 201554 382046 201622 382102
rect 201678 382046 201774 382102
rect 201154 381978 201774 382046
rect 201154 381922 201250 381978
rect 201306 381922 201374 381978
rect 201430 381922 201498 381978
rect 201554 381922 201622 381978
rect 201678 381922 201774 381978
rect 201154 364350 201774 381922
rect 204448 382350 204768 382384
rect 204448 382294 204518 382350
rect 204574 382294 204642 382350
rect 204698 382294 204768 382350
rect 204448 382226 204768 382294
rect 204448 382170 204518 382226
rect 204574 382170 204642 382226
rect 204698 382170 204768 382226
rect 204448 382102 204768 382170
rect 204448 382046 204518 382102
rect 204574 382046 204642 382102
rect 204698 382046 204768 382102
rect 204448 381978 204768 382046
rect 204448 381922 204518 381978
rect 204574 381922 204642 381978
rect 204698 381922 204768 381978
rect 204448 381888 204768 381922
rect 235168 382350 235488 382384
rect 235168 382294 235238 382350
rect 235294 382294 235362 382350
rect 235418 382294 235488 382350
rect 235168 382226 235488 382294
rect 235168 382170 235238 382226
rect 235294 382170 235362 382226
rect 235418 382170 235488 382226
rect 235168 382102 235488 382170
rect 235168 382046 235238 382102
rect 235294 382046 235362 382102
rect 235418 382046 235488 382102
rect 235168 381978 235488 382046
rect 235168 381922 235238 381978
rect 235294 381922 235362 381978
rect 235418 381922 235488 381978
rect 235168 381888 235488 381922
rect 265888 382350 266208 382384
rect 265888 382294 265958 382350
rect 266014 382294 266082 382350
rect 266138 382294 266208 382350
rect 265888 382226 266208 382294
rect 265888 382170 265958 382226
rect 266014 382170 266082 382226
rect 266138 382170 266208 382226
rect 265888 382102 266208 382170
rect 265888 382046 265958 382102
rect 266014 382046 266082 382102
rect 266138 382046 266208 382102
rect 265888 381978 266208 382046
rect 265888 381922 265958 381978
rect 266014 381922 266082 381978
rect 266138 381922 266208 381978
rect 265888 381888 266208 381922
rect 296608 382350 296928 382384
rect 296608 382294 296678 382350
rect 296734 382294 296802 382350
rect 296858 382294 296928 382350
rect 296608 382226 296928 382294
rect 296608 382170 296678 382226
rect 296734 382170 296802 382226
rect 296858 382170 296928 382226
rect 296608 382102 296928 382170
rect 296608 382046 296678 382102
rect 296734 382046 296802 382102
rect 296858 382046 296928 382102
rect 296608 381978 296928 382046
rect 296608 381922 296678 381978
rect 296734 381922 296802 381978
rect 296858 381922 296928 381978
rect 296608 381888 296928 381922
rect 327328 382350 327648 382384
rect 327328 382294 327398 382350
rect 327454 382294 327522 382350
rect 327578 382294 327648 382350
rect 327328 382226 327648 382294
rect 327328 382170 327398 382226
rect 327454 382170 327522 382226
rect 327578 382170 327648 382226
rect 327328 382102 327648 382170
rect 327328 382046 327398 382102
rect 327454 382046 327522 382102
rect 327578 382046 327648 382102
rect 327328 381978 327648 382046
rect 327328 381922 327398 381978
rect 327454 381922 327522 381978
rect 327578 381922 327648 381978
rect 327328 381888 327648 381922
rect 358048 382350 358368 382384
rect 358048 382294 358118 382350
rect 358174 382294 358242 382350
rect 358298 382294 358368 382350
rect 358048 382226 358368 382294
rect 358048 382170 358118 382226
rect 358174 382170 358242 382226
rect 358298 382170 358368 382226
rect 358048 382102 358368 382170
rect 358048 382046 358118 382102
rect 358174 382046 358242 382102
rect 358298 382046 358368 382102
rect 358048 381978 358368 382046
rect 358048 381922 358118 381978
rect 358174 381922 358242 381978
rect 358298 381922 358368 381978
rect 358048 381888 358368 381922
rect 388768 382350 389088 382384
rect 388768 382294 388838 382350
rect 388894 382294 388962 382350
rect 389018 382294 389088 382350
rect 388768 382226 389088 382294
rect 388768 382170 388838 382226
rect 388894 382170 388962 382226
rect 389018 382170 389088 382226
rect 388768 382102 389088 382170
rect 388768 382046 388838 382102
rect 388894 382046 388962 382102
rect 389018 382046 389088 382102
rect 388768 381978 389088 382046
rect 388768 381922 388838 381978
rect 388894 381922 388962 381978
rect 389018 381922 389088 381978
rect 388768 381888 389088 381922
rect 419488 382350 419808 382384
rect 419488 382294 419558 382350
rect 419614 382294 419682 382350
rect 419738 382294 419808 382350
rect 419488 382226 419808 382294
rect 419488 382170 419558 382226
rect 419614 382170 419682 382226
rect 419738 382170 419808 382226
rect 419488 382102 419808 382170
rect 419488 382046 419558 382102
rect 419614 382046 419682 382102
rect 419738 382046 419808 382102
rect 419488 381978 419808 382046
rect 419488 381922 419558 381978
rect 419614 381922 419682 381978
rect 419738 381922 419808 381978
rect 419488 381888 419808 381922
rect 450208 382350 450528 382384
rect 450208 382294 450278 382350
rect 450334 382294 450402 382350
rect 450458 382294 450528 382350
rect 450208 382226 450528 382294
rect 450208 382170 450278 382226
rect 450334 382170 450402 382226
rect 450458 382170 450528 382226
rect 450208 382102 450528 382170
rect 450208 382046 450278 382102
rect 450334 382046 450402 382102
rect 450458 382046 450528 382102
rect 450208 381978 450528 382046
rect 450208 381922 450278 381978
rect 450334 381922 450402 381978
rect 450458 381922 450528 381978
rect 450208 381888 450528 381922
rect 480928 382350 481248 382384
rect 480928 382294 480998 382350
rect 481054 382294 481122 382350
rect 481178 382294 481248 382350
rect 480928 382226 481248 382294
rect 480928 382170 480998 382226
rect 481054 382170 481122 382226
rect 481178 382170 481248 382226
rect 480928 382102 481248 382170
rect 480928 382046 480998 382102
rect 481054 382046 481122 382102
rect 481178 382046 481248 382102
rect 480928 381978 481248 382046
rect 480928 381922 480998 381978
rect 481054 381922 481122 381978
rect 481178 381922 481248 381978
rect 480928 381888 481248 381922
rect 507154 382350 507774 399922
rect 507154 382294 507250 382350
rect 507306 382294 507374 382350
rect 507430 382294 507498 382350
rect 507554 382294 507622 382350
rect 507678 382294 507774 382350
rect 507154 382226 507774 382294
rect 507154 382170 507250 382226
rect 507306 382170 507374 382226
rect 507430 382170 507498 382226
rect 507554 382170 507622 382226
rect 507678 382170 507774 382226
rect 507154 382102 507774 382170
rect 507154 382046 507250 382102
rect 507306 382046 507374 382102
rect 507430 382046 507498 382102
rect 507554 382046 507622 382102
rect 507678 382046 507774 382102
rect 507154 381978 507774 382046
rect 507154 381922 507250 381978
rect 507306 381922 507374 381978
rect 507430 381922 507498 381978
rect 507554 381922 507622 381978
rect 507678 381922 507774 381978
rect 219808 370350 220128 370384
rect 219808 370294 219878 370350
rect 219934 370294 220002 370350
rect 220058 370294 220128 370350
rect 219808 370226 220128 370294
rect 219808 370170 219878 370226
rect 219934 370170 220002 370226
rect 220058 370170 220128 370226
rect 219808 370102 220128 370170
rect 219808 370046 219878 370102
rect 219934 370046 220002 370102
rect 220058 370046 220128 370102
rect 219808 369978 220128 370046
rect 219808 369922 219878 369978
rect 219934 369922 220002 369978
rect 220058 369922 220128 369978
rect 219808 369888 220128 369922
rect 250528 370350 250848 370384
rect 250528 370294 250598 370350
rect 250654 370294 250722 370350
rect 250778 370294 250848 370350
rect 250528 370226 250848 370294
rect 250528 370170 250598 370226
rect 250654 370170 250722 370226
rect 250778 370170 250848 370226
rect 250528 370102 250848 370170
rect 250528 370046 250598 370102
rect 250654 370046 250722 370102
rect 250778 370046 250848 370102
rect 250528 369978 250848 370046
rect 250528 369922 250598 369978
rect 250654 369922 250722 369978
rect 250778 369922 250848 369978
rect 250528 369888 250848 369922
rect 281248 370350 281568 370384
rect 281248 370294 281318 370350
rect 281374 370294 281442 370350
rect 281498 370294 281568 370350
rect 281248 370226 281568 370294
rect 281248 370170 281318 370226
rect 281374 370170 281442 370226
rect 281498 370170 281568 370226
rect 281248 370102 281568 370170
rect 281248 370046 281318 370102
rect 281374 370046 281442 370102
rect 281498 370046 281568 370102
rect 281248 369978 281568 370046
rect 281248 369922 281318 369978
rect 281374 369922 281442 369978
rect 281498 369922 281568 369978
rect 281248 369888 281568 369922
rect 311968 370350 312288 370384
rect 311968 370294 312038 370350
rect 312094 370294 312162 370350
rect 312218 370294 312288 370350
rect 311968 370226 312288 370294
rect 311968 370170 312038 370226
rect 312094 370170 312162 370226
rect 312218 370170 312288 370226
rect 311968 370102 312288 370170
rect 311968 370046 312038 370102
rect 312094 370046 312162 370102
rect 312218 370046 312288 370102
rect 311968 369978 312288 370046
rect 311968 369922 312038 369978
rect 312094 369922 312162 369978
rect 312218 369922 312288 369978
rect 311968 369888 312288 369922
rect 342688 370350 343008 370384
rect 342688 370294 342758 370350
rect 342814 370294 342882 370350
rect 342938 370294 343008 370350
rect 342688 370226 343008 370294
rect 342688 370170 342758 370226
rect 342814 370170 342882 370226
rect 342938 370170 343008 370226
rect 342688 370102 343008 370170
rect 342688 370046 342758 370102
rect 342814 370046 342882 370102
rect 342938 370046 343008 370102
rect 342688 369978 343008 370046
rect 342688 369922 342758 369978
rect 342814 369922 342882 369978
rect 342938 369922 343008 369978
rect 342688 369888 343008 369922
rect 373408 370350 373728 370384
rect 373408 370294 373478 370350
rect 373534 370294 373602 370350
rect 373658 370294 373728 370350
rect 373408 370226 373728 370294
rect 373408 370170 373478 370226
rect 373534 370170 373602 370226
rect 373658 370170 373728 370226
rect 373408 370102 373728 370170
rect 373408 370046 373478 370102
rect 373534 370046 373602 370102
rect 373658 370046 373728 370102
rect 373408 369978 373728 370046
rect 373408 369922 373478 369978
rect 373534 369922 373602 369978
rect 373658 369922 373728 369978
rect 373408 369888 373728 369922
rect 404128 370350 404448 370384
rect 404128 370294 404198 370350
rect 404254 370294 404322 370350
rect 404378 370294 404448 370350
rect 404128 370226 404448 370294
rect 404128 370170 404198 370226
rect 404254 370170 404322 370226
rect 404378 370170 404448 370226
rect 404128 370102 404448 370170
rect 404128 370046 404198 370102
rect 404254 370046 404322 370102
rect 404378 370046 404448 370102
rect 404128 369978 404448 370046
rect 404128 369922 404198 369978
rect 404254 369922 404322 369978
rect 404378 369922 404448 369978
rect 404128 369888 404448 369922
rect 434848 370350 435168 370384
rect 434848 370294 434918 370350
rect 434974 370294 435042 370350
rect 435098 370294 435168 370350
rect 434848 370226 435168 370294
rect 434848 370170 434918 370226
rect 434974 370170 435042 370226
rect 435098 370170 435168 370226
rect 434848 370102 435168 370170
rect 434848 370046 434918 370102
rect 434974 370046 435042 370102
rect 435098 370046 435168 370102
rect 434848 369978 435168 370046
rect 434848 369922 434918 369978
rect 434974 369922 435042 369978
rect 435098 369922 435168 369978
rect 434848 369888 435168 369922
rect 465568 370350 465888 370384
rect 465568 370294 465638 370350
rect 465694 370294 465762 370350
rect 465818 370294 465888 370350
rect 465568 370226 465888 370294
rect 465568 370170 465638 370226
rect 465694 370170 465762 370226
rect 465818 370170 465888 370226
rect 465568 370102 465888 370170
rect 465568 370046 465638 370102
rect 465694 370046 465762 370102
rect 465818 370046 465888 370102
rect 465568 369978 465888 370046
rect 465568 369922 465638 369978
rect 465694 369922 465762 369978
rect 465818 369922 465888 369978
rect 465568 369888 465888 369922
rect 496288 370350 496608 370384
rect 496288 370294 496358 370350
rect 496414 370294 496482 370350
rect 496538 370294 496608 370350
rect 496288 370226 496608 370294
rect 496288 370170 496358 370226
rect 496414 370170 496482 370226
rect 496538 370170 496608 370226
rect 496288 370102 496608 370170
rect 496288 370046 496358 370102
rect 496414 370046 496482 370102
rect 496538 370046 496608 370102
rect 496288 369978 496608 370046
rect 496288 369922 496358 369978
rect 496414 369922 496482 369978
rect 496538 369922 496608 369978
rect 496288 369888 496608 369922
rect 201154 364294 201250 364350
rect 201306 364294 201374 364350
rect 201430 364294 201498 364350
rect 201554 364294 201622 364350
rect 201678 364294 201774 364350
rect 201154 364226 201774 364294
rect 201154 364170 201250 364226
rect 201306 364170 201374 364226
rect 201430 364170 201498 364226
rect 201554 364170 201622 364226
rect 201678 364170 201774 364226
rect 201154 364102 201774 364170
rect 201154 364046 201250 364102
rect 201306 364046 201374 364102
rect 201430 364046 201498 364102
rect 201554 364046 201622 364102
rect 201678 364046 201774 364102
rect 201154 363978 201774 364046
rect 201154 363922 201250 363978
rect 201306 363922 201374 363978
rect 201430 363922 201498 363978
rect 201554 363922 201622 363978
rect 201678 363922 201774 363978
rect 201154 346350 201774 363922
rect 204448 364350 204768 364384
rect 204448 364294 204518 364350
rect 204574 364294 204642 364350
rect 204698 364294 204768 364350
rect 204448 364226 204768 364294
rect 204448 364170 204518 364226
rect 204574 364170 204642 364226
rect 204698 364170 204768 364226
rect 204448 364102 204768 364170
rect 204448 364046 204518 364102
rect 204574 364046 204642 364102
rect 204698 364046 204768 364102
rect 204448 363978 204768 364046
rect 204448 363922 204518 363978
rect 204574 363922 204642 363978
rect 204698 363922 204768 363978
rect 204448 363888 204768 363922
rect 235168 364350 235488 364384
rect 235168 364294 235238 364350
rect 235294 364294 235362 364350
rect 235418 364294 235488 364350
rect 235168 364226 235488 364294
rect 235168 364170 235238 364226
rect 235294 364170 235362 364226
rect 235418 364170 235488 364226
rect 235168 364102 235488 364170
rect 235168 364046 235238 364102
rect 235294 364046 235362 364102
rect 235418 364046 235488 364102
rect 235168 363978 235488 364046
rect 235168 363922 235238 363978
rect 235294 363922 235362 363978
rect 235418 363922 235488 363978
rect 235168 363888 235488 363922
rect 265888 364350 266208 364384
rect 265888 364294 265958 364350
rect 266014 364294 266082 364350
rect 266138 364294 266208 364350
rect 265888 364226 266208 364294
rect 265888 364170 265958 364226
rect 266014 364170 266082 364226
rect 266138 364170 266208 364226
rect 265888 364102 266208 364170
rect 265888 364046 265958 364102
rect 266014 364046 266082 364102
rect 266138 364046 266208 364102
rect 265888 363978 266208 364046
rect 265888 363922 265958 363978
rect 266014 363922 266082 363978
rect 266138 363922 266208 363978
rect 265888 363888 266208 363922
rect 296608 364350 296928 364384
rect 296608 364294 296678 364350
rect 296734 364294 296802 364350
rect 296858 364294 296928 364350
rect 296608 364226 296928 364294
rect 296608 364170 296678 364226
rect 296734 364170 296802 364226
rect 296858 364170 296928 364226
rect 296608 364102 296928 364170
rect 296608 364046 296678 364102
rect 296734 364046 296802 364102
rect 296858 364046 296928 364102
rect 296608 363978 296928 364046
rect 296608 363922 296678 363978
rect 296734 363922 296802 363978
rect 296858 363922 296928 363978
rect 296608 363888 296928 363922
rect 327328 364350 327648 364384
rect 327328 364294 327398 364350
rect 327454 364294 327522 364350
rect 327578 364294 327648 364350
rect 327328 364226 327648 364294
rect 327328 364170 327398 364226
rect 327454 364170 327522 364226
rect 327578 364170 327648 364226
rect 327328 364102 327648 364170
rect 327328 364046 327398 364102
rect 327454 364046 327522 364102
rect 327578 364046 327648 364102
rect 327328 363978 327648 364046
rect 327328 363922 327398 363978
rect 327454 363922 327522 363978
rect 327578 363922 327648 363978
rect 327328 363888 327648 363922
rect 358048 364350 358368 364384
rect 358048 364294 358118 364350
rect 358174 364294 358242 364350
rect 358298 364294 358368 364350
rect 358048 364226 358368 364294
rect 358048 364170 358118 364226
rect 358174 364170 358242 364226
rect 358298 364170 358368 364226
rect 358048 364102 358368 364170
rect 358048 364046 358118 364102
rect 358174 364046 358242 364102
rect 358298 364046 358368 364102
rect 358048 363978 358368 364046
rect 358048 363922 358118 363978
rect 358174 363922 358242 363978
rect 358298 363922 358368 363978
rect 358048 363888 358368 363922
rect 388768 364350 389088 364384
rect 388768 364294 388838 364350
rect 388894 364294 388962 364350
rect 389018 364294 389088 364350
rect 388768 364226 389088 364294
rect 388768 364170 388838 364226
rect 388894 364170 388962 364226
rect 389018 364170 389088 364226
rect 388768 364102 389088 364170
rect 388768 364046 388838 364102
rect 388894 364046 388962 364102
rect 389018 364046 389088 364102
rect 388768 363978 389088 364046
rect 388768 363922 388838 363978
rect 388894 363922 388962 363978
rect 389018 363922 389088 363978
rect 388768 363888 389088 363922
rect 419488 364350 419808 364384
rect 419488 364294 419558 364350
rect 419614 364294 419682 364350
rect 419738 364294 419808 364350
rect 419488 364226 419808 364294
rect 419488 364170 419558 364226
rect 419614 364170 419682 364226
rect 419738 364170 419808 364226
rect 419488 364102 419808 364170
rect 419488 364046 419558 364102
rect 419614 364046 419682 364102
rect 419738 364046 419808 364102
rect 419488 363978 419808 364046
rect 419488 363922 419558 363978
rect 419614 363922 419682 363978
rect 419738 363922 419808 363978
rect 419488 363888 419808 363922
rect 450208 364350 450528 364384
rect 450208 364294 450278 364350
rect 450334 364294 450402 364350
rect 450458 364294 450528 364350
rect 450208 364226 450528 364294
rect 450208 364170 450278 364226
rect 450334 364170 450402 364226
rect 450458 364170 450528 364226
rect 450208 364102 450528 364170
rect 450208 364046 450278 364102
rect 450334 364046 450402 364102
rect 450458 364046 450528 364102
rect 450208 363978 450528 364046
rect 450208 363922 450278 363978
rect 450334 363922 450402 363978
rect 450458 363922 450528 363978
rect 450208 363888 450528 363922
rect 480928 364350 481248 364384
rect 480928 364294 480998 364350
rect 481054 364294 481122 364350
rect 481178 364294 481248 364350
rect 480928 364226 481248 364294
rect 480928 364170 480998 364226
rect 481054 364170 481122 364226
rect 481178 364170 481248 364226
rect 480928 364102 481248 364170
rect 480928 364046 480998 364102
rect 481054 364046 481122 364102
rect 481178 364046 481248 364102
rect 480928 363978 481248 364046
rect 480928 363922 480998 363978
rect 481054 363922 481122 363978
rect 481178 363922 481248 363978
rect 480928 363888 481248 363922
rect 507154 364350 507774 381922
rect 507154 364294 507250 364350
rect 507306 364294 507374 364350
rect 507430 364294 507498 364350
rect 507554 364294 507622 364350
rect 507678 364294 507774 364350
rect 507154 364226 507774 364294
rect 507154 364170 507250 364226
rect 507306 364170 507374 364226
rect 507430 364170 507498 364226
rect 507554 364170 507622 364226
rect 507678 364170 507774 364226
rect 507154 364102 507774 364170
rect 507154 364046 507250 364102
rect 507306 364046 507374 364102
rect 507430 364046 507498 364102
rect 507554 364046 507622 364102
rect 507678 364046 507774 364102
rect 507154 363978 507774 364046
rect 507154 363922 507250 363978
rect 507306 363922 507374 363978
rect 507430 363922 507498 363978
rect 507554 363922 507622 363978
rect 507678 363922 507774 363978
rect 219808 352350 220128 352384
rect 219808 352294 219878 352350
rect 219934 352294 220002 352350
rect 220058 352294 220128 352350
rect 219808 352226 220128 352294
rect 219808 352170 219878 352226
rect 219934 352170 220002 352226
rect 220058 352170 220128 352226
rect 219808 352102 220128 352170
rect 219808 352046 219878 352102
rect 219934 352046 220002 352102
rect 220058 352046 220128 352102
rect 219808 351978 220128 352046
rect 219808 351922 219878 351978
rect 219934 351922 220002 351978
rect 220058 351922 220128 351978
rect 219808 351888 220128 351922
rect 250528 352350 250848 352384
rect 250528 352294 250598 352350
rect 250654 352294 250722 352350
rect 250778 352294 250848 352350
rect 250528 352226 250848 352294
rect 250528 352170 250598 352226
rect 250654 352170 250722 352226
rect 250778 352170 250848 352226
rect 250528 352102 250848 352170
rect 250528 352046 250598 352102
rect 250654 352046 250722 352102
rect 250778 352046 250848 352102
rect 250528 351978 250848 352046
rect 250528 351922 250598 351978
rect 250654 351922 250722 351978
rect 250778 351922 250848 351978
rect 250528 351888 250848 351922
rect 281248 352350 281568 352384
rect 281248 352294 281318 352350
rect 281374 352294 281442 352350
rect 281498 352294 281568 352350
rect 281248 352226 281568 352294
rect 281248 352170 281318 352226
rect 281374 352170 281442 352226
rect 281498 352170 281568 352226
rect 281248 352102 281568 352170
rect 281248 352046 281318 352102
rect 281374 352046 281442 352102
rect 281498 352046 281568 352102
rect 281248 351978 281568 352046
rect 281248 351922 281318 351978
rect 281374 351922 281442 351978
rect 281498 351922 281568 351978
rect 281248 351888 281568 351922
rect 311968 352350 312288 352384
rect 311968 352294 312038 352350
rect 312094 352294 312162 352350
rect 312218 352294 312288 352350
rect 311968 352226 312288 352294
rect 311968 352170 312038 352226
rect 312094 352170 312162 352226
rect 312218 352170 312288 352226
rect 311968 352102 312288 352170
rect 311968 352046 312038 352102
rect 312094 352046 312162 352102
rect 312218 352046 312288 352102
rect 311968 351978 312288 352046
rect 311968 351922 312038 351978
rect 312094 351922 312162 351978
rect 312218 351922 312288 351978
rect 311968 351888 312288 351922
rect 342688 352350 343008 352384
rect 342688 352294 342758 352350
rect 342814 352294 342882 352350
rect 342938 352294 343008 352350
rect 342688 352226 343008 352294
rect 342688 352170 342758 352226
rect 342814 352170 342882 352226
rect 342938 352170 343008 352226
rect 342688 352102 343008 352170
rect 342688 352046 342758 352102
rect 342814 352046 342882 352102
rect 342938 352046 343008 352102
rect 342688 351978 343008 352046
rect 342688 351922 342758 351978
rect 342814 351922 342882 351978
rect 342938 351922 343008 351978
rect 342688 351888 343008 351922
rect 373408 352350 373728 352384
rect 373408 352294 373478 352350
rect 373534 352294 373602 352350
rect 373658 352294 373728 352350
rect 373408 352226 373728 352294
rect 373408 352170 373478 352226
rect 373534 352170 373602 352226
rect 373658 352170 373728 352226
rect 373408 352102 373728 352170
rect 373408 352046 373478 352102
rect 373534 352046 373602 352102
rect 373658 352046 373728 352102
rect 373408 351978 373728 352046
rect 373408 351922 373478 351978
rect 373534 351922 373602 351978
rect 373658 351922 373728 351978
rect 373408 351888 373728 351922
rect 404128 352350 404448 352384
rect 404128 352294 404198 352350
rect 404254 352294 404322 352350
rect 404378 352294 404448 352350
rect 404128 352226 404448 352294
rect 404128 352170 404198 352226
rect 404254 352170 404322 352226
rect 404378 352170 404448 352226
rect 404128 352102 404448 352170
rect 404128 352046 404198 352102
rect 404254 352046 404322 352102
rect 404378 352046 404448 352102
rect 404128 351978 404448 352046
rect 404128 351922 404198 351978
rect 404254 351922 404322 351978
rect 404378 351922 404448 351978
rect 404128 351888 404448 351922
rect 434848 352350 435168 352384
rect 434848 352294 434918 352350
rect 434974 352294 435042 352350
rect 435098 352294 435168 352350
rect 434848 352226 435168 352294
rect 434848 352170 434918 352226
rect 434974 352170 435042 352226
rect 435098 352170 435168 352226
rect 434848 352102 435168 352170
rect 434848 352046 434918 352102
rect 434974 352046 435042 352102
rect 435098 352046 435168 352102
rect 434848 351978 435168 352046
rect 434848 351922 434918 351978
rect 434974 351922 435042 351978
rect 435098 351922 435168 351978
rect 434848 351888 435168 351922
rect 465568 352350 465888 352384
rect 465568 352294 465638 352350
rect 465694 352294 465762 352350
rect 465818 352294 465888 352350
rect 465568 352226 465888 352294
rect 465568 352170 465638 352226
rect 465694 352170 465762 352226
rect 465818 352170 465888 352226
rect 465568 352102 465888 352170
rect 465568 352046 465638 352102
rect 465694 352046 465762 352102
rect 465818 352046 465888 352102
rect 465568 351978 465888 352046
rect 465568 351922 465638 351978
rect 465694 351922 465762 351978
rect 465818 351922 465888 351978
rect 465568 351888 465888 351922
rect 496288 352350 496608 352384
rect 496288 352294 496358 352350
rect 496414 352294 496482 352350
rect 496538 352294 496608 352350
rect 496288 352226 496608 352294
rect 496288 352170 496358 352226
rect 496414 352170 496482 352226
rect 496538 352170 496608 352226
rect 496288 352102 496608 352170
rect 496288 352046 496358 352102
rect 496414 352046 496482 352102
rect 496538 352046 496608 352102
rect 496288 351978 496608 352046
rect 496288 351922 496358 351978
rect 496414 351922 496482 351978
rect 496538 351922 496608 351978
rect 496288 351888 496608 351922
rect 201154 346294 201250 346350
rect 201306 346294 201374 346350
rect 201430 346294 201498 346350
rect 201554 346294 201622 346350
rect 201678 346294 201774 346350
rect 201154 346226 201774 346294
rect 201154 346170 201250 346226
rect 201306 346170 201374 346226
rect 201430 346170 201498 346226
rect 201554 346170 201622 346226
rect 201678 346170 201774 346226
rect 201154 346102 201774 346170
rect 201154 346046 201250 346102
rect 201306 346046 201374 346102
rect 201430 346046 201498 346102
rect 201554 346046 201622 346102
rect 201678 346046 201774 346102
rect 201154 345978 201774 346046
rect 201154 345922 201250 345978
rect 201306 345922 201374 345978
rect 201430 345922 201498 345978
rect 201554 345922 201622 345978
rect 201678 345922 201774 345978
rect 201154 328350 201774 345922
rect 204448 346350 204768 346384
rect 204448 346294 204518 346350
rect 204574 346294 204642 346350
rect 204698 346294 204768 346350
rect 204448 346226 204768 346294
rect 204448 346170 204518 346226
rect 204574 346170 204642 346226
rect 204698 346170 204768 346226
rect 204448 346102 204768 346170
rect 204448 346046 204518 346102
rect 204574 346046 204642 346102
rect 204698 346046 204768 346102
rect 204448 345978 204768 346046
rect 204448 345922 204518 345978
rect 204574 345922 204642 345978
rect 204698 345922 204768 345978
rect 204448 345888 204768 345922
rect 235168 346350 235488 346384
rect 235168 346294 235238 346350
rect 235294 346294 235362 346350
rect 235418 346294 235488 346350
rect 235168 346226 235488 346294
rect 235168 346170 235238 346226
rect 235294 346170 235362 346226
rect 235418 346170 235488 346226
rect 235168 346102 235488 346170
rect 235168 346046 235238 346102
rect 235294 346046 235362 346102
rect 235418 346046 235488 346102
rect 235168 345978 235488 346046
rect 235168 345922 235238 345978
rect 235294 345922 235362 345978
rect 235418 345922 235488 345978
rect 235168 345888 235488 345922
rect 265888 346350 266208 346384
rect 265888 346294 265958 346350
rect 266014 346294 266082 346350
rect 266138 346294 266208 346350
rect 265888 346226 266208 346294
rect 265888 346170 265958 346226
rect 266014 346170 266082 346226
rect 266138 346170 266208 346226
rect 265888 346102 266208 346170
rect 265888 346046 265958 346102
rect 266014 346046 266082 346102
rect 266138 346046 266208 346102
rect 265888 345978 266208 346046
rect 265888 345922 265958 345978
rect 266014 345922 266082 345978
rect 266138 345922 266208 345978
rect 265888 345888 266208 345922
rect 296608 346350 296928 346384
rect 296608 346294 296678 346350
rect 296734 346294 296802 346350
rect 296858 346294 296928 346350
rect 296608 346226 296928 346294
rect 296608 346170 296678 346226
rect 296734 346170 296802 346226
rect 296858 346170 296928 346226
rect 296608 346102 296928 346170
rect 296608 346046 296678 346102
rect 296734 346046 296802 346102
rect 296858 346046 296928 346102
rect 296608 345978 296928 346046
rect 296608 345922 296678 345978
rect 296734 345922 296802 345978
rect 296858 345922 296928 345978
rect 296608 345888 296928 345922
rect 327328 346350 327648 346384
rect 327328 346294 327398 346350
rect 327454 346294 327522 346350
rect 327578 346294 327648 346350
rect 327328 346226 327648 346294
rect 327328 346170 327398 346226
rect 327454 346170 327522 346226
rect 327578 346170 327648 346226
rect 327328 346102 327648 346170
rect 327328 346046 327398 346102
rect 327454 346046 327522 346102
rect 327578 346046 327648 346102
rect 327328 345978 327648 346046
rect 327328 345922 327398 345978
rect 327454 345922 327522 345978
rect 327578 345922 327648 345978
rect 327328 345888 327648 345922
rect 358048 346350 358368 346384
rect 358048 346294 358118 346350
rect 358174 346294 358242 346350
rect 358298 346294 358368 346350
rect 358048 346226 358368 346294
rect 358048 346170 358118 346226
rect 358174 346170 358242 346226
rect 358298 346170 358368 346226
rect 358048 346102 358368 346170
rect 358048 346046 358118 346102
rect 358174 346046 358242 346102
rect 358298 346046 358368 346102
rect 358048 345978 358368 346046
rect 358048 345922 358118 345978
rect 358174 345922 358242 345978
rect 358298 345922 358368 345978
rect 358048 345888 358368 345922
rect 388768 346350 389088 346384
rect 388768 346294 388838 346350
rect 388894 346294 388962 346350
rect 389018 346294 389088 346350
rect 388768 346226 389088 346294
rect 388768 346170 388838 346226
rect 388894 346170 388962 346226
rect 389018 346170 389088 346226
rect 388768 346102 389088 346170
rect 388768 346046 388838 346102
rect 388894 346046 388962 346102
rect 389018 346046 389088 346102
rect 388768 345978 389088 346046
rect 388768 345922 388838 345978
rect 388894 345922 388962 345978
rect 389018 345922 389088 345978
rect 388768 345888 389088 345922
rect 419488 346350 419808 346384
rect 419488 346294 419558 346350
rect 419614 346294 419682 346350
rect 419738 346294 419808 346350
rect 419488 346226 419808 346294
rect 419488 346170 419558 346226
rect 419614 346170 419682 346226
rect 419738 346170 419808 346226
rect 419488 346102 419808 346170
rect 419488 346046 419558 346102
rect 419614 346046 419682 346102
rect 419738 346046 419808 346102
rect 419488 345978 419808 346046
rect 419488 345922 419558 345978
rect 419614 345922 419682 345978
rect 419738 345922 419808 345978
rect 419488 345888 419808 345922
rect 450208 346350 450528 346384
rect 450208 346294 450278 346350
rect 450334 346294 450402 346350
rect 450458 346294 450528 346350
rect 450208 346226 450528 346294
rect 450208 346170 450278 346226
rect 450334 346170 450402 346226
rect 450458 346170 450528 346226
rect 450208 346102 450528 346170
rect 450208 346046 450278 346102
rect 450334 346046 450402 346102
rect 450458 346046 450528 346102
rect 450208 345978 450528 346046
rect 450208 345922 450278 345978
rect 450334 345922 450402 345978
rect 450458 345922 450528 345978
rect 450208 345888 450528 345922
rect 480928 346350 481248 346384
rect 480928 346294 480998 346350
rect 481054 346294 481122 346350
rect 481178 346294 481248 346350
rect 480928 346226 481248 346294
rect 480928 346170 480998 346226
rect 481054 346170 481122 346226
rect 481178 346170 481248 346226
rect 480928 346102 481248 346170
rect 480928 346046 480998 346102
rect 481054 346046 481122 346102
rect 481178 346046 481248 346102
rect 480928 345978 481248 346046
rect 480928 345922 480998 345978
rect 481054 345922 481122 345978
rect 481178 345922 481248 345978
rect 480928 345888 481248 345922
rect 507154 346350 507774 363922
rect 507154 346294 507250 346350
rect 507306 346294 507374 346350
rect 507430 346294 507498 346350
rect 507554 346294 507622 346350
rect 507678 346294 507774 346350
rect 507154 346226 507774 346294
rect 507154 346170 507250 346226
rect 507306 346170 507374 346226
rect 507430 346170 507498 346226
rect 507554 346170 507622 346226
rect 507678 346170 507774 346226
rect 507154 346102 507774 346170
rect 507154 346046 507250 346102
rect 507306 346046 507374 346102
rect 507430 346046 507498 346102
rect 507554 346046 507622 346102
rect 507678 346046 507774 346102
rect 507154 345978 507774 346046
rect 507154 345922 507250 345978
rect 507306 345922 507374 345978
rect 507430 345922 507498 345978
rect 507554 345922 507622 345978
rect 507678 345922 507774 345978
rect 219808 334350 220128 334384
rect 219808 334294 219878 334350
rect 219934 334294 220002 334350
rect 220058 334294 220128 334350
rect 219808 334226 220128 334294
rect 219808 334170 219878 334226
rect 219934 334170 220002 334226
rect 220058 334170 220128 334226
rect 219808 334102 220128 334170
rect 219808 334046 219878 334102
rect 219934 334046 220002 334102
rect 220058 334046 220128 334102
rect 219808 333978 220128 334046
rect 219808 333922 219878 333978
rect 219934 333922 220002 333978
rect 220058 333922 220128 333978
rect 219808 333888 220128 333922
rect 250528 334350 250848 334384
rect 250528 334294 250598 334350
rect 250654 334294 250722 334350
rect 250778 334294 250848 334350
rect 250528 334226 250848 334294
rect 250528 334170 250598 334226
rect 250654 334170 250722 334226
rect 250778 334170 250848 334226
rect 250528 334102 250848 334170
rect 250528 334046 250598 334102
rect 250654 334046 250722 334102
rect 250778 334046 250848 334102
rect 250528 333978 250848 334046
rect 250528 333922 250598 333978
rect 250654 333922 250722 333978
rect 250778 333922 250848 333978
rect 250528 333888 250848 333922
rect 281248 334350 281568 334384
rect 281248 334294 281318 334350
rect 281374 334294 281442 334350
rect 281498 334294 281568 334350
rect 281248 334226 281568 334294
rect 281248 334170 281318 334226
rect 281374 334170 281442 334226
rect 281498 334170 281568 334226
rect 281248 334102 281568 334170
rect 281248 334046 281318 334102
rect 281374 334046 281442 334102
rect 281498 334046 281568 334102
rect 281248 333978 281568 334046
rect 281248 333922 281318 333978
rect 281374 333922 281442 333978
rect 281498 333922 281568 333978
rect 281248 333888 281568 333922
rect 311968 334350 312288 334384
rect 311968 334294 312038 334350
rect 312094 334294 312162 334350
rect 312218 334294 312288 334350
rect 311968 334226 312288 334294
rect 311968 334170 312038 334226
rect 312094 334170 312162 334226
rect 312218 334170 312288 334226
rect 311968 334102 312288 334170
rect 311968 334046 312038 334102
rect 312094 334046 312162 334102
rect 312218 334046 312288 334102
rect 311968 333978 312288 334046
rect 311968 333922 312038 333978
rect 312094 333922 312162 333978
rect 312218 333922 312288 333978
rect 311968 333888 312288 333922
rect 342688 334350 343008 334384
rect 342688 334294 342758 334350
rect 342814 334294 342882 334350
rect 342938 334294 343008 334350
rect 342688 334226 343008 334294
rect 342688 334170 342758 334226
rect 342814 334170 342882 334226
rect 342938 334170 343008 334226
rect 342688 334102 343008 334170
rect 342688 334046 342758 334102
rect 342814 334046 342882 334102
rect 342938 334046 343008 334102
rect 342688 333978 343008 334046
rect 342688 333922 342758 333978
rect 342814 333922 342882 333978
rect 342938 333922 343008 333978
rect 342688 333888 343008 333922
rect 373408 334350 373728 334384
rect 373408 334294 373478 334350
rect 373534 334294 373602 334350
rect 373658 334294 373728 334350
rect 373408 334226 373728 334294
rect 373408 334170 373478 334226
rect 373534 334170 373602 334226
rect 373658 334170 373728 334226
rect 373408 334102 373728 334170
rect 373408 334046 373478 334102
rect 373534 334046 373602 334102
rect 373658 334046 373728 334102
rect 373408 333978 373728 334046
rect 373408 333922 373478 333978
rect 373534 333922 373602 333978
rect 373658 333922 373728 333978
rect 373408 333888 373728 333922
rect 404128 334350 404448 334384
rect 404128 334294 404198 334350
rect 404254 334294 404322 334350
rect 404378 334294 404448 334350
rect 404128 334226 404448 334294
rect 404128 334170 404198 334226
rect 404254 334170 404322 334226
rect 404378 334170 404448 334226
rect 404128 334102 404448 334170
rect 404128 334046 404198 334102
rect 404254 334046 404322 334102
rect 404378 334046 404448 334102
rect 404128 333978 404448 334046
rect 404128 333922 404198 333978
rect 404254 333922 404322 333978
rect 404378 333922 404448 333978
rect 404128 333888 404448 333922
rect 434848 334350 435168 334384
rect 434848 334294 434918 334350
rect 434974 334294 435042 334350
rect 435098 334294 435168 334350
rect 434848 334226 435168 334294
rect 434848 334170 434918 334226
rect 434974 334170 435042 334226
rect 435098 334170 435168 334226
rect 434848 334102 435168 334170
rect 434848 334046 434918 334102
rect 434974 334046 435042 334102
rect 435098 334046 435168 334102
rect 434848 333978 435168 334046
rect 434848 333922 434918 333978
rect 434974 333922 435042 333978
rect 435098 333922 435168 333978
rect 434848 333888 435168 333922
rect 465568 334350 465888 334384
rect 465568 334294 465638 334350
rect 465694 334294 465762 334350
rect 465818 334294 465888 334350
rect 465568 334226 465888 334294
rect 465568 334170 465638 334226
rect 465694 334170 465762 334226
rect 465818 334170 465888 334226
rect 465568 334102 465888 334170
rect 465568 334046 465638 334102
rect 465694 334046 465762 334102
rect 465818 334046 465888 334102
rect 465568 333978 465888 334046
rect 465568 333922 465638 333978
rect 465694 333922 465762 333978
rect 465818 333922 465888 333978
rect 465568 333888 465888 333922
rect 496288 334350 496608 334384
rect 496288 334294 496358 334350
rect 496414 334294 496482 334350
rect 496538 334294 496608 334350
rect 496288 334226 496608 334294
rect 496288 334170 496358 334226
rect 496414 334170 496482 334226
rect 496538 334170 496608 334226
rect 496288 334102 496608 334170
rect 496288 334046 496358 334102
rect 496414 334046 496482 334102
rect 496538 334046 496608 334102
rect 496288 333978 496608 334046
rect 496288 333922 496358 333978
rect 496414 333922 496482 333978
rect 496538 333922 496608 333978
rect 496288 333888 496608 333922
rect 201154 328294 201250 328350
rect 201306 328294 201374 328350
rect 201430 328294 201498 328350
rect 201554 328294 201622 328350
rect 201678 328294 201774 328350
rect 201154 328226 201774 328294
rect 201154 328170 201250 328226
rect 201306 328170 201374 328226
rect 201430 328170 201498 328226
rect 201554 328170 201622 328226
rect 201678 328170 201774 328226
rect 201154 328102 201774 328170
rect 201154 328046 201250 328102
rect 201306 328046 201374 328102
rect 201430 328046 201498 328102
rect 201554 328046 201622 328102
rect 201678 328046 201774 328102
rect 201154 327978 201774 328046
rect 201154 327922 201250 327978
rect 201306 327922 201374 327978
rect 201430 327922 201498 327978
rect 201554 327922 201622 327978
rect 201678 327922 201774 327978
rect 201154 310350 201774 327922
rect 204448 328350 204768 328384
rect 204448 328294 204518 328350
rect 204574 328294 204642 328350
rect 204698 328294 204768 328350
rect 204448 328226 204768 328294
rect 204448 328170 204518 328226
rect 204574 328170 204642 328226
rect 204698 328170 204768 328226
rect 204448 328102 204768 328170
rect 204448 328046 204518 328102
rect 204574 328046 204642 328102
rect 204698 328046 204768 328102
rect 204448 327978 204768 328046
rect 204448 327922 204518 327978
rect 204574 327922 204642 327978
rect 204698 327922 204768 327978
rect 204448 327888 204768 327922
rect 235168 328350 235488 328384
rect 235168 328294 235238 328350
rect 235294 328294 235362 328350
rect 235418 328294 235488 328350
rect 235168 328226 235488 328294
rect 235168 328170 235238 328226
rect 235294 328170 235362 328226
rect 235418 328170 235488 328226
rect 235168 328102 235488 328170
rect 235168 328046 235238 328102
rect 235294 328046 235362 328102
rect 235418 328046 235488 328102
rect 235168 327978 235488 328046
rect 235168 327922 235238 327978
rect 235294 327922 235362 327978
rect 235418 327922 235488 327978
rect 235168 327888 235488 327922
rect 265888 328350 266208 328384
rect 265888 328294 265958 328350
rect 266014 328294 266082 328350
rect 266138 328294 266208 328350
rect 265888 328226 266208 328294
rect 265888 328170 265958 328226
rect 266014 328170 266082 328226
rect 266138 328170 266208 328226
rect 265888 328102 266208 328170
rect 265888 328046 265958 328102
rect 266014 328046 266082 328102
rect 266138 328046 266208 328102
rect 265888 327978 266208 328046
rect 265888 327922 265958 327978
rect 266014 327922 266082 327978
rect 266138 327922 266208 327978
rect 265888 327888 266208 327922
rect 296608 328350 296928 328384
rect 296608 328294 296678 328350
rect 296734 328294 296802 328350
rect 296858 328294 296928 328350
rect 296608 328226 296928 328294
rect 296608 328170 296678 328226
rect 296734 328170 296802 328226
rect 296858 328170 296928 328226
rect 296608 328102 296928 328170
rect 296608 328046 296678 328102
rect 296734 328046 296802 328102
rect 296858 328046 296928 328102
rect 296608 327978 296928 328046
rect 296608 327922 296678 327978
rect 296734 327922 296802 327978
rect 296858 327922 296928 327978
rect 296608 327888 296928 327922
rect 327328 328350 327648 328384
rect 327328 328294 327398 328350
rect 327454 328294 327522 328350
rect 327578 328294 327648 328350
rect 327328 328226 327648 328294
rect 327328 328170 327398 328226
rect 327454 328170 327522 328226
rect 327578 328170 327648 328226
rect 327328 328102 327648 328170
rect 327328 328046 327398 328102
rect 327454 328046 327522 328102
rect 327578 328046 327648 328102
rect 327328 327978 327648 328046
rect 327328 327922 327398 327978
rect 327454 327922 327522 327978
rect 327578 327922 327648 327978
rect 327328 327888 327648 327922
rect 358048 328350 358368 328384
rect 358048 328294 358118 328350
rect 358174 328294 358242 328350
rect 358298 328294 358368 328350
rect 358048 328226 358368 328294
rect 358048 328170 358118 328226
rect 358174 328170 358242 328226
rect 358298 328170 358368 328226
rect 358048 328102 358368 328170
rect 358048 328046 358118 328102
rect 358174 328046 358242 328102
rect 358298 328046 358368 328102
rect 358048 327978 358368 328046
rect 358048 327922 358118 327978
rect 358174 327922 358242 327978
rect 358298 327922 358368 327978
rect 358048 327888 358368 327922
rect 388768 328350 389088 328384
rect 388768 328294 388838 328350
rect 388894 328294 388962 328350
rect 389018 328294 389088 328350
rect 388768 328226 389088 328294
rect 388768 328170 388838 328226
rect 388894 328170 388962 328226
rect 389018 328170 389088 328226
rect 388768 328102 389088 328170
rect 388768 328046 388838 328102
rect 388894 328046 388962 328102
rect 389018 328046 389088 328102
rect 388768 327978 389088 328046
rect 388768 327922 388838 327978
rect 388894 327922 388962 327978
rect 389018 327922 389088 327978
rect 388768 327888 389088 327922
rect 419488 328350 419808 328384
rect 419488 328294 419558 328350
rect 419614 328294 419682 328350
rect 419738 328294 419808 328350
rect 419488 328226 419808 328294
rect 419488 328170 419558 328226
rect 419614 328170 419682 328226
rect 419738 328170 419808 328226
rect 419488 328102 419808 328170
rect 419488 328046 419558 328102
rect 419614 328046 419682 328102
rect 419738 328046 419808 328102
rect 419488 327978 419808 328046
rect 419488 327922 419558 327978
rect 419614 327922 419682 327978
rect 419738 327922 419808 327978
rect 419488 327888 419808 327922
rect 450208 328350 450528 328384
rect 450208 328294 450278 328350
rect 450334 328294 450402 328350
rect 450458 328294 450528 328350
rect 450208 328226 450528 328294
rect 450208 328170 450278 328226
rect 450334 328170 450402 328226
rect 450458 328170 450528 328226
rect 450208 328102 450528 328170
rect 450208 328046 450278 328102
rect 450334 328046 450402 328102
rect 450458 328046 450528 328102
rect 450208 327978 450528 328046
rect 450208 327922 450278 327978
rect 450334 327922 450402 327978
rect 450458 327922 450528 327978
rect 450208 327888 450528 327922
rect 480928 328350 481248 328384
rect 480928 328294 480998 328350
rect 481054 328294 481122 328350
rect 481178 328294 481248 328350
rect 480928 328226 481248 328294
rect 480928 328170 480998 328226
rect 481054 328170 481122 328226
rect 481178 328170 481248 328226
rect 480928 328102 481248 328170
rect 480928 328046 480998 328102
rect 481054 328046 481122 328102
rect 481178 328046 481248 328102
rect 480928 327978 481248 328046
rect 480928 327922 480998 327978
rect 481054 327922 481122 327978
rect 481178 327922 481248 327978
rect 480928 327888 481248 327922
rect 507154 328350 507774 345922
rect 507154 328294 507250 328350
rect 507306 328294 507374 328350
rect 507430 328294 507498 328350
rect 507554 328294 507622 328350
rect 507678 328294 507774 328350
rect 507154 328226 507774 328294
rect 507154 328170 507250 328226
rect 507306 328170 507374 328226
rect 507430 328170 507498 328226
rect 507554 328170 507622 328226
rect 507678 328170 507774 328226
rect 507154 328102 507774 328170
rect 507154 328046 507250 328102
rect 507306 328046 507374 328102
rect 507430 328046 507498 328102
rect 507554 328046 507622 328102
rect 507678 328046 507774 328102
rect 507154 327978 507774 328046
rect 507154 327922 507250 327978
rect 507306 327922 507374 327978
rect 507430 327922 507498 327978
rect 507554 327922 507622 327978
rect 507678 327922 507774 327978
rect 219808 316350 220128 316384
rect 219808 316294 219878 316350
rect 219934 316294 220002 316350
rect 220058 316294 220128 316350
rect 219808 316226 220128 316294
rect 219808 316170 219878 316226
rect 219934 316170 220002 316226
rect 220058 316170 220128 316226
rect 219808 316102 220128 316170
rect 219808 316046 219878 316102
rect 219934 316046 220002 316102
rect 220058 316046 220128 316102
rect 219808 315978 220128 316046
rect 219808 315922 219878 315978
rect 219934 315922 220002 315978
rect 220058 315922 220128 315978
rect 219808 315888 220128 315922
rect 250528 316350 250848 316384
rect 250528 316294 250598 316350
rect 250654 316294 250722 316350
rect 250778 316294 250848 316350
rect 250528 316226 250848 316294
rect 250528 316170 250598 316226
rect 250654 316170 250722 316226
rect 250778 316170 250848 316226
rect 250528 316102 250848 316170
rect 250528 316046 250598 316102
rect 250654 316046 250722 316102
rect 250778 316046 250848 316102
rect 250528 315978 250848 316046
rect 250528 315922 250598 315978
rect 250654 315922 250722 315978
rect 250778 315922 250848 315978
rect 250528 315888 250848 315922
rect 281248 316350 281568 316384
rect 281248 316294 281318 316350
rect 281374 316294 281442 316350
rect 281498 316294 281568 316350
rect 281248 316226 281568 316294
rect 281248 316170 281318 316226
rect 281374 316170 281442 316226
rect 281498 316170 281568 316226
rect 281248 316102 281568 316170
rect 281248 316046 281318 316102
rect 281374 316046 281442 316102
rect 281498 316046 281568 316102
rect 281248 315978 281568 316046
rect 281248 315922 281318 315978
rect 281374 315922 281442 315978
rect 281498 315922 281568 315978
rect 281248 315888 281568 315922
rect 311968 316350 312288 316384
rect 311968 316294 312038 316350
rect 312094 316294 312162 316350
rect 312218 316294 312288 316350
rect 311968 316226 312288 316294
rect 311968 316170 312038 316226
rect 312094 316170 312162 316226
rect 312218 316170 312288 316226
rect 311968 316102 312288 316170
rect 311968 316046 312038 316102
rect 312094 316046 312162 316102
rect 312218 316046 312288 316102
rect 311968 315978 312288 316046
rect 311968 315922 312038 315978
rect 312094 315922 312162 315978
rect 312218 315922 312288 315978
rect 311968 315888 312288 315922
rect 342688 316350 343008 316384
rect 342688 316294 342758 316350
rect 342814 316294 342882 316350
rect 342938 316294 343008 316350
rect 342688 316226 343008 316294
rect 342688 316170 342758 316226
rect 342814 316170 342882 316226
rect 342938 316170 343008 316226
rect 342688 316102 343008 316170
rect 342688 316046 342758 316102
rect 342814 316046 342882 316102
rect 342938 316046 343008 316102
rect 342688 315978 343008 316046
rect 342688 315922 342758 315978
rect 342814 315922 342882 315978
rect 342938 315922 343008 315978
rect 342688 315888 343008 315922
rect 373408 316350 373728 316384
rect 373408 316294 373478 316350
rect 373534 316294 373602 316350
rect 373658 316294 373728 316350
rect 373408 316226 373728 316294
rect 373408 316170 373478 316226
rect 373534 316170 373602 316226
rect 373658 316170 373728 316226
rect 373408 316102 373728 316170
rect 373408 316046 373478 316102
rect 373534 316046 373602 316102
rect 373658 316046 373728 316102
rect 373408 315978 373728 316046
rect 373408 315922 373478 315978
rect 373534 315922 373602 315978
rect 373658 315922 373728 315978
rect 373408 315888 373728 315922
rect 404128 316350 404448 316384
rect 404128 316294 404198 316350
rect 404254 316294 404322 316350
rect 404378 316294 404448 316350
rect 404128 316226 404448 316294
rect 404128 316170 404198 316226
rect 404254 316170 404322 316226
rect 404378 316170 404448 316226
rect 404128 316102 404448 316170
rect 404128 316046 404198 316102
rect 404254 316046 404322 316102
rect 404378 316046 404448 316102
rect 404128 315978 404448 316046
rect 404128 315922 404198 315978
rect 404254 315922 404322 315978
rect 404378 315922 404448 315978
rect 404128 315888 404448 315922
rect 434848 316350 435168 316384
rect 434848 316294 434918 316350
rect 434974 316294 435042 316350
rect 435098 316294 435168 316350
rect 434848 316226 435168 316294
rect 434848 316170 434918 316226
rect 434974 316170 435042 316226
rect 435098 316170 435168 316226
rect 434848 316102 435168 316170
rect 434848 316046 434918 316102
rect 434974 316046 435042 316102
rect 435098 316046 435168 316102
rect 434848 315978 435168 316046
rect 434848 315922 434918 315978
rect 434974 315922 435042 315978
rect 435098 315922 435168 315978
rect 434848 315888 435168 315922
rect 465568 316350 465888 316384
rect 465568 316294 465638 316350
rect 465694 316294 465762 316350
rect 465818 316294 465888 316350
rect 465568 316226 465888 316294
rect 465568 316170 465638 316226
rect 465694 316170 465762 316226
rect 465818 316170 465888 316226
rect 465568 316102 465888 316170
rect 465568 316046 465638 316102
rect 465694 316046 465762 316102
rect 465818 316046 465888 316102
rect 465568 315978 465888 316046
rect 465568 315922 465638 315978
rect 465694 315922 465762 315978
rect 465818 315922 465888 315978
rect 465568 315888 465888 315922
rect 496288 316350 496608 316384
rect 496288 316294 496358 316350
rect 496414 316294 496482 316350
rect 496538 316294 496608 316350
rect 496288 316226 496608 316294
rect 496288 316170 496358 316226
rect 496414 316170 496482 316226
rect 496538 316170 496608 316226
rect 496288 316102 496608 316170
rect 496288 316046 496358 316102
rect 496414 316046 496482 316102
rect 496538 316046 496608 316102
rect 496288 315978 496608 316046
rect 496288 315922 496358 315978
rect 496414 315922 496482 315978
rect 496538 315922 496608 315978
rect 496288 315888 496608 315922
rect 201154 310294 201250 310350
rect 201306 310294 201374 310350
rect 201430 310294 201498 310350
rect 201554 310294 201622 310350
rect 201678 310294 201774 310350
rect 201154 310226 201774 310294
rect 201154 310170 201250 310226
rect 201306 310170 201374 310226
rect 201430 310170 201498 310226
rect 201554 310170 201622 310226
rect 201678 310170 201774 310226
rect 201154 310102 201774 310170
rect 201154 310046 201250 310102
rect 201306 310046 201374 310102
rect 201430 310046 201498 310102
rect 201554 310046 201622 310102
rect 201678 310046 201774 310102
rect 201154 309978 201774 310046
rect 201154 309922 201250 309978
rect 201306 309922 201374 309978
rect 201430 309922 201498 309978
rect 201554 309922 201622 309978
rect 201678 309922 201774 309978
rect 201154 292350 201774 309922
rect 204448 310350 204768 310384
rect 204448 310294 204518 310350
rect 204574 310294 204642 310350
rect 204698 310294 204768 310350
rect 204448 310226 204768 310294
rect 204448 310170 204518 310226
rect 204574 310170 204642 310226
rect 204698 310170 204768 310226
rect 204448 310102 204768 310170
rect 204448 310046 204518 310102
rect 204574 310046 204642 310102
rect 204698 310046 204768 310102
rect 204448 309978 204768 310046
rect 204448 309922 204518 309978
rect 204574 309922 204642 309978
rect 204698 309922 204768 309978
rect 204448 309888 204768 309922
rect 235168 310350 235488 310384
rect 235168 310294 235238 310350
rect 235294 310294 235362 310350
rect 235418 310294 235488 310350
rect 235168 310226 235488 310294
rect 235168 310170 235238 310226
rect 235294 310170 235362 310226
rect 235418 310170 235488 310226
rect 235168 310102 235488 310170
rect 235168 310046 235238 310102
rect 235294 310046 235362 310102
rect 235418 310046 235488 310102
rect 235168 309978 235488 310046
rect 235168 309922 235238 309978
rect 235294 309922 235362 309978
rect 235418 309922 235488 309978
rect 235168 309888 235488 309922
rect 265888 310350 266208 310384
rect 265888 310294 265958 310350
rect 266014 310294 266082 310350
rect 266138 310294 266208 310350
rect 265888 310226 266208 310294
rect 265888 310170 265958 310226
rect 266014 310170 266082 310226
rect 266138 310170 266208 310226
rect 265888 310102 266208 310170
rect 265888 310046 265958 310102
rect 266014 310046 266082 310102
rect 266138 310046 266208 310102
rect 265888 309978 266208 310046
rect 265888 309922 265958 309978
rect 266014 309922 266082 309978
rect 266138 309922 266208 309978
rect 265888 309888 266208 309922
rect 296608 310350 296928 310384
rect 296608 310294 296678 310350
rect 296734 310294 296802 310350
rect 296858 310294 296928 310350
rect 296608 310226 296928 310294
rect 296608 310170 296678 310226
rect 296734 310170 296802 310226
rect 296858 310170 296928 310226
rect 296608 310102 296928 310170
rect 296608 310046 296678 310102
rect 296734 310046 296802 310102
rect 296858 310046 296928 310102
rect 296608 309978 296928 310046
rect 296608 309922 296678 309978
rect 296734 309922 296802 309978
rect 296858 309922 296928 309978
rect 296608 309888 296928 309922
rect 327328 310350 327648 310384
rect 327328 310294 327398 310350
rect 327454 310294 327522 310350
rect 327578 310294 327648 310350
rect 327328 310226 327648 310294
rect 327328 310170 327398 310226
rect 327454 310170 327522 310226
rect 327578 310170 327648 310226
rect 327328 310102 327648 310170
rect 327328 310046 327398 310102
rect 327454 310046 327522 310102
rect 327578 310046 327648 310102
rect 327328 309978 327648 310046
rect 327328 309922 327398 309978
rect 327454 309922 327522 309978
rect 327578 309922 327648 309978
rect 327328 309888 327648 309922
rect 358048 310350 358368 310384
rect 358048 310294 358118 310350
rect 358174 310294 358242 310350
rect 358298 310294 358368 310350
rect 358048 310226 358368 310294
rect 358048 310170 358118 310226
rect 358174 310170 358242 310226
rect 358298 310170 358368 310226
rect 358048 310102 358368 310170
rect 358048 310046 358118 310102
rect 358174 310046 358242 310102
rect 358298 310046 358368 310102
rect 358048 309978 358368 310046
rect 358048 309922 358118 309978
rect 358174 309922 358242 309978
rect 358298 309922 358368 309978
rect 358048 309888 358368 309922
rect 388768 310350 389088 310384
rect 388768 310294 388838 310350
rect 388894 310294 388962 310350
rect 389018 310294 389088 310350
rect 388768 310226 389088 310294
rect 388768 310170 388838 310226
rect 388894 310170 388962 310226
rect 389018 310170 389088 310226
rect 388768 310102 389088 310170
rect 388768 310046 388838 310102
rect 388894 310046 388962 310102
rect 389018 310046 389088 310102
rect 388768 309978 389088 310046
rect 388768 309922 388838 309978
rect 388894 309922 388962 309978
rect 389018 309922 389088 309978
rect 388768 309888 389088 309922
rect 419488 310350 419808 310384
rect 419488 310294 419558 310350
rect 419614 310294 419682 310350
rect 419738 310294 419808 310350
rect 419488 310226 419808 310294
rect 419488 310170 419558 310226
rect 419614 310170 419682 310226
rect 419738 310170 419808 310226
rect 419488 310102 419808 310170
rect 419488 310046 419558 310102
rect 419614 310046 419682 310102
rect 419738 310046 419808 310102
rect 419488 309978 419808 310046
rect 419488 309922 419558 309978
rect 419614 309922 419682 309978
rect 419738 309922 419808 309978
rect 419488 309888 419808 309922
rect 450208 310350 450528 310384
rect 450208 310294 450278 310350
rect 450334 310294 450402 310350
rect 450458 310294 450528 310350
rect 450208 310226 450528 310294
rect 450208 310170 450278 310226
rect 450334 310170 450402 310226
rect 450458 310170 450528 310226
rect 450208 310102 450528 310170
rect 450208 310046 450278 310102
rect 450334 310046 450402 310102
rect 450458 310046 450528 310102
rect 450208 309978 450528 310046
rect 450208 309922 450278 309978
rect 450334 309922 450402 309978
rect 450458 309922 450528 309978
rect 450208 309888 450528 309922
rect 480928 310350 481248 310384
rect 480928 310294 480998 310350
rect 481054 310294 481122 310350
rect 481178 310294 481248 310350
rect 480928 310226 481248 310294
rect 480928 310170 480998 310226
rect 481054 310170 481122 310226
rect 481178 310170 481248 310226
rect 480928 310102 481248 310170
rect 480928 310046 480998 310102
rect 481054 310046 481122 310102
rect 481178 310046 481248 310102
rect 480928 309978 481248 310046
rect 480928 309922 480998 309978
rect 481054 309922 481122 309978
rect 481178 309922 481248 309978
rect 480928 309888 481248 309922
rect 507154 310350 507774 327922
rect 507154 310294 507250 310350
rect 507306 310294 507374 310350
rect 507430 310294 507498 310350
rect 507554 310294 507622 310350
rect 507678 310294 507774 310350
rect 507154 310226 507774 310294
rect 507154 310170 507250 310226
rect 507306 310170 507374 310226
rect 507430 310170 507498 310226
rect 507554 310170 507622 310226
rect 507678 310170 507774 310226
rect 507154 310102 507774 310170
rect 507154 310046 507250 310102
rect 507306 310046 507374 310102
rect 507430 310046 507498 310102
rect 507554 310046 507622 310102
rect 507678 310046 507774 310102
rect 507154 309978 507774 310046
rect 507154 309922 507250 309978
rect 507306 309922 507374 309978
rect 507430 309922 507498 309978
rect 507554 309922 507622 309978
rect 507678 309922 507774 309978
rect 219808 298350 220128 298384
rect 219808 298294 219878 298350
rect 219934 298294 220002 298350
rect 220058 298294 220128 298350
rect 219808 298226 220128 298294
rect 219808 298170 219878 298226
rect 219934 298170 220002 298226
rect 220058 298170 220128 298226
rect 219808 298102 220128 298170
rect 219808 298046 219878 298102
rect 219934 298046 220002 298102
rect 220058 298046 220128 298102
rect 219808 297978 220128 298046
rect 219808 297922 219878 297978
rect 219934 297922 220002 297978
rect 220058 297922 220128 297978
rect 219808 297888 220128 297922
rect 250528 298350 250848 298384
rect 250528 298294 250598 298350
rect 250654 298294 250722 298350
rect 250778 298294 250848 298350
rect 250528 298226 250848 298294
rect 250528 298170 250598 298226
rect 250654 298170 250722 298226
rect 250778 298170 250848 298226
rect 250528 298102 250848 298170
rect 250528 298046 250598 298102
rect 250654 298046 250722 298102
rect 250778 298046 250848 298102
rect 250528 297978 250848 298046
rect 250528 297922 250598 297978
rect 250654 297922 250722 297978
rect 250778 297922 250848 297978
rect 250528 297888 250848 297922
rect 281248 298350 281568 298384
rect 281248 298294 281318 298350
rect 281374 298294 281442 298350
rect 281498 298294 281568 298350
rect 281248 298226 281568 298294
rect 281248 298170 281318 298226
rect 281374 298170 281442 298226
rect 281498 298170 281568 298226
rect 281248 298102 281568 298170
rect 281248 298046 281318 298102
rect 281374 298046 281442 298102
rect 281498 298046 281568 298102
rect 281248 297978 281568 298046
rect 281248 297922 281318 297978
rect 281374 297922 281442 297978
rect 281498 297922 281568 297978
rect 281248 297888 281568 297922
rect 311968 298350 312288 298384
rect 311968 298294 312038 298350
rect 312094 298294 312162 298350
rect 312218 298294 312288 298350
rect 311968 298226 312288 298294
rect 311968 298170 312038 298226
rect 312094 298170 312162 298226
rect 312218 298170 312288 298226
rect 311968 298102 312288 298170
rect 311968 298046 312038 298102
rect 312094 298046 312162 298102
rect 312218 298046 312288 298102
rect 311968 297978 312288 298046
rect 311968 297922 312038 297978
rect 312094 297922 312162 297978
rect 312218 297922 312288 297978
rect 311968 297888 312288 297922
rect 342688 298350 343008 298384
rect 342688 298294 342758 298350
rect 342814 298294 342882 298350
rect 342938 298294 343008 298350
rect 342688 298226 343008 298294
rect 342688 298170 342758 298226
rect 342814 298170 342882 298226
rect 342938 298170 343008 298226
rect 342688 298102 343008 298170
rect 342688 298046 342758 298102
rect 342814 298046 342882 298102
rect 342938 298046 343008 298102
rect 342688 297978 343008 298046
rect 342688 297922 342758 297978
rect 342814 297922 342882 297978
rect 342938 297922 343008 297978
rect 342688 297888 343008 297922
rect 373408 298350 373728 298384
rect 373408 298294 373478 298350
rect 373534 298294 373602 298350
rect 373658 298294 373728 298350
rect 373408 298226 373728 298294
rect 373408 298170 373478 298226
rect 373534 298170 373602 298226
rect 373658 298170 373728 298226
rect 373408 298102 373728 298170
rect 373408 298046 373478 298102
rect 373534 298046 373602 298102
rect 373658 298046 373728 298102
rect 373408 297978 373728 298046
rect 373408 297922 373478 297978
rect 373534 297922 373602 297978
rect 373658 297922 373728 297978
rect 373408 297888 373728 297922
rect 404128 298350 404448 298384
rect 404128 298294 404198 298350
rect 404254 298294 404322 298350
rect 404378 298294 404448 298350
rect 404128 298226 404448 298294
rect 404128 298170 404198 298226
rect 404254 298170 404322 298226
rect 404378 298170 404448 298226
rect 404128 298102 404448 298170
rect 404128 298046 404198 298102
rect 404254 298046 404322 298102
rect 404378 298046 404448 298102
rect 404128 297978 404448 298046
rect 404128 297922 404198 297978
rect 404254 297922 404322 297978
rect 404378 297922 404448 297978
rect 404128 297888 404448 297922
rect 434848 298350 435168 298384
rect 434848 298294 434918 298350
rect 434974 298294 435042 298350
rect 435098 298294 435168 298350
rect 434848 298226 435168 298294
rect 434848 298170 434918 298226
rect 434974 298170 435042 298226
rect 435098 298170 435168 298226
rect 434848 298102 435168 298170
rect 434848 298046 434918 298102
rect 434974 298046 435042 298102
rect 435098 298046 435168 298102
rect 434848 297978 435168 298046
rect 434848 297922 434918 297978
rect 434974 297922 435042 297978
rect 435098 297922 435168 297978
rect 434848 297888 435168 297922
rect 465568 298350 465888 298384
rect 465568 298294 465638 298350
rect 465694 298294 465762 298350
rect 465818 298294 465888 298350
rect 465568 298226 465888 298294
rect 465568 298170 465638 298226
rect 465694 298170 465762 298226
rect 465818 298170 465888 298226
rect 465568 298102 465888 298170
rect 465568 298046 465638 298102
rect 465694 298046 465762 298102
rect 465818 298046 465888 298102
rect 465568 297978 465888 298046
rect 465568 297922 465638 297978
rect 465694 297922 465762 297978
rect 465818 297922 465888 297978
rect 465568 297888 465888 297922
rect 496288 298350 496608 298384
rect 496288 298294 496358 298350
rect 496414 298294 496482 298350
rect 496538 298294 496608 298350
rect 496288 298226 496608 298294
rect 496288 298170 496358 298226
rect 496414 298170 496482 298226
rect 496538 298170 496608 298226
rect 496288 298102 496608 298170
rect 496288 298046 496358 298102
rect 496414 298046 496482 298102
rect 496538 298046 496608 298102
rect 496288 297978 496608 298046
rect 496288 297922 496358 297978
rect 496414 297922 496482 297978
rect 496538 297922 496608 297978
rect 496288 297888 496608 297922
rect 201154 292294 201250 292350
rect 201306 292294 201374 292350
rect 201430 292294 201498 292350
rect 201554 292294 201622 292350
rect 201678 292294 201774 292350
rect 201154 292226 201774 292294
rect 201154 292170 201250 292226
rect 201306 292170 201374 292226
rect 201430 292170 201498 292226
rect 201554 292170 201622 292226
rect 201678 292170 201774 292226
rect 201154 292102 201774 292170
rect 201154 292046 201250 292102
rect 201306 292046 201374 292102
rect 201430 292046 201498 292102
rect 201554 292046 201622 292102
rect 201678 292046 201774 292102
rect 201154 291978 201774 292046
rect 201154 291922 201250 291978
rect 201306 291922 201374 291978
rect 201430 291922 201498 291978
rect 201554 291922 201622 291978
rect 201678 291922 201774 291978
rect 201154 274350 201774 291922
rect 204448 292350 204768 292384
rect 204448 292294 204518 292350
rect 204574 292294 204642 292350
rect 204698 292294 204768 292350
rect 204448 292226 204768 292294
rect 204448 292170 204518 292226
rect 204574 292170 204642 292226
rect 204698 292170 204768 292226
rect 204448 292102 204768 292170
rect 204448 292046 204518 292102
rect 204574 292046 204642 292102
rect 204698 292046 204768 292102
rect 204448 291978 204768 292046
rect 204448 291922 204518 291978
rect 204574 291922 204642 291978
rect 204698 291922 204768 291978
rect 204448 291888 204768 291922
rect 235168 292350 235488 292384
rect 235168 292294 235238 292350
rect 235294 292294 235362 292350
rect 235418 292294 235488 292350
rect 235168 292226 235488 292294
rect 235168 292170 235238 292226
rect 235294 292170 235362 292226
rect 235418 292170 235488 292226
rect 235168 292102 235488 292170
rect 235168 292046 235238 292102
rect 235294 292046 235362 292102
rect 235418 292046 235488 292102
rect 235168 291978 235488 292046
rect 235168 291922 235238 291978
rect 235294 291922 235362 291978
rect 235418 291922 235488 291978
rect 235168 291888 235488 291922
rect 265888 292350 266208 292384
rect 265888 292294 265958 292350
rect 266014 292294 266082 292350
rect 266138 292294 266208 292350
rect 265888 292226 266208 292294
rect 265888 292170 265958 292226
rect 266014 292170 266082 292226
rect 266138 292170 266208 292226
rect 265888 292102 266208 292170
rect 265888 292046 265958 292102
rect 266014 292046 266082 292102
rect 266138 292046 266208 292102
rect 265888 291978 266208 292046
rect 265888 291922 265958 291978
rect 266014 291922 266082 291978
rect 266138 291922 266208 291978
rect 265888 291888 266208 291922
rect 296608 292350 296928 292384
rect 296608 292294 296678 292350
rect 296734 292294 296802 292350
rect 296858 292294 296928 292350
rect 296608 292226 296928 292294
rect 296608 292170 296678 292226
rect 296734 292170 296802 292226
rect 296858 292170 296928 292226
rect 296608 292102 296928 292170
rect 296608 292046 296678 292102
rect 296734 292046 296802 292102
rect 296858 292046 296928 292102
rect 296608 291978 296928 292046
rect 296608 291922 296678 291978
rect 296734 291922 296802 291978
rect 296858 291922 296928 291978
rect 296608 291888 296928 291922
rect 327328 292350 327648 292384
rect 327328 292294 327398 292350
rect 327454 292294 327522 292350
rect 327578 292294 327648 292350
rect 327328 292226 327648 292294
rect 327328 292170 327398 292226
rect 327454 292170 327522 292226
rect 327578 292170 327648 292226
rect 327328 292102 327648 292170
rect 327328 292046 327398 292102
rect 327454 292046 327522 292102
rect 327578 292046 327648 292102
rect 327328 291978 327648 292046
rect 327328 291922 327398 291978
rect 327454 291922 327522 291978
rect 327578 291922 327648 291978
rect 327328 291888 327648 291922
rect 358048 292350 358368 292384
rect 358048 292294 358118 292350
rect 358174 292294 358242 292350
rect 358298 292294 358368 292350
rect 358048 292226 358368 292294
rect 358048 292170 358118 292226
rect 358174 292170 358242 292226
rect 358298 292170 358368 292226
rect 358048 292102 358368 292170
rect 358048 292046 358118 292102
rect 358174 292046 358242 292102
rect 358298 292046 358368 292102
rect 358048 291978 358368 292046
rect 358048 291922 358118 291978
rect 358174 291922 358242 291978
rect 358298 291922 358368 291978
rect 358048 291888 358368 291922
rect 388768 292350 389088 292384
rect 388768 292294 388838 292350
rect 388894 292294 388962 292350
rect 389018 292294 389088 292350
rect 388768 292226 389088 292294
rect 388768 292170 388838 292226
rect 388894 292170 388962 292226
rect 389018 292170 389088 292226
rect 388768 292102 389088 292170
rect 388768 292046 388838 292102
rect 388894 292046 388962 292102
rect 389018 292046 389088 292102
rect 388768 291978 389088 292046
rect 388768 291922 388838 291978
rect 388894 291922 388962 291978
rect 389018 291922 389088 291978
rect 388768 291888 389088 291922
rect 419488 292350 419808 292384
rect 419488 292294 419558 292350
rect 419614 292294 419682 292350
rect 419738 292294 419808 292350
rect 419488 292226 419808 292294
rect 419488 292170 419558 292226
rect 419614 292170 419682 292226
rect 419738 292170 419808 292226
rect 419488 292102 419808 292170
rect 419488 292046 419558 292102
rect 419614 292046 419682 292102
rect 419738 292046 419808 292102
rect 419488 291978 419808 292046
rect 419488 291922 419558 291978
rect 419614 291922 419682 291978
rect 419738 291922 419808 291978
rect 419488 291888 419808 291922
rect 450208 292350 450528 292384
rect 450208 292294 450278 292350
rect 450334 292294 450402 292350
rect 450458 292294 450528 292350
rect 450208 292226 450528 292294
rect 450208 292170 450278 292226
rect 450334 292170 450402 292226
rect 450458 292170 450528 292226
rect 450208 292102 450528 292170
rect 450208 292046 450278 292102
rect 450334 292046 450402 292102
rect 450458 292046 450528 292102
rect 450208 291978 450528 292046
rect 450208 291922 450278 291978
rect 450334 291922 450402 291978
rect 450458 291922 450528 291978
rect 450208 291888 450528 291922
rect 480928 292350 481248 292384
rect 480928 292294 480998 292350
rect 481054 292294 481122 292350
rect 481178 292294 481248 292350
rect 480928 292226 481248 292294
rect 480928 292170 480998 292226
rect 481054 292170 481122 292226
rect 481178 292170 481248 292226
rect 480928 292102 481248 292170
rect 480928 292046 480998 292102
rect 481054 292046 481122 292102
rect 481178 292046 481248 292102
rect 480928 291978 481248 292046
rect 480928 291922 480998 291978
rect 481054 291922 481122 291978
rect 481178 291922 481248 291978
rect 480928 291888 481248 291922
rect 507154 292350 507774 309922
rect 507154 292294 507250 292350
rect 507306 292294 507374 292350
rect 507430 292294 507498 292350
rect 507554 292294 507622 292350
rect 507678 292294 507774 292350
rect 507154 292226 507774 292294
rect 507154 292170 507250 292226
rect 507306 292170 507374 292226
rect 507430 292170 507498 292226
rect 507554 292170 507622 292226
rect 507678 292170 507774 292226
rect 507154 292102 507774 292170
rect 507154 292046 507250 292102
rect 507306 292046 507374 292102
rect 507430 292046 507498 292102
rect 507554 292046 507622 292102
rect 507678 292046 507774 292102
rect 507154 291978 507774 292046
rect 507154 291922 507250 291978
rect 507306 291922 507374 291978
rect 507430 291922 507498 291978
rect 507554 291922 507622 291978
rect 507678 291922 507774 291978
rect 219808 280350 220128 280384
rect 219808 280294 219878 280350
rect 219934 280294 220002 280350
rect 220058 280294 220128 280350
rect 219808 280226 220128 280294
rect 219808 280170 219878 280226
rect 219934 280170 220002 280226
rect 220058 280170 220128 280226
rect 219808 280102 220128 280170
rect 219808 280046 219878 280102
rect 219934 280046 220002 280102
rect 220058 280046 220128 280102
rect 219808 279978 220128 280046
rect 219808 279922 219878 279978
rect 219934 279922 220002 279978
rect 220058 279922 220128 279978
rect 219808 279888 220128 279922
rect 250528 280350 250848 280384
rect 250528 280294 250598 280350
rect 250654 280294 250722 280350
rect 250778 280294 250848 280350
rect 250528 280226 250848 280294
rect 250528 280170 250598 280226
rect 250654 280170 250722 280226
rect 250778 280170 250848 280226
rect 250528 280102 250848 280170
rect 250528 280046 250598 280102
rect 250654 280046 250722 280102
rect 250778 280046 250848 280102
rect 250528 279978 250848 280046
rect 250528 279922 250598 279978
rect 250654 279922 250722 279978
rect 250778 279922 250848 279978
rect 250528 279888 250848 279922
rect 281248 280350 281568 280384
rect 281248 280294 281318 280350
rect 281374 280294 281442 280350
rect 281498 280294 281568 280350
rect 281248 280226 281568 280294
rect 281248 280170 281318 280226
rect 281374 280170 281442 280226
rect 281498 280170 281568 280226
rect 281248 280102 281568 280170
rect 281248 280046 281318 280102
rect 281374 280046 281442 280102
rect 281498 280046 281568 280102
rect 281248 279978 281568 280046
rect 281248 279922 281318 279978
rect 281374 279922 281442 279978
rect 281498 279922 281568 279978
rect 281248 279888 281568 279922
rect 311968 280350 312288 280384
rect 311968 280294 312038 280350
rect 312094 280294 312162 280350
rect 312218 280294 312288 280350
rect 311968 280226 312288 280294
rect 311968 280170 312038 280226
rect 312094 280170 312162 280226
rect 312218 280170 312288 280226
rect 311968 280102 312288 280170
rect 311968 280046 312038 280102
rect 312094 280046 312162 280102
rect 312218 280046 312288 280102
rect 311968 279978 312288 280046
rect 311968 279922 312038 279978
rect 312094 279922 312162 279978
rect 312218 279922 312288 279978
rect 311968 279888 312288 279922
rect 342688 280350 343008 280384
rect 342688 280294 342758 280350
rect 342814 280294 342882 280350
rect 342938 280294 343008 280350
rect 342688 280226 343008 280294
rect 342688 280170 342758 280226
rect 342814 280170 342882 280226
rect 342938 280170 343008 280226
rect 342688 280102 343008 280170
rect 342688 280046 342758 280102
rect 342814 280046 342882 280102
rect 342938 280046 343008 280102
rect 342688 279978 343008 280046
rect 342688 279922 342758 279978
rect 342814 279922 342882 279978
rect 342938 279922 343008 279978
rect 342688 279888 343008 279922
rect 373408 280350 373728 280384
rect 373408 280294 373478 280350
rect 373534 280294 373602 280350
rect 373658 280294 373728 280350
rect 373408 280226 373728 280294
rect 373408 280170 373478 280226
rect 373534 280170 373602 280226
rect 373658 280170 373728 280226
rect 373408 280102 373728 280170
rect 373408 280046 373478 280102
rect 373534 280046 373602 280102
rect 373658 280046 373728 280102
rect 373408 279978 373728 280046
rect 373408 279922 373478 279978
rect 373534 279922 373602 279978
rect 373658 279922 373728 279978
rect 373408 279888 373728 279922
rect 404128 280350 404448 280384
rect 404128 280294 404198 280350
rect 404254 280294 404322 280350
rect 404378 280294 404448 280350
rect 404128 280226 404448 280294
rect 404128 280170 404198 280226
rect 404254 280170 404322 280226
rect 404378 280170 404448 280226
rect 404128 280102 404448 280170
rect 404128 280046 404198 280102
rect 404254 280046 404322 280102
rect 404378 280046 404448 280102
rect 404128 279978 404448 280046
rect 404128 279922 404198 279978
rect 404254 279922 404322 279978
rect 404378 279922 404448 279978
rect 404128 279888 404448 279922
rect 434848 280350 435168 280384
rect 434848 280294 434918 280350
rect 434974 280294 435042 280350
rect 435098 280294 435168 280350
rect 434848 280226 435168 280294
rect 434848 280170 434918 280226
rect 434974 280170 435042 280226
rect 435098 280170 435168 280226
rect 434848 280102 435168 280170
rect 434848 280046 434918 280102
rect 434974 280046 435042 280102
rect 435098 280046 435168 280102
rect 434848 279978 435168 280046
rect 434848 279922 434918 279978
rect 434974 279922 435042 279978
rect 435098 279922 435168 279978
rect 434848 279888 435168 279922
rect 465568 280350 465888 280384
rect 465568 280294 465638 280350
rect 465694 280294 465762 280350
rect 465818 280294 465888 280350
rect 465568 280226 465888 280294
rect 465568 280170 465638 280226
rect 465694 280170 465762 280226
rect 465818 280170 465888 280226
rect 465568 280102 465888 280170
rect 465568 280046 465638 280102
rect 465694 280046 465762 280102
rect 465818 280046 465888 280102
rect 465568 279978 465888 280046
rect 465568 279922 465638 279978
rect 465694 279922 465762 279978
rect 465818 279922 465888 279978
rect 465568 279888 465888 279922
rect 496288 280350 496608 280384
rect 496288 280294 496358 280350
rect 496414 280294 496482 280350
rect 496538 280294 496608 280350
rect 496288 280226 496608 280294
rect 496288 280170 496358 280226
rect 496414 280170 496482 280226
rect 496538 280170 496608 280226
rect 496288 280102 496608 280170
rect 496288 280046 496358 280102
rect 496414 280046 496482 280102
rect 496538 280046 496608 280102
rect 496288 279978 496608 280046
rect 496288 279922 496358 279978
rect 496414 279922 496482 279978
rect 496538 279922 496608 279978
rect 496288 279888 496608 279922
rect 201154 274294 201250 274350
rect 201306 274294 201374 274350
rect 201430 274294 201498 274350
rect 201554 274294 201622 274350
rect 201678 274294 201774 274350
rect 201154 274226 201774 274294
rect 201154 274170 201250 274226
rect 201306 274170 201374 274226
rect 201430 274170 201498 274226
rect 201554 274170 201622 274226
rect 201678 274170 201774 274226
rect 201154 274102 201774 274170
rect 201154 274046 201250 274102
rect 201306 274046 201374 274102
rect 201430 274046 201498 274102
rect 201554 274046 201622 274102
rect 201678 274046 201774 274102
rect 201154 273978 201774 274046
rect 201154 273922 201250 273978
rect 201306 273922 201374 273978
rect 201430 273922 201498 273978
rect 201554 273922 201622 273978
rect 201678 273922 201774 273978
rect 201154 256350 201774 273922
rect 204448 274350 204768 274384
rect 204448 274294 204518 274350
rect 204574 274294 204642 274350
rect 204698 274294 204768 274350
rect 204448 274226 204768 274294
rect 204448 274170 204518 274226
rect 204574 274170 204642 274226
rect 204698 274170 204768 274226
rect 204448 274102 204768 274170
rect 204448 274046 204518 274102
rect 204574 274046 204642 274102
rect 204698 274046 204768 274102
rect 204448 273978 204768 274046
rect 204448 273922 204518 273978
rect 204574 273922 204642 273978
rect 204698 273922 204768 273978
rect 204448 273888 204768 273922
rect 235168 274350 235488 274384
rect 235168 274294 235238 274350
rect 235294 274294 235362 274350
rect 235418 274294 235488 274350
rect 235168 274226 235488 274294
rect 235168 274170 235238 274226
rect 235294 274170 235362 274226
rect 235418 274170 235488 274226
rect 235168 274102 235488 274170
rect 235168 274046 235238 274102
rect 235294 274046 235362 274102
rect 235418 274046 235488 274102
rect 235168 273978 235488 274046
rect 235168 273922 235238 273978
rect 235294 273922 235362 273978
rect 235418 273922 235488 273978
rect 235168 273888 235488 273922
rect 265888 274350 266208 274384
rect 265888 274294 265958 274350
rect 266014 274294 266082 274350
rect 266138 274294 266208 274350
rect 265888 274226 266208 274294
rect 265888 274170 265958 274226
rect 266014 274170 266082 274226
rect 266138 274170 266208 274226
rect 265888 274102 266208 274170
rect 265888 274046 265958 274102
rect 266014 274046 266082 274102
rect 266138 274046 266208 274102
rect 265888 273978 266208 274046
rect 265888 273922 265958 273978
rect 266014 273922 266082 273978
rect 266138 273922 266208 273978
rect 265888 273888 266208 273922
rect 296608 274350 296928 274384
rect 296608 274294 296678 274350
rect 296734 274294 296802 274350
rect 296858 274294 296928 274350
rect 296608 274226 296928 274294
rect 296608 274170 296678 274226
rect 296734 274170 296802 274226
rect 296858 274170 296928 274226
rect 296608 274102 296928 274170
rect 296608 274046 296678 274102
rect 296734 274046 296802 274102
rect 296858 274046 296928 274102
rect 296608 273978 296928 274046
rect 296608 273922 296678 273978
rect 296734 273922 296802 273978
rect 296858 273922 296928 273978
rect 296608 273888 296928 273922
rect 327328 274350 327648 274384
rect 327328 274294 327398 274350
rect 327454 274294 327522 274350
rect 327578 274294 327648 274350
rect 327328 274226 327648 274294
rect 327328 274170 327398 274226
rect 327454 274170 327522 274226
rect 327578 274170 327648 274226
rect 327328 274102 327648 274170
rect 327328 274046 327398 274102
rect 327454 274046 327522 274102
rect 327578 274046 327648 274102
rect 327328 273978 327648 274046
rect 327328 273922 327398 273978
rect 327454 273922 327522 273978
rect 327578 273922 327648 273978
rect 327328 273888 327648 273922
rect 358048 274350 358368 274384
rect 358048 274294 358118 274350
rect 358174 274294 358242 274350
rect 358298 274294 358368 274350
rect 358048 274226 358368 274294
rect 358048 274170 358118 274226
rect 358174 274170 358242 274226
rect 358298 274170 358368 274226
rect 358048 274102 358368 274170
rect 358048 274046 358118 274102
rect 358174 274046 358242 274102
rect 358298 274046 358368 274102
rect 358048 273978 358368 274046
rect 358048 273922 358118 273978
rect 358174 273922 358242 273978
rect 358298 273922 358368 273978
rect 358048 273888 358368 273922
rect 388768 274350 389088 274384
rect 388768 274294 388838 274350
rect 388894 274294 388962 274350
rect 389018 274294 389088 274350
rect 388768 274226 389088 274294
rect 388768 274170 388838 274226
rect 388894 274170 388962 274226
rect 389018 274170 389088 274226
rect 388768 274102 389088 274170
rect 388768 274046 388838 274102
rect 388894 274046 388962 274102
rect 389018 274046 389088 274102
rect 388768 273978 389088 274046
rect 388768 273922 388838 273978
rect 388894 273922 388962 273978
rect 389018 273922 389088 273978
rect 388768 273888 389088 273922
rect 419488 274350 419808 274384
rect 419488 274294 419558 274350
rect 419614 274294 419682 274350
rect 419738 274294 419808 274350
rect 419488 274226 419808 274294
rect 419488 274170 419558 274226
rect 419614 274170 419682 274226
rect 419738 274170 419808 274226
rect 419488 274102 419808 274170
rect 419488 274046 419558 274102
rect 419614 274046 419682 274102
rect 419738 274046 419808 274102
rect 419488 273978 419808 274046
rect 419488 273922 419558 273978
rect 419614 273922 419682 273978
rect 419738 273922 419808 273978
rect 419488 273888 419808 273922
rect 450208 274350 450528 274384
rect 450208 274294 450278 274350
rect 450334 274294 450402 274350
rect 450458 274294 450528 274350
rect 450208 274226 450528 274294
rect 450208 274170 450278 274226
rect 450334 274170 450402 274226
rect 450458 274170 450528 274226
rect 450208 274102 450528 274170
rect 450208 274046 450278 274102
rect 450334 274046 450402 274102
rect 450458 274046 450528 274102
rect 450208 273978 450528 274046
rect 450208 273922 450278 273978
rect 450334 273922 450402 273978
rect 450458 273922 450528 273978
rect 450208 273888 450528 273922
rect 480928 274350 481248 274384
rect 480928 274294 480998 274350
rect 481054 274294 481122 274350
rect 481178 274294 481248 274350
rect 480928 274226 481248 274294
rect 480928 274170 480998 274226
rect 481054 274170 481122 274226
rect 481178 274170 481248 274226
rect 480928 274102 481248 274170
rect 480928 274046 480998 274102
rect 481054 274046 481122 274102
rect 481178 274046 481248 274102
rect 480928 273978 481248 274046
rect 480928 273922 480998 273978
rect 481054 273922 481122 273978
rect 481178 273922 481248 273978
rect 480928 273888 481248 273922
rect 507154 274350 507774 291922
rect 507154 274294 507250 274350
rect 507306 274294 507374 274350
rect 507430 274294 507498 274350
rect 507554 274294 507622 274350
rect 507678 274294 507774 274350
rect 507154 274226 507774 274294
rect 507154 274170 507250 274226
rect 507306 274170 507374 274226
rect 507430 274170 507498 274226
rect 507554 274170 507622 274226
rect 507678 274170 507774 274226
rect 507154 274102 507774 274170
rect 507154 274046 507250 274102
rect 507306 274046 507374 274102
rect 507430 274046 507498 274102
rect 507554 274046 507622 274102
rect 507678 274046 507774 274102
rect 507154 273978 507774 274046
rect 507154 273922 507250 273978
rect 507306 273922 507374 273978
rect 507430 273922 507498 273978
rect 507554 273922 507622 273978
rect 507678 273922 507774 273978
rect 219808 262350 220128 262384
rect 219808 262294 219878 262350
rect 219934 262294 220002 262350
rect 220058 262294 220128 262350
rect 219808 262226 220128 262294
rect 219808 262170 219878 262226
rect 219934 262170 220002 262226
rect 220058 262170 220128 262226
rect 219808 262102 220128 262170
rect 219808 262046 219878 262102
rect 219934 262046 220002 262102
rect 220058 262046 220128 262102
rect 219808 261978 220128 262046
rect 219808 261922 219878 261978
rect 219934 261922 220002 261978
rect 220058 261922 220128 261978
rect 219808 261888 220128 261922
rect 250528 262350 250848 262384
rect 250528 262294 250598 262350
rect 250654 262294 250722 262350
rect 250778 262294 250848 262350
rect 250528 262226 250848 262294
rect 250528 262170 250598 262226
rect 250654 262170 250722 262226
rect 250778 262170 250848 262226
rect 250528 262102 250848 262170
rect 250528 262046 250598 262102
rect 250654 262046 250722 262102
rect 250778 262046 250848 262102
rect 250528 261978 250848 262046
rect 250528 261922 250598 261978
rect 250654 261922 250722 261978
rect 250778 261922 250848 261978
rect 250528 261888 250848 261922
rect 281248 262350 281568 262384
rect 281248 262294 281318 262350
rect 281374 262294 281442 262350
rect 281498 262294 281568 262350
rect 281248 262226 281568 262294
rect 281248 262170 281318 262226
rect 281374 262170 281442 262226
rect 281498 262170 281568 262226
rect 281248 262102 281568 262170
rect 281248 262046 281318 262102
rect 281374 262046 281442 262102
rect 281498 262046 281568 262102
rect 281248 261978 281568 262046
rect 281248 261922 281318 261978
rect 281374 261922 281442 261978
rect 281498 261922 281568 261978
rect 281248 261888 281568 261922
rect 311968 262350 312288 262384
rect 311968 262294 312038 262350
rect 312094 262294 312162 262350
rect 312218 262294 312288 262350
rect 311968 262226 312288 262294
rect 311968 262170 312038 262226
rect 312094 262170 312162 262226
rect 312218 262170 312288 262226
rect 311968 262102 312288 262170
rect 311968 262046 312038 262102
rect 312094 262046 312162 262102
rect 312218 262046 312288 262102
rect 311968 261978 312288 262046
rect 311968 261922 312038 261978
rect 312094 261922 312162 261978
rect 312218 261922 312288 261978
rect 311968 261888 312288 261922
rect 342688 262350 343008 262384
rect 342688 262294 342758 262350
rect 342814 262294 342882 262350
rect 342938 262294 343008 262350
rect 342688 262226 343008 262294
rect 342688 262170 342758 262226
rect 342814 262170 342882 262226
rect 342938 262170 343008 262226
rect 342688 262102 343008 262170
rect 342688 262046 342758 262102
rect 342814 262046 342882 262102
rect 342938 262046 343008 262102
rect 342688 261978 343008 262046
rect 342688 261922 342758 261978
rect 342814 261922 342882 261978
rect 342938 261922 343008 261978
rect 342688 261888 343008 261922
rect 373408 262350 373728 262384
rect 373408 262294 373478 262350
rect 373534 262294 373602 262350
rect 373658 262294 373728 262350
rect 373408 262226 373728 262294
rect 373408 262170 373478 262226
rect 373534 262170 373602 262226
rect 373658 262170 373728 262226
rect 373408 262102 373728 262170
rect 373408 262046 373478 262102
rect 373534 262046 373602 262102
rect 373658 262046 373728 262102
rect 373408 261978 373728 262046
rect 373408 261922 373478 261978
rect 373534 261922 373602 261978
rect 373658 261922 373728 261978
rect 373408 261888 373728 261922
rect 404128 262350 404448 262384
rect 404128 262294 404198 262350
rect 404254 262294 404322 262350
rect 404378 262294 404448 262350
rect 404128 262226 404448 262294
rect 404128 262170 404198 262226
rect 404254 262170 404322 262226
rect 404378 262170 404448 262226
rect 404128 262102 404448 262170
rect 404128 262046 404198 262102
rect 404254 262046 404322 262102
rect 404378 262046 404448 262102
rect 404128 261978 404448 262046
rect 404128 261922 404198 261978
rect 404254 261922 404322 261978
rect 404378 261922 404448 261978
rect 404128 261888 404448 261922
rect 434848 262350 435168 262384
rect 434848 262294 434918 262350
rect 434974 262294 435042 262350
rect 435098 262294 435168 262350
rect 434848 262226 435168 262294
rect 434848 262170 434918 262226
rect 434974 262170 435042 262226
rect 435098 262170 435168 262226
rect 434848 262102 435168 262170
rect 434848 262046 434918 262102
rect 434974 262046 435042 262102
rect 435098 262046 435168 262102
rect 434848 261978 435168 262046
rect 434848 261922 434918 261978
rect 434974 261922 435042 261978
rect 435098 261922 435168 261978
rect 434848 261888 435168 261922
rect 465568 262350 465888 262384
rect 465568 262294 465638 262350
rect 465694 262294 465762 262350
rect 465818 262294 465888 262350
rect 465568 262226 465888 262294
rect 465568 262170 465638 262226
rect 465694 262170 465762 262226
rect 465818 262170 465888 262226
rect 465568 262102 465888 262170
rect 465568 262046 465638 262102
rect 465694 262046 465762 262102
rect 465818 262046 465888 262102
rect 465568 261978 465888 262046
rect 465568 261922 465638 261978
rect 465694 261922 465762 261978
rect 465818 261922 465888 261978
rect 465568 261888 465888 261922
rect 496288 262350 496608 262384
rect 496288 262294 496358 262350
rect 496414 262294 496482 262350
rect 496538 262294 496608 262350
rect 496288 262226 496608 262294
rect 496288 262170 496358 262226
rect 496414 262170 496482 262226
rect 496538 262170 496608 262226
rect 496288 262102 496608 262170
rect 496288 262046 496358 262102
rect 496414 262046 496482 262102
rect 496538 262046 496608 262102
rect 496288 261978 496608 262046
rect 496288 261922 496358 261978
rect 496414 261922 496482 261978
rect 496538 261922 496608 261978
rect 496288 261888 496608 261922
rect 201154 256294 201250 256350
rect 201306 256294 201374 256350
rect 201430 256294 201498 256350
rect 201554 256294 201622 256350
rect 201678 256294 201774 256350
rect 201154 256226 201774 256294
rect 201154 256170 201250 256226
rect 201306 256170 201374 256226
rect 201430 256170 201498 256226
rect 201554 256170 201622 256226
rect 201678 256170 201774 256226
rect 201154 256102 201774 256170
rect 201154 256046 201250 256102
rect 201306 256046 201374 256102
rect 201430 256046 201498 256102
rect 201554 256046 201622 256102
rect 201678 256046 201774 256102
rect 201154 255978 201774 256046
rect 201154 255922 201250 255978
rect 201306 255922 201374 255978
rect 201430 255922 201498 255978
rect 201554 255922 201622 255978
rect 201678 255922 201774 255978
rect 201154 238350 201774 255922
rect 204448 256350 204768 256384
rect 204448 256294 204518 256350
rect 204574 256294 204642 256350
rect 204698 256294 204768 256350
rect 204448 256226 204768 256294
rect 204448 256170 204518 256226
rect 204574 256170 204642 256226
rect 204698 256170 204768 256226
rect 204448 256102 204768 256170
rect 204448 256046 204518 256102
rect 204574 256046 204642 256102
rect 204698 256046 204768 256102
rect 204448 255978 204768 256046
rect 204448 255922 204518 255978
rect 204574 255922 204642 255978
rect 204698 255922 204768 255978
rect 204448 255888 204768 255922
rect 235168 256350 235488 256384
rect 235168 256294 235238 256350
rect 235294 256294 235362 256350
rect 235418 256294 235488 256350
rect 235168 256226 235488 256294
rect 235168 256170 235238 256226
rect 235294 256170 235362 256226
rect 235418 256170 235488 256226
rect 235168 256102 235488 256170
rect 235168 256046 235238 256102
rect 235294 256046 235362 256102
rect 235418 256046 235488 256102
rect 235168 255978 235488 256046
rect 235168 255922 235238 255978
rect 235294 255922 235362 255978
rect 235418 255922 235488 255978
rect 235168 255888 235488 255922
rect 265888 256350 266208 256384
rect 265888 256294 265958 256350
rect 266014 256294 266082 256350
rect 266138 256294 266208 256350
rect 265888 256226 266208 256294
rect 265888 256170 265958 256226
rect 266014 256170 266082 256226
rect 266138 256170 266208 256226
rect 265888 256102 266208 256170
rect 265888 256046 265958 256102
rect 266014 256046 266082 256102
rect 266138 256046 266208 256102
rect 265888 255978 266208 256046
rect 265888 255922 265958 255978
rect 266014 255922 266082 255978
rect 266138 255922 266208 255978
rect 265888 255888 266208 255922
rect 296608 256350 296928 256384
rect 296608 256294 296678 256350
rect 296734 256294 296802 256350
rect 296858 256294 296928 256350
rect 296608 256226 296928 256294
rect 296608 256170 296678 256226
rect 296734 256170 296802 256226
rect 296858 256170 296928 256226
rect 296608 256102 296928 256170
rect 296608 256046 296678 256102
rect 296734 256046 296802 256102
rect 296858 256046 296928 256102
rect 296608 255978 296928 256046
rect 296608 255922 296678 255978
rect 296734 255922 296802 255978
rect 296858 255922 296928 255978
rect 296608 255888 296928 255922
rect 327328 256350 327648 256384
rect 327328 256294 327398 256350
rect 327454 256294 327522 256350
rect 327578 256294 327648 256350
rect 327328 256226 327648 256294
rect 327328 256170 327398 256226
rect 327454 256170 327522 256226
rect 327578 256170 327648 256226
rect 327328 256102 327648 256170
rect 327328 256046 327398 256102
rect 327454 256046 327522 256102
rect 327578 256046 327648 256102
rect 327328 255978 327648 256046
rect 327328 255922 327398 255978
rect 327454 255922 327522 255978
rect 327578 255922 327648 255978
rect 327328 255888 327648 255922
rect 358048 256350 358368 256384
rect 358048 256294 358118 256350
rect 358174 256294 358242 256350
rect 358298 256294 358368 256350
rect 358048 256226 358368 256294
rect 358048 256170 358118 256226
rect 358174 256170 358242 256226
rect 358298 256170 358368 256226
rect 358048 256102 358368 256170
rect 358048 256046 358118 256102
rect 358174 256046 358242 256102
rect 358298 256046 358368 256102
rect 358048 255978 358368 256046
rect 358048 255922 358118 255978
rect 358174 255922 358242 255978
rect 358298 255922 358368 255978
rect 358048 255888 358368 255922
rect 388768 256350 389088 256384
rect 388768 256294 388838 256350
rect 388894 256294 388962 256350
rect 389018 256294 389088 256350
rect 388768 256226 389088 256294
rect 388768 256170 388838 256226
rect 388894 256170 388962 256226
rect 389018 256170 389088 256226
rect 388768 256102 389088 256170
rect 388768 256046 388838 256102
rect 388894 256046 388962 256102
rect 389018 256046 389088 256102
rect 388768 255978 389088 256046
rect 388768 255922 388838 255978
rect 388894 255922 388962 255978
rect 389018 255922 389088 255978
rect 388768 255888 389088 255922
rect 419488 256350 419808 256384
rect 419488 256294 419558 256350
rect 419614 256294 419682 256350
rect 419738 256294 419808 256350
rect 419488 256226 419808 256294
rect 419488 256170 419558 256226
rect 419614 256170 419682 256226
rect 419738 256170 419808 256226
rect 419488 256102 419808 256170
rect 419488 256046 419558 256102
rect 419614 256046 419682 256102
rect 419738 256046 419808 256102
rect 419488 255978 419808 256046
rect 419488 255922 419558 255978
rect 419614 255922 419682 255978
rect 419738 255922 419808 255978
rect 419488 255888 419808 255922
rect 450208 256350 450528 256384
rect 450208 256294 450278 256350
rect 450334 256294 450402 256350
rect 450458 256294 450528 256350
rect 450208 256226 450528 256294
rect 450208 256170 450278 256226
rect 450334 256170 450402 256226
rect 450458 256170 450528 256226
rect 450208 256102 450528 256170
rect 450208 256046 450278 256102
rect 450334 256046 450402 256102
rect 450458 256046 450528 256102
rect 450208 255978 450528 256046
rect 450208 255922 450278 255978
rect 450334 255922 450402 255978
rect 450458 255922 450528 255978
rect 450208 255888 450528 255922
rect 480928 256350 481248 256384
rect 480928 256294 480998 256350
rect 481054 256294 481122 256350
rect 481178 256294 481248 256350
rect 480928 256226 481248 256294
rect 480928 256170 480998 256226
rect 481054 256170 481122 256226
rect 481178 256170 481248 256226
rect 480928 256102 481248 256170
rect 480928 256046 480998 256102
rect 481054 256046 481122 256102
rect 481178 256046 481248 256102
rect 480928 255978 481248 256046
rect 480928 255922 480998 255978
rect 481054 255922 481122 255978
rect 481178 255922 481248 255978
rect 480928 255888 481248 255922
rect 507154 256350 507774 273922
rect 507154 256294 507250 256350
rect 507306 256294 507374 256350
rect 507430 256294 507498 256350
rect 507554 256294 507622 256350
rect 507678 256294 507774 256350
rect 507154 256226 507774 256294
rect 507154 256170 507250 256226
rect 507306 256170 507374 256226
rect 507430 256170 507498 256226
rect 507554 256170 507622 256226
rect 507678 256170 507774 256226
rect 507154 256102 507774 256170
rect 507154 256046 507250 256102
rect 507306 256046 507374 256102
rect 507430 256046 507498 256102
rect 507554 256046 507622 256102
rect 507678 256046 507774 256102
rect 507154 255978 507774 256046
rect 507154 255922 507250 255978
rect 507306 255922 507374 255978
rect 507430 255922 507498 255978
rect 507554 255922 507622 255978
rect 507678 255922 507774 255978
rect 219808 244350 220128 244384
rect 219808 244294 219878 244350
rect 219934 244294 220002 244350
rect 220058 244294 220128 244350
rect 219808 244226 220128 244294
rect 219808 244170 219878 244226
rect 219934 244170 220002 244226
rect 220058 244170 220128 244226
rect 219808 244102 220128 244170
rect 219808 244046 219878 244102
rect 219934 244046 220002 244102
rect 220058 244046 220128 244102
rect 219808 243978 220128 244046
rect 219808 243922 219878 243978
rect 219934 243922 220002 243978
rect 220058 243922 220128 243978
rect 219808 243888 220128 243922
rect 250528 244350 250848 244384
rect 250528 244294 250598 244350
rect 250654 244294 250722 244350
rect 250778 244294 250848 244350
rect 250528 244226 250848 244294
rect 250528 244170 250598 244226
rect 250654 244170 250722 244226
rect 250778 244170 250848 244226
rect 250528 244102 250848 244170
rect 250528 244046 250598 244102
rect 250654 244046 250722 244102
rect 250778 244046 250848 244102
rect 250528 243978 250848 244046
rect 250528 243922 250598 243978
rect 250654 243922 250722 243978
rect 250778 243922 250848 243978
rect 250528 243888 250848 243922
rect 281248 244350 281568 244384
rect 281248 244294 281318 244350
rect 281374 244294 281442 244350
rect 281498 244294 281568 244350
rect 281248 244226 281568 244294
rect 281248 244170 281318 244226
rect 281374 244170 281442 244226
rect 281498 244170 281568 244226
rect 281248 244102 281568 244170
rect 281248 244046 281318 244102
rect 281374 244046 281442 244102
rect 281498 244046 281568 244102
rect 281248 243978 281568 244046
rect 281248 243922 281318 243978
rect 281374 243922 281442 243978
rect 281498 243922 281568 243978
rect 281248 243888 281568 243922
rect 311968 244350 312288 244384
rect 311968 244294 312038 244350
rect 312094 244294 312162 244350
rect 312218 244294 312288 244350
rect 311968 244226 312288 244294
rect 311968 244170 312038 244226
rect 312094 244170 312162 244226
rect 312218 244170 312288 244226
rect 311968 244102 312288 244170
rect 311968 244046 312038 244102
rect 312094 244046 312162 244102
rect 312218 244046 312288 244102
rect 311968 243978 312288 244046
rect 311968 243922 312038 243978
rect 312094 243922 312162 243978
rect 312218 243922 312288 243978
rect 311968 243888 312288 243922
rect 342688 244350 343008 244384
rect 342688 244294 342758 244350
rect 342814 244294 342882 244350
rect 342938 244294 343008 244350
rect 342688 244226 343008 244294
rect 342688 244170 342758 244226
rect 342814 244170 342882 244226
rect 342938 244170 343008 244226
rect 342688 244102 343008 244170
rect 342688 244046 342758 244102
rect 342814 244046 342882 244102
rect 342938 244046 343008 244102
rect 342688 243978 343008 244046
rect 342688 243922 342758 243978
rect 342814 243922 342882 243978
rect 342938 243922 343008 243978
rect 342688 243888 343008 243922
rect 373408 244350 373728 244384
rect 373408 244294 373478 244350
rect 373534 244294 373602 244350
rect 373658 244294 373728 244350
rect 373408 244226 373728 244294
rect 373408 244170 373478 244226
rect 373534 244170 373602 244226
rect 373658 244170 373728 244226
rect 373408 244102 373728 244170
rect 373408 244046 373478 244102
rect 373534 244046 373602 244102
rect 373658 244046 373728 244102
rect 373408 243978 373728 244046
rect 373408 243922 373478 243978
rect 373534 243922 373602 243978
rect 373658 243922 373728 243978
rect 373408 243888 373728 243922
rect 404128 244350 404448 244384
rect 404128 244294 404198 244350
rect 404254 244294 404322 244350
rect 404378 244294 404448 244350
rect 404128 244226 404448 244294
rect 404128 244170 404198 244226
rect 404254 244170 404322 244226
rect 404378 244170 404448 244226
rect 404128 244102 404448 244170
rect 404128 244046 404198 244102
rect 404254 244046 404322 244102
rect 404378 244046 404448 244102
rect 404128 243978 404448 244046
rect 404128 243922 404198 243978
rect 404254 243922 404322 243978
rect 404378 243922 404448 243978
rect 404128 243888 404448 243922
rect 434848 244350 435168 244384
rect 434848 244294 434918 244350
rect 434974 244294 435042 244350
rect 435098 244294 435168 244350
rect 434848 244226 435168 244294
rect 434848 244170 434918 244226
rect 434974 244170 435042 244226
rect 435098 244170 435168 244226
rect 434848 244102 435168 244170
rect 434848 244046 434918 244102
rect 434974 244046 435042 244102
rect 435098 244046 435168 244102
rect 434848 243978 435168 244046
rect 434848 243922 434918 243978
rect 434974 243922 435042 243978
rect 435098 243922 435168 243978
rect 434848 243888 435168 243922
rect 465568 244350 465888 244384
rect 465568 244294 465638 244350
rect 465694 244294 465762 244350
rect 465818 244294 465888 244350
rect 465568 244226 465888 244294
rect 465568 244170 465638 244226
rect 465694 244170 465762 244226
rect 465818 244170 465888 244226
rect 465568 244102 465888 244170
rect 465568 244046 465638 244102
rect 465694 244046 465762 244102
rect 465818 244046 465888 244102
rect 465568 243978 465888 244046
rect 465568 243922 465638 243978
rect 465694 243922 465762 243978
rect 465818 243922 465888 243978
rect 465568 243888 465888 243922
rect 496288 244350 496608 244384
rect 496288 244294 496358 244350
rect 496414 244294 496482 244350
rect 496538 244294 496608 244350
rect 496288 244226 496608 244294
rect 496288 244170 496358 244226
rect 496414 244170 496482 244226
rect 496538 244170 496608 244226
rect 496288 244102 496608 244170
rect 496288 244046 496358 244102
rect 496414 244046 496482 244102
rect 496538 244046 496608 244102
rect 496288 243978 496608 244046
rect 496288 243922 496358 243978
rect 496414 243922 496482 243978
rect 496538 243922 496608 243978
rect 496288 243888 496608 243922
rect 201154 238294 201250 238350
rect 201306 238294 201374 238350
rect 201430 238294 201498 238350
rect 201554 238294 201622 238350
rect 201678 238294 201774 238350
rect 201154 238226 201774 238294
rect 201154 238170 201250 238226
rect 201306 238170 201374 238226
rect 201430 238170 201498 238226
rect 201554 238170 201622 238226
rect 201678 238170 201774 238226
rect 201154 238102 201774 238170
rect 201154 238046 201250 238102
rect 201306 238046 201374 238102
rect 201430 238046 201498 238102
rect 201554 238046 201622 238102
rect 201678 238046 201774 238102
rect 201154 237978 201774 238046
rect 201154 237922 201250 237978
rect 201306 237922 201374 237978
rect 201430 237922 201498 237978
rect 201554 237922 201622 237978
rect 201678 237922 201774 237978
rect 201154 220350 201774 237922
rect 204448 238350 204768 238384
rect 204448 238294 204518 238350
rect 204574 238294 204642 238350
rect 204698 238294 204768 238350
rect 204448 238226 204768 238294
rect 204448 238170 204518 238226
rect 204574 238170 204642 238226
rect 204698 238170 204768 238226
rect 204448 238102 204768 238170
rect 204448 238046 204518 238102
rect 204574 238046 204642 238102
rect 204698 238046 204768 238102
rect 204448 237978 204768 238046
rect 204448 237922 204518 237978
rect 204574 237922 204642 237978
rect 204698 237922 204768 237978
rect 204448 237888 204768 237922
rect 235168 238350 235488 238384
rect 235168 238294 235238 238350
rect 235294 238294 235362 238350
rect 235418 238294 235488 238350
rect 235168 238226 235488 238294
rect 235168 238170 235238 238226
rect 235294 238170 235362 238226
rect 235418 238170 235488 238226
rect 235168 238102 235488 238170
rect 235168 238046 235238 238102
rect 235294 238046 235362 238102
rect 235418 238046 235488 238102
rect 235168 237978 235488 238046
rect 235168 237922 235238 237978
rect 235294 237922 235362 237978
rect 235418 237922 235488 237978
rect 235168 237888 235488 237922
rect 265888 238350 266208 238384
rect 265888 238294 265958 238350
rect 266014 238294 266082 238350
rect 266138 238294 266208 238350
rect 265888 238226 266208 238294
rect 265888 238170 265958 238226
rect 266014 238170 266082 238226
rect 266138 238170 266208 238226
rect 265888 238102 266208 238170
rect 265888 238046 265958 238102
rect 266014 238046 266082 238102
rect 266138 238046 266208 238102
rect 265888 237978 266208 238046
rect 265888 237922 265958 237978
rect 266014 237922 266082 237978
rect 266138 237922 266208 237978
rect 265888 237888 266208 237922
rect 296608 238350 296928 238384
rect 296608 238294 296678 238350
rect 296734 238294 296802 238350
rect 296858 238294 296928 238350
rect 296608 238226 296928 238294
rect 296608 238170 296678 238226
rect 296734 238170 296802 238226
rect 296858 238170 296928 238226
rect 296608 238102 296928 238170
rect 296608 238046 296678 238102
rect 296734 238046 296802 238102
rect 296858 238046 296928 238102
rect 296608 237978 296928 238046
rect 296608 237922 296678 237978
rect 296734 237922 296802 237978
rect 296858 237922 296928 237978
rect 296608 237888 296928 237922
rect 327328 238350 327648 238384
rect 327328 238294 327398 238350
rect 327454 238294 327522 238350
rect 327578 238294 327648 238350
rect 327328 238226 327648 238294
rect 327328 238170 327398 238226
rect 327454 238170 327522 238226
rect 327578 238170 327648 238226
rect 327328 238102 327648 238170
rect 327328 238046 327398 238102
rect 327454 238046 327522 238102
rect 327578 238046 327648 238102
rect 327328 237978 327648 238046
rect 327328 237922 327398 237978
rect 327454 237922 327522 237978
rect 327578 237922 327648 237978
rect 327328 237888 327648 237922
rect 358048 238350 358368 238384
rect 358048 238294 358118 238350
rect 358174 238294 358242 238350
rect 358298 238294 358368 238350
rect 358048 238226 358368 238294
rect 358048 238170 358118 238226
rect 358174 238170 358242 238226
rect 358298 238170 358368 238226
rect 358048 238102 358368 238170
rect 358048 238046 358118 238102
rect 358174 238046 358242 238102
rect 358298 238046 358368 238102
rect 358048 237978 358368 238046
rect 358048 237922 358118 237978
rect 358174 237922 358242 237978
rect 358298 237922 358368 237978
rect 358048 237888 358368 237922
rect 388768 238350 389088 238384
rect 388768 238294 388838 238350
rect 388894 238294 388962 238350
rect 389018 238294 389088 238350
rect 388768 238226 389088 238294
rect 388768 238170 388838 238226
rect 388894 238170 388962 238226
rect 389018 238170 389088 238226
rect 388768 238102 389088 238170
rect 388768 238046 388838 238102
rect 388894 238046 388962 238102
rect 389018 238046 389088 238102
rect 388768 237978 389088 238046
rect 388768 237922 388838 237978
rect 388894 237922 388962 237978
rect 389018 237922 389088 237978
rect 388768 237888 389088 237922
rect 419488 238350 419808 238384
rect 419488 238294 419558 238350
rect 419614 238294 419682 238350
rect 419738 238294 419808 238350
rect 419488 238226 419808 238294
rect 419488 238170 419558 238226
rect 419614 238170 419682 238226
rect 419738 238170 419808 238226
rect 419488 238102 419808 238170
rect 419488 238046 419558 238102
rect 419614 238046 419682 238102
rect 419738 238046 419808 238102
rect 419488 237978 419808 238046
rect 419488 237922 419558 237978
rect 419614 237922 419682 237978
rect 419738 237922 419808 237978
rect 419488 237888 419808 237922
rect 450208 238350 450528 238384
rect 450208 238294 450278 238350
rect 450334 238294 450402 238350
rect 450458 238294 450528 238350
rect 450208 238226 450528 238294
rect 450208 238170 450278 238226
rect 450334 238170 450402 238226
rect 450458 238170 450528 238226
rect 450208 238102 450528 238170
rect 450208 238046 450278 238102
rect 450334 238046 450402 238102
rect 450458 238046 450528 238102
rect 450208 237978 450528 238046
rect 450208 237922 450278 237978
rect 450334 237922 450402 237978
rect 450458 237922 450528 237978
rect 450208 237888 450528 237922
rect 480928 238350 481248 238384
rect 480928 238294 480998 238350
rect 481054 238294 481122 238350
rect 481178 238294 481248 238350
rect 480928 238226 481248 238294
rect 480928 238170 480998 238226
rect 481054 238170 481122 238226
rect 481178 238170 481248 238226
rect 480928 238102 481248 238170
rect 480928 238046 480998 238102
rect 481054 238046 481122 238102
rect 481178 238046 481248 238102
rect 480928 237978 481248 238046
rect 480928 237922 480998 237978
rect 481054 237922 481122 237978
rect 481178 237922 481248 237978
rect 480928 237888 481248 237922
rect 507154 238350 507774 255922
rect 507154 238294 507250 238350
rect 507306 238294 507374 238350
rect 507430 238294 507498 238350
rect 507554 238294 507622 238350
rect 507678 238294 507774 238350
rect 507154 238226 507774 238294
rect 507154 238170 507250 238226
rect 507306 238170 507374 238226
rect 507430 238170 507498 238226
rect 507554 238170 507622 238226
rect 507678 238170 507774 238226
rect 507154 238102 507774 238170
rect 507154 238046 507250 238102
rect 507306 238046 507374 238102
rect 507430 238046 507498 238102
rect 507554 238046 507622 238102
rect 507678 238046 507774 238102
rect 507154 237978 507774 238046
rect 507154 237922 507250 237978
rect 507306 237922 507374 237978
rect 507430 237922 507498 237978
rect 507554 237922 507622 237978
rect 507678 237922 507774 237978
rect 219808 226350 220128 226384
rect 219808 226294 219878 226350
rect 219934 226294 220002 226350
rect 220058 226294 220128 226350
rect 219808 226226 220128 226294
rect 219808 226170 219878 226226
rect 219934 226170 220002 226226
rect 220058 226170 220128 226226
rect 219808 226102 220128 226170
rect 219808 226046 219878 226102
rect 219934 226046 220002 226102
rect 220058 226046 220128 226102
rect 219808 225978 220128 226046
rect 219808 225922 219878 225978
rect 219934 225922 220002 225978
rect 220058 225922 220128 225978
rect 219808 225888 220128 225922
rect 250528 226350 250848 226384
rect 250528 226294 250598 226350
rect 250654 226294 250722 226350
rect 250778 226294 250848 226350
rect 250528 226226 250848 226294
rect 250528 226170 250598 226226
rect 250654 226170 250722 226226
rect 250778 226170 250848 226226
rect 250528 226102 250848 226170
rect 250528 226046 250598 226102
rect 250654 226046 250722 226102
rect 250778 226046 250848 226102
rect 250528 225978 250848 226046
rect 250528 225922 250598 225978
rect 250654 225922 250722 225978
rect 250778 225922 250848 225978
rect 250528 225888 250848 225922
rect 281248 226350 281568 226384
rect 281248 226294 281318 226350
rect 281374 226294 281442 226350
rect 281498 226294 281568 226350
rect 281248 226226 281568 226294
rect 281248 226170 281318 226226
rect 281374 226170 281442 226226
rect 281498 226170 281568 226226
rect 281248 226102 281568 226170
rect 281248 226046 281318 226102
rect 281374 226046 281442 226102
rect 281498 226046 281568 226102
rect 281248 225978 281568 226046
rect 281248 225922 281318 225978
rect 281374 225922 281442 225978
rect 281498 225922 281568 225978
rect 281248 225888 281568 225922
rect 311968 226350 312288 226384
rect 311968 226294 312038 226350
rect 312094 226294 312162 226350
rect 312218 226294 312288 226350
rect 311968 226226 312288 226294
rect 311968 226170 312038 226226
rect 312094 226170 312162 226226
rect 312218 226170 312288 226226
rect 311968 226102 312288 226170
rect 311968 226046 312038 226102
rect 312094 226046 312162 226102
rect 312218 226046 312288 226102
rect 311968 225978 312288 226046
rect 311968 225922 312038 225978
rect 312094 225922 312162 225978
rect 312218 225922 312288 225978
rect 311968 225888 312288 225922
rect 342688 226350 343008 226384
rect 342688 226294 342758 226350
rect 342814 226294 342882 226350
rect 342938 226294 343008 226350
rect 342688 226226 343008 226294
rect 342688 226170 342758 226226
rect 342814 226170 342882 226226
rect 342938 226170 343008 226226
rect 342688 226102 343008 226170
rect 342688 226046 342758 226102
rect 342814 226046 342882 226102
rect 342938 226046 343008 226102
rect 342688 225978 343008 226046
rect 342688 225922 342758 225978
rect 342814 225922 342882 225978
rect 342938 225922 343008 225978
rect 342688 225888 343008 225922
rect 373408 226350 373728 226384
rect 373408 226294 373478 226350
rect 373534 226294 373602 226350
rect 373658 226294 373728 226350
rect 373408 226226 373728 226294
rect 373408 226170 373478 226226
rect 373534 226170 373602 226226
rect 373658 226170 373728 226226
rect 373408 226102 373728 226170
rect 373408 226046 373478 226102
rect 373534 226046 373602 226102
rect 373658 226046 373728 226102
rect 373408 225978 373728 226046
rect 373408 225922 373478 225978
rect 373534 225922 373602 225978
rect 373658 225922 373728 225978
rect 373408 225888 373728 225922
rect 404128 226350 404448 226384
rect 404128 226294 404198 226350
rect 404254 226294 404322 226350
rect 404378 226294 404448 226350
rect 404128 226226 404448 226294
rect 404128 226170 404198 226226
rect 404254 226170 404322 226226
rect 404378 226170 404448 226226
rect 404128 226102 404448 226170
rect 404128 226046 404198 226102
rect 404254 226046 404322 226102
rect 404378 226046 404448 226102
rect 404128 225978 404448 226046
rect 404128 225922 404198 225978
rect 404254 225922 404322 225978
rect 404378 225922 404448 225978
rect 404128 225888 404448 225922
rect 434848 226350 435168 226384
rect 434848 226294 434918 226350
rect 434974 226294 435042 226350
rect 435098 226294 435168 226350
rect 434848 226226 435168 226294
rect 434848 226170 434918 226226
rect 434974 226170 435042 226226
rect 435098 226170 435168 226226
rect 434848 226102 435168 226170
rect 434848 226046 434918 226102
rect 434974 226046 435042 226102
rect 435098 226046 435168 226102
rect 434848 225978 435168 226046
rect 434848 225922 434918 225978
rect 434974 225922 435042 225978
rect 435098 225922 435168 225978
rect 434848 225888 435168 225922
rect 465568 226350 465888 226384
rect 465568 226294 465638 226350
rect 465694 226294 465762 226350
rect 465818 226294 465888 226350
rect 465568 226226 465888 226294
rect 465568 226170 465638 226226
rect 465694 226170 465762 226226
rect 465818 226170 465888 226226
rect 465568 226102 465888 226170
rect 465568 226046 465638 226102
rect 465694 226046 465762 226102
rect 465818 226046 465888 226102
rect 465568 225978 465888 226046
rect 465568 225922 465638 225978
rect 465694 225922 465762 225978
rect 465818 225922 465888 225978
rect 465568 225888 465888 225922
rect 496288 226350 496608 226384
rect 496288 226294 496358 226350
rect 496414 226294 496482 226350
rect 496538 226294 496608 226350
rect 496288 226226 496608 226294
rect 496288 226170 496358 226226
rect 496414 226170 496482 226226
rect 496538 226170 496608 226226
rect 496288 226102 496608 226170
rect 496288 226046 496358 226102
rect 496414 226046 496482 226102
rect 496538 226046 496608 226102
rect 496288 225978 496608 226046
rect 496288 225922 496358 225978
rect 496414 225922 496482 225978
rect 496538 225922 496608 225978
rect 496288 225888 496608 225922
rect 201154 220294 201250 220350
rect 201306 220294 201374 220350
rect 201430 220294 201498 220350
rect 201554 220294 201622 220350
rect 201678 220294 201774 220350
rect 201154 220226 201774 220294
rect 201154 220170 201250 220226
rect 201306 220170 201374 220226
rect 201430 220170 201498 220226
rect 201554 220170 201622 220226
rect 201678 220170 201774 220226
rect 201154 220102 201774 220170
rect 201154 220046 201250 220102
rect 201306 220046 201374 220102
rect 201430 220046 201498 220102
rect 201554 220046 201622 220102
rect 201678 220046 201774 220102
rect 201154 219978 201774 220046
rect 201154 219922 201250 219978
rect 201306 219922 201374 219978
rect 201430 219922 201498 219978
rect 201554 219922 201622 219978
rect 201678 219922 201774 219978
rect 201154 202350 201774 219922
rect 204448 220350 204768 220384
rect 204448 220294 204518 220350
rect 204574 220294 204642 220350
rect 204698 220294 204768 220350
rect 204448 220226 204768 220294
rect 204448 220170 204518 220226
rect 204574 220170 204642 220226
rect 204698 220170 204768 220226
rect 204448 220102 204768 220170
rect 204448 220046 204518 220102
rect 204574 220046 204642 220102
rect 204698 220046 204768 220102
rect 204448 219978 204768 220046
rect 204448 219922 204518 219978
rect 204574 219922 204642 219978
rect 204698 219922 204768 219978
rect 204448 219888 204768 219922
rect 235168 220350 235488 220384
rect 235168 220294 235238 220350
rect 235294 220294 235362 220350
rect 235418 220294 235488 220350
rect 235168 220226 235488 220294
rect 235168 220170 235238 220226
rect 235294 220170 235362 220226
rect 235418 220170 235488 220226
rect 235168 220102 235488 220170
rect 235168 220046 235238 220102
rect 235294 220046 235362 220102
rect 235418 220046 235488 220102
rect 235168 219978 235488 220046
rect 235168 219922 235238 219978
rect 235294 219922 235362 219978
rect 235418 219922 235488 219978
rect 235168 219888 235488 219922
rect 265888 220350 266208 220384
rect 265888 220294 265958 220350
rect 266014 220294 266082 220350
rect 266138 220294 266208 220350
rect 265888 220226 266208 220294
rect 265888 220170 265958 220226
rect 266014 220170 266082 220226
rect 266138 220170 266208 220226
rect 265888 220102 266208 220170
rect 265888 220046 265958 220102
rect 266014 220046 266082 220102
rect 266138 220046 266208 220102
rect 265888 219978 266208 220046
rect 265888 219922 265958 219978
rect 266014 219922 266082 219978
rect 266138 219922 266208 219978
rect 265888 219888 266208 219922
rect 296608 220350 296928 220384
rect 296608 220294 296678 220350
rect 296734 220294 296802 220350
rect 296858 220294 296928 220350
rect 296608 220226 296928 220294
rect 296608 220170 296678 220226
rect 296734 220170 296802 220226
rect 296858 220170 296928 220226
rect 296608 220102 296928 220170
rect 296608 220046 296678 220102
rect 296734 220046 296802 220102
rect 296858 220046 296928 220102
rect 296608 219978 296928 220046
rect 296608 219922 296678 219978
rect 296734 219922 296802 219978
rect 296858 219922 296928 219978
rect 296608 219888 296928 219922
rect 327328 220350 327648 220384
rect 327328 220294 327398 220350
rect 327454 220294 327522 220350
rect 327578 220294 327648 220350
rect 327328 220226 327648 220294
rect 327328 220170 327398 220226
rect 327454 220170 327522 220226
rect 327578 220170 327648 220226
rect 327328 220102 327648 220170
rect 327328 220046 327398 220102
rect 327454 220046 327522 220102
rect 327578 220046 327648 220102
rect 327328 219978 327648 220046
rect 327328 219922 327398 219978
rect 327454 219922 327522 219978
rect 327578 219922 327648 219978
rect 327328 219888 327648 219922
rect 358048 220350 358368 220384
rect 358048 220294 358118 220350
rect 358174 220294 358242 220350
rect 358298 220294 358368 220350
rect 358048 220226 358368 220294
rect 358048 220170 358118 220226
rect 358174 220170 358242 220226
rect 358298 220170 358368 220226
rect 358048 220102 358368 220170
rect 358048 220046 358118 220102
rect 358174 220046 358242 220102
rect 358298 220046 358368 220102
rect 358048 219978 358368 220046
rect 358048 219922 358118 219978
rect 358174 219922 358242 219978
rect 358298 219922 358368 219978
rect 358048 219888 358368 219922
rect 388768 220350 389088 220384
rect 388768 220294 388838 220350
rect 388894 220294 388962 220350
rect 389018 220294 389088 220350
rect 388768 220226 389088 220294
rect 388768 220170 388838 220226
rect 388894 220170 388962 220226
rect 389018 220170 389088 220226
rect 388768 220102 389088 220170
rect 388768 220046 388838 220102
rect 388894 220046 388962 220102
rect 389018 220046 389088 220102
rect 388768 219978 389088 220046
rect 388768 219922 388838 219978
rect 388894 219922 388962 219978
rect 389018 219922 389088 219978
rect 388768 219888 389088 219922
rect 419488 220350 419808 220384
rect 419488 220294 419558 220350
rect 419614 220294 419682 220350
rect 419738 220294 419808 220350
rect 419488 220226 419808 220294
rect 419488 220170 419558 220226
rect 419614 220170 419682 220226
rect 419738 220170 419808 220226
rect 419488 220102 419808 220170
rect 419488 220046 419558 220102
rect 419614 220046 419682 220102
rect 419738 220046 419808 220102
rect 419488 219978 419808 220046
rect 419488 219922 419558 219978
rect 419614 219922 419682 219978
rect 419738 219922 419808 219978
rect 419488 219888 419808 219922
rect 450208 220350 450528 220384
rect 450208 220294 450278 220350
rect 450334 220294 450402 220350
rect 450458 220294 450528 220350
rect 450208 220226 450528 220294
rect 450208 220170 450278 220226
rect 450334 220170 450402 220226
rect 450458 220170 450528 220226
rect 450208 220102 450528 220170
rect 450208 220046 450278 220102
rect 450334 220046 450402 220102
rect 450458 220046 450528 220102
rect 450208 219978 450528 220046
rect 450208 219922 450278 219978
rect 450334 219922 450402 219978
rect 450458 219922 450528 219978
rect 450208 219888 450528 219922
rect 480928 220350 481248 220384
rect 480928 220294 480998 220350
rect 481054 220294 481122 220350
rect 481178 220294 481248 220350
rect 480928 220226 481248 220294
rect 480928 220170 480998 220226
rect 481054 220170 481122 220226
rect 481178 220170 481248 220226
rect 480928 220102 481248 220170
rect 480928 220046 480998 220102
rect 481054 220046 481122 220102
rect 481178 220046 481248 220102
rect 480928 219978 481248 220046
rect 480928 219922 480998 219978
rect 481054 219922 481122 219978
rect 481178 219922 481248 219978
rect 480928 219888 481248 219922
rect 507154 220350 507774 237922
rect 507154 220294 507250 220350
rect 507306 220294 507374 220350
rect 507430 220294 507498 220350
rect 507554 220294 507622 220350
rect 507678 220294 507774 220350
rect 507154 220226 507774 220294
rect 507154 220170 507250 220226
rect 507306 220170 507374 220226
rect 507430 220170 507498 220226
rect 507554 220170 507622 220226
rect 507678 220170 507774 220226
rect 507154 220102 507774 220170
rect 507154 220046 507250 220102
rect 507306 220046 507374 220102
rect 507430 220046 507498 220102
rect 507554 220046 507622 220102
rect 507678 220046 507774 220102
rect 507154 219978 507774 220046
rect 507154 219922 507250 219978
rect 507306 219922 507374 219978
rect 507430 219922 507498 219978
rect 507554 219922 507622 219978
rect 507678 219922 507774 219978
rect 201154 202294 201250 202350
rect 201306 202294 201374 202350
rect 201430 202294 201498 202350
rect 201554 202294 201622 202350
rect 201678 202294 201774 202350
rect 201154 202226 201774 202294
rect 201154 202170 201250 202226
rect 201306 202170 201374 202226
rect 201430 202170 201498 202226
rect 201554 202170 201622 202226
rect 201678 202170 201774 202226
rect 201154 202102 201774 202170
rect 201154 202046 201250 202102
rect 201306 202046 201374 202102
rect 201430 202046 201498 202102
rect 201554 202046 201622 202102
rect 201678 202046 201774 202102
rect 201154 201978 201774 202046
rect 201154 201922 201250 201978
rect 201306 201922 201374 201978
rect 201430 201922 201498 201978
rect 201554 201922 201622 201978
rect 201678 201922 201774 201978
rect 201154 184350 201774 201922
rect 201154 184294 201250 184350
rect 201306 184294 201374 184350
rect 201430 184294 201498 184350
rect 201554 184294 201622 184350
rect 201678 184294 201774 184350
rect 201154 184226 201774 184294
rect 201154 184170 201250 184226
rect 201306 184170 201374 184226
rect 201430 184170 201498 184226
rect 201554 184170 201622 184226
rect 201678 184170 201774 184226
rect 201154 184102 201774 184170
rect 201154 184046 201250 184102
rect 201306 184046 201374 184102
rect 201430 184046 201498 184102
rect 201554 184046 201622 184102
rect 201678 184046 201774 184102
rect 201154 183978 201774 184046
rect 201154 183922 201250 183978
rect 201306 183922 201374 183978
rect 201430 183922 201498 183978
rect 201554 183922 201622 183978
rect 201678 183922 201774 183978
rect 201154 166350 201774 183922
rect 201154 166294 201250 166350
rect 201306 166294 201374 166350
rect 201430 166294 201498 166350
rect 201554 166294 201622 166350
rect 201678 166294 201774 166350
rect 201154 166226 201774 166294
rect 201154 166170 201250 166226
rect 201306 166170 201374 166226
rect 201430 166170 201498 166226
rect 201554 166170 201622 166226
rect 201678 166170 201774 166226
rect 201154 166102 201774 166170
rect 201154 166046 201250 166102
rect 201306 166046 201374 166102
rect 201430 166046 201498 166102
rect 201554 166046 201622 166102
rect 201678 166046 201774 166102
rect 201154 165978 201774 166046
rect 201154 165922 201250 165978
rect 201306 165922 201374 165978
rect 201430 165922 201498 165978
rect 201554 165922 201622 165978
rect 201678 165922 201774 165978
rect 201154 148350 201774 165922
rect 201154 148294 201250 148350
rect 201306 148294 201374 148350
rect 201430 148294 201498 148350
rect 201554 148294 201622 148350
rect 201678 148294 201774 148350
rect 201154 148226 201774 148294
rect 201154 148170 201250 148226
rect 201306 148170 201374 148226
rect 201430 148170 201498 148226
rect 201554 148170 201622 148226
rect 201678 148170 201774 148226
rect 201154 148102 201774 148170
rect 201154 148046 201250 148102
rect 201306 148046 201374 148102
rect 201430 148046 201498 148102
rect 201554 148046 201622 148102
rect 201678 148046 201774 148102
rect 201154 147978 201774 148046
rect 201154 147922 201250 147978
rect 201306 147922 201374 147978
rect 201430 147922 201498 147978
rect 201554 147922 201622 147978
rect 201678 147922 201774 147978
rect 201154 130350 201774 147922
rect 201154 130294 201250 130350
rect 201306 130294 201374 130350
rect 201430 130294 201498 130350
rect 201554 130294 201622 130350
rect 201678 130294 201774 130350
rect 201154 130226 201774 130294
rect 201154 130170 201250 130226
rect 201306 130170 201374 130226
rect 201430 130170 201498 130226
rect 201554 130170 201622 130226
rect 201678 130170 201774 130226
rect 201154 130102 201774 130170
rect 201154 130046 201250 130102
rect 201306 130046 201374 130102
rect 201430 130046 201498 130102
rect 201554 130046 201622 130102
rect 201678 130046 201774 130102
rect 201154 129978 201774 130046
rect 201154 129922 201250 129978
rect 201306 129922 201374 129978
rect 201430 129922 201498 129978
rect 201554 129922 201622 129978
rect 201678 129922 201774 129978
rect 201154 112350 201774 129922
rect 201154 112294 201250 112350
rect 201306 112294 201374 112350
rect 201430 112294 201498 112350
rect 201554 112294 201622 112350
rect 201678 112294 201774 112350
rect 201154 112226 201774 112294
rect 201154 112170 201250 112226
rect 201306 112170 201374 112226
rect 201430 112170 201498 112226
rect 201554 112170 201622 112226
rect 201678 112170 201774 112226
rect 201154 112102 201774 112170
rect 201154 112046 201250 112102
rect 201306 112046 201374 112102
rect 201430 112046 201498 112102
rect 201554 112046 201622 112102
rect 201678 112046 201774 112102
rect 201154 111978 201774 112046
rect 201154 111922 201250 111978
rect 201306 111922 201374 111978
rect 201430 111922 201498 111978
rect 201554 111922 201622 111978
rect 201678 111922 201774 111978
rect 201154 94350 201774 111922
rect 201154 94294 201250 94350
rect 201306 94294 201374 94350
rect 201430 94294 201498 94350
rect 201554 94294 201622 94350
rect 201678 94294 201774 94350
rect 201154 94226 201774 94294
rect 201154 94170 201250 94226
rect 201306 94170 201374 94226
rect 201430 94170 201498 94226
rect 201554 94170 201622 94226
rect 201678 94170 201774 94226
rect 201154 94102 201774 94170
rect 201154 94046 201250 94102
rect 201306 94046 201374 94102
rect 201430 94046 201498 94102
rect 201554 94046 201622 94102
rect 201678 94046 201774 94102
rect 201154 93978 201774 94046
rect 201154 93922 201250 93978
rect 201306 93922 201374 93978
rect 201430 93922 201498 93978
rect 201554 93922 201622 93978
rect 201678 93922 201774 93978
rect 201154 76350 201774 93922
rect 201154 76294 201250 76350
rect 201306 76294 201374 76350
rect 201430 76294 201498 76350
rect 201554 76294 201622 76350
rect 201678 76294 201774 76350
rect 201154 76226 201774 76294
rect 201154 76170 201250 76226
rect 201306 76170 201374 76226
rect 201430 76170 201498 76226
rect 201554 76170 201622 76226
rect 201678 76170 201774 76226
rect 201154 76102 201774 76170
rect 201154 76046 201250 76102
rect 201306 76046 201374 76102
rect 201430 76046 201498 76102
rect 201554 76046 201622 76102
rect 201678 76046 201774 76102
rect 201154 75978 201774 76046
rect 201154 75922 201250 75978
rect 201306 75922 201374 75978
rect 201430 75922 201498 75978
rect 201554 75922 201622 75978
rect 201678 75922 201774 75978
rect 201154 58350 201774 75922
rect 201154 58294 201250 58350
rect 201306 58294 201374 58350
rect 201430 58294 201498 58350
rect 201554 58294 201622 58350
rect 201678 58294 201774 58350
rect 201154 58226 201774 58294
rect 201154 58170 201250 58226
rect 201306 58170 201374 58226
rect 201430 58170 201498 58226
rect 201554 58170 201622 58226
rect 201678 58170 201774 58226
rect 201154 58102 201774 58170
rect 201154 58046 201250 58102
rect 201306 58046 201374 58102
rect 201430 58046 201498 58102
rect 201554 58046 201622 58102
rect 201678 58046 201774 58102
rect 201154 57978 201774 58046
rect 201154 57922 201250 57978
rect 201306 57922 201374 57978
rect 201430 57922 201498 57978
rect 201554 57922 201622 57978
rect 201678 57922 201774 57978
rect 201154 40350 201774 57922
rect 201154 40294 201250 40350
rect 201306 40294 201374 40350
rect 201430 40294 201498 40350
rect 201554 40294 201622 40350
rect 201678 40294 201774 40350
rect 201154 40226 201774 40294
rect 201154 40170 201250 40226
rect 201306 40170 201374 40226
rect 201430 40170 201498 40226
rect 201554 40170 201622 40226
rect 201678 40170 201774 40226
rect 201154 40102 201774 40170
rect 201154 40046 201250 40102
rect 201306 40046 201374 40102
rect 201430 40046 201498 40102
rect 201554 40046 201622 40102
rect 201678 40046 201774 40102
rect 201154 39978 201774 40046
rect 201154 39922 201250 39978
rect 201306 39922 201374 39978
rect 201430 39922 201498 39978
rect 201554 39922 201622 39978
rect 201678 39922 201774 39978
rect 201154 22350 201774 39922
rect 201154 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 201774 22350
rect 201154 22226 201774 22294
rect 201154 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 201774 22226
rect 201154 22102 201774 22170
rect 201154 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 201774 22102
rect 201154 21978 201774 22046
rect 201154 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 201774 21978
rect 201154 4350 201774 21922
rect 201154 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 201774 4350
rect 201154 4226 201774 4294
rect 201154 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 201774 4226
rect 201154 4102 201774 4170
rect 201154 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 201774 4102
rect 201154 3978 201774 4046
rect 201154 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 201774 3978
rect 201154 -160 201774 3922
rect 201154 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 201774 -160
rect 201154 -284 201774 -216
rect 201154 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 201774 -284
rect 201154 -408 201774 -340
rect 201154 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 201774 -408
rect 201154 -532 201774 -464
rect 201154 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 201774 -532
rect 201154 -1644 201774 -588
rect 204874 208350 205494 210842
rect 204874 208294 204970 208350
rect 205026 208294 205094 208350
rect 205150 208294 205218 208350
rect 205274 208294 205342 208350
rect 205398 208294 205494 208350
rect 204874 208226 205494 208294
rect 204874 208170 204970 208226
rect 205026 208170 205094 208226
rect 205150 208170 205218 208226
rect 205274 208170 205342 208226
rect 205398 208170 205494 208226
rect 204874 208102 205494 208170
rect 204874 208046 204970 208102
rect 205026 208046 205094 208102
rect 205150 208046 205218 208102
rect 205274 208046 205342 208102
rect 205398 208046 205494 208102
rect 204874 207978 205494 208046
rect 204874 207922 204970 207978
rect 205026 207922 205094 207978
rect 205150 207922 205218 207978
rect 205274 207922 205342 207978
rect 205398 207922 205494 207978
rect 204874 190350 205494 207922
rect 219808 208350 220128 208384
rect 219808 208294 219878 208350
rect 219934 208294 220002 208350
rect 220058 208294 220128 208350
rect 219808 208226 220128 208294
rect 219808 208170 219878 208226
rect 219934 208170 220002 208226
rect 220058 208170 220128 208226
rect 219808 208102 220128 208170
rect 219808 208046 219878 208102
rect 219934 208046 220002 208102
rect 220058 208046 220128 208102
rect 219808 207978 220128 208046
rect 219808 207922 219878 207978
rect 219934 207922 220002 207978
rect 220058 207922 220128 207978
rect 219808 207888 220128 207922
rect 222874 208350 223494 210842
rect 222874 208294 222970 208350
rect 223026 208294 223094 208350
rect 223150 208294 223218 208350
rect 223274 208294 223342 208350
rect 223398 208294 223494 208350
rect 222874 208226 223494 208294
rect 222874 208170 222970 208226
rect 223026 208170 223094 208226
rect 223150 208170 223218 208226
rect 223274 208170 223342 208226
rect 223398 208170 223494 208226
rect 222874 208102 223494 208170
rect 222874 208046 222970 208102
rect 223026 208046 223094 208102
rect 223150 208046 223218 208102
rect 223274 208046 223342 208102
rect 223398 208046 223494 208102
rect 222874 207978 223494 208046
rect 222874 207922 222970 207978
rect 223026 207922 223094 207978
rect 223150 207922 223218 207978
rect 223274 207922 223342 207978
rect 223398 207922 223494 207978
rect 204874 190294 204970 190350
rect 205026 190294 205094 190350
rect 205150 190294 205218 190350
rect 205274 190294 205342 190350
rect 205398 190294 205494 190350
rect 204874 190226 205494 190294
rect 204874 190170 204970 190226
rect 205026 190170 205094 190226
rect 205150 190170 205218 190226
rect 205274 190170 205342 190226
rect 205398 190170 205494 190226
rect 204874 190102 205494 190170
rect 204874 190046 204970 190102
rect 205026 190046 205094 190102
rect 205150 190046 205218 190102
rect 205274 190046 205342 190102
rect 205398 190046 205494 190102
rect 204874 189978 205494 190046
rect 204874 189922 204970 189978
rect 205026 189922 205094 189978
rect 205150 189922 205218 189978
rect 205274 189922 205342 189978
rect 205398 189922 205494 189978
rect 204874 172350 205494 189922
rect 204874 172294 204970 172350
rect 205026 172294 205094 172350
rect 205150 172294 205218 172350
rect 205274 172294 205342 172350
rect 205398 172294 205494 172350
rect 204874 172226 205494 172294
rect 204874 172170 204970 172226
rect 205026 172170 205094 172226
rect 205150 172170 205218 172226
rect 205274 172170 205342 172226
rect 205398 172170 205494 172226
rect 204874 172102 205494 172170
rect 204874 172046 204970 172102
rect 205026 172046 205094 172102
rect 205150 172046 205218 172102
rect 205274 172046 205342 172102
rect 205398 172046 205494 172102
rect 204874 171978 205494 172046
rect 204874 171922 204970 171978
rect 205026 171922 205094 171978
rect 205150 171922 205218 171978
rect 205274 171922 205342 171978
rect 205398 171922 205494 171978
rect 204874 154350 205494 171922
rect 204874 154294 204970 154350
rect 205026 154294 205094 154350
rect 205150 154294 205218 154350
rect 205274 154294 205342 154350
rect 205398 154294 205494 154350
rect 204874 154226 205494 154294
rect 204874 154170 204970 154226
rect 205026 154170 205094 154226
rect 205150 154170 205218 154226
rect 205274 154170 205342 154226
rect 205398 154170 205494 154226
rect 204874 154102 205494 154170
rect 204874 154046 204970 154102
rect 205026 154046 205094 154102
rect 205150 154046 205218 154102
rect 205274 154046 205342 154102
rect 205398 154046 205494 154102
rect 204874 153978 205494 154046
rect 204874 153922 204970 153978
rect 205026 153922 205094 153978
rect 205150 153922 205218 153978
rect 205274 153922 205342 153978
rect 205398 153922 205494 153978
rect 204874 136350 205494 153922
rect 204874 136294 204970 136350
rect 205026 136294 205094 136350
rect 205150 136294 205218 136350
rect 205274 136294 205342 136350
rect 205398 136294 205494 136350
rect 204874 136226 205494 136294
rect 204874 136170 204970 136226
rect 205026 136170 205094 136226
rect 205150 136170 205218 136226
rect 205274 136170 205342 136226
rect 205398 136170 205494 136226
rect 204874 136102 205494 136170
rect 204874 136046 204970 136102
rect 205026 136046 205094 136102
rect 205150 136046 205218 136102
rect 205274 136046 205342 136102
rect 205398 136046 205494 136102
rect 204874 135978 205494 136046
rect 204874 135922 204970 135978
rect 205026 135922 205094 135978
rect 205150 135922 205218 135978
rect 205274 135922 205342 135978
rect 205398 135922 205494 135978
rect 204874 118350 205494 135922
rect 204874 118294 204970 118350
rect 205026 118294 205094 118350
rect 205150 118294 205218 118350
rect 205274 118294 205342 118350
rect 205398 118294 205494 118350
rect 204874 118226 205494 118294
rect 204874 118170 204970 118226
rect 205026 118170 205094 118226
rect 205150 118170 205218 118226
rect 205274 118170 205342 118226
rect 205398 118170 205494 118226
rect 204874 118102 205494 118170
rect 204874 118046 204970 118102
rect 205026 118046 205094 118102
rect 205150 118046 205218 118102
rect 205274 118046 205342 118102
rect 205398 118046 205494 118102
rect 204874 117978 205494 118046
rect 204874 117922 204970 117978
rect 205026 117922 205094 117978
rect 205150 117922 205218 117978
rect 205274 117922 205342 117978
rect 205398 117922 205494 117978
rect 204874 100350 205494 117922
rect 204874 100294 204970 100350
rect 205026 100294 205094 100350
rect 205150 100294 205218 100350
rect 205274 100294 205342 100350
rect 205398 100294 205494 100350
rect 204874 100226 205494 100294
rect 204874 100170 204970 100226
rect 205026 100170 205094 100226
rect 205150 100170 205218 100226
rect 205274 100170 205342 100226
rect 205398 100170 205494 100226
rect 204874 100102 205494 100170
rect 204874 100046 204970 100102
rect 205026 100046 205094 100102
rect 205150 100046 205218 100102
rect 205274 100046 205342 100102
rect 205398 100046 205494 100102
rect 204874 99978 205494 100046
rect 204874 99922 204970 99978
rect 205026 99922 205094 99978
rect 205150 99922 205218 99978
rect 205274 99922 205342 99978
rect 205398 99922 205494 99978
rect 204874 82350 205494 99922
rect 204874 82294 204970 82350
rect 205026 82294 205094 82350
rect 205150 82294 205218 82350
rect 205274 82294 205342 82350
rect 205398 82294 205494 82350
rect 204874 82226 205494 82294
rect 204874 82170 204970 82226
rect 205026 82170 205094 82226
rect 205150 82170 205218 82226
rect 205274 82170 205342 82226
rect 205398 82170 205494 82226
rect 204874 82102 205494 82170
rect 204874 82046 204970 82102
rect 205026 82046 205094 82102
rect 205150 82046 205218 82102
rect 205274 82046 205342 82102
rect 205398 82046 205494 82102
rect 204874 81978 205494 82046
rect 204874 81922 204970 81978
rect 205026 81922 205094 81978
rect 205150 81922 205218 81978
rect 205274 81922 205342 81978
rect 205398 81922 205494 81978
rect 204874 64350 205494 81922
rect 204874 64294 204970 64350
rect 205026 64294 205094 64350
rect 205150 64294 205218 64350
rect 205274 64294 205342 64350
rect 205398 64294 205494 64350
rect 204874 64226 205494 64294
rect 204874 64170 204970 64226
rect 205026 64170 205094 64226
rect 205150 64170 205218 64226
rect 205274 64170 205342 64226
rect 205398 64170 205494 64226
rect 204874 64102 205494 64170
rect 204874 64046 204970 64102
rect 205026 64046 205094 64102
rect 205150 64046 205218 64102
rect 205274 64046 205342 64102
rect 205398 64046 205494 64102
rect 204874 63978 205494 64046
rect 204874 63922 204970 63978
rect 205026 63922 205094 63978
rect 205150 63922 205218 63978
rect 205274 63922 205342 63978
rect 205398 63922 205494 63978
rect 204874 46350 205494 63922
rect 204874 46294 204970 46350
rect 205026 46294 205094 46350
rect 205150 46294 205218 46350
rect 205274 46294 205342 46350
rect 205398 46294 205494 46350
rect 204874 46226 205494 46294
rect 204874 46170 204970 46226
rect 205026 46170 205094 46226
rect 205150 46170 205218 46226
rect 205274 46170 205342 46226
rect 205398 46170 205494 46226
rect 204874 46102 205494 46170
rect 204874 46046 204970 46102
rect 205026 46046 205094 46102
rect 205150 46046 205218 46102
rect 205274 46046 205342 46102
rect 205398 46046 205494 46102
rect 204874 45978 205494 46046
rect 204874 45922 204970 45978
rect 205026 45922 205094 45978
rect 205150 45922 205218 45978
rect 205274 45922 205342 45978
rect 205398 45922 205494 45978
rect 204874 28350 205494 45922
rect 204874 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 205494 28350
rect 204874 28226 205494 28294
rect 204874 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 205494 28226
rect 204874 28102 205494 28170
rect 204874 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 205494 28102
rect 204874 27978 205494 28046
rect 204874 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 205494 27978
rect 204874 10350 205494 27922
rect 204874 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 205494 10350
rect 204874 10226 205494 10294
rect 204874 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 205494 10226
rect 204874 10102 205494 10170
rect 204874 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 205494 10102
rect 204874 9978 205494 10046
rect 204874 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 205494 9978
rect 204874 -1120 205494 9922
rect 204874 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 205494 -1120
rect 204874 -1244 205494 -1176
rect 204874 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 205494 -1244
rect 204874 -1368 205494 -1300
rect 204874 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 205494 -1368
rect 204874 -1492 205494 -1424
rect 204874 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 205494 -1492
rect 204874 -1644 205494 -1548
rect 219154 184350 219774 201020
rect 219154 184294 219250 184350
rect 219306 184294 219374 184350
rect 219430 184294 219498 184350
rect 219554 184294 219622 184350
rect 219678 184294 219774 184350
rect 219154 184226 219774 184294
rect 219154 184170 219250 184226
rect 219306 184170 219374 184226
rect 219430 184170 219498 184226
rect 219554 184170 219622 184226
rect 219678 184170 219774 184226
rect 219154 184102 219774 184170
rect 219154 184046 219250 184102
rect 219306 184046 219374 184102
rect 219430 184046 219498 184102
rect 219554 184046 219622 184102
rect 219678 184046 219774 184102
rect 219154 183978 219774 184046
rect 219154 183922 219250 183978
rect 219306 183922 219374 183978
rect 219430 183922 219498 183978
rect 219554 183922 219622 183978
rect 219678 183922 219774 183978
rect 219154 166350 219774 183922
rect 219154 166294 219250 166350
rect 219306 166294 219374 166350
rect 219430 166294 219498 166350
rect 219554 166294 219622 166350
rect 219678 166294 219774 166350
rect 219154 166226 219774 166294
rect 219154 166170 219250 166226
rect 219306 166170 219374 166226
rect 219430 166170 219498 166226
rect 219554 166170 219622 166226
rect 219678 166170 219774 166226
rect 219154 166102 219774 166170
rect 219154 166046 219250 166102
rect 219306 166046 219374 166102
rect 219430 166046 219498 166102
rect 219554 166046 219622 166102
rect 219678 166046 219774 166102
rect 219154 165978 219774 166046
rect 219154 165922 219250 165978
rect 219306 165922 219374 165978
rect 219430 165922 219498 165978
rect 219554 165922 219622 165978
rect 219678 165922 219774 165978
rect 219154 148350 219774 165922
rect 219154 148294 219250 148350
rect 219306 148294 219374 148350
rect 219430 148294 219498 148350
rect 219554 148294 219622 148350
rect 219678 148294 219774 148350
rect 219154 148226 219774 148294
rect 219154 148170 219250 148226
rect 219306 148170 219374 148226
rect 219430 148170 219498 148226
rect 219554 148170 219622 148226
rect 219678 148170 219774 148226
rect 219154 148102 219774 148170
rect 219154 148046 219250 148102
rect 219306 148046 219374 148102
rect 219430 148046 219498 148102
rect 219554 148046 219622 148102
rect 219678 148046 219774 148102
rect 219154 147978 219774 148046
rect 219154 147922 219250 147978
rect 219306 147922 219374 147978
rect 219430 147922 219498 147978
rect 219554 147922 219622 147978
rect 219678 147922 219774 147978
rect 219154 130350 219774 147922
rect 219154 130294 219250 130350
rect 219306 130294 219374 130350
rect 219430 130294 219498 130350
rect 219554 130294 219622 130350
rect 219678 130294 219774 130350
rect 219154 130226 219774 130294
rect 219154 130170 219250 130226
rect 219306 130170 219374 130226
rect 219430 130170 219498 130226
rect 219554 130170 219622 130226
rect 219678 130170 219774 130226
rect 219154 130102 219774 130170
rect 219154 130046 219250 130102
rect 219306 130046 219374 130102
rect 219430 130046 219498 130102
rect 219554 130046 219622 130102
rect 219678 130046 219774 130102
rect 219154 129978 219774 130046
rect 219154 129922 219250 129978
rect 219306 129922 219374 129978
rect 219430 129922 219498 129978
rect 219554 129922 219622 129978
rect 219678 129922 219774 129978
rect 219154 112350 219774 129922
rect 219154 112294 219250 112350
rect 219306 112294 219374 112350
rect 219430 112294 219498 112350
rect 219554 112294 219622 112350
rect 219678 112294 219774 112350
rect 219154 112226 219774 112294
rect 219154 112170 219250 112226
rect 219306 112170 219374 112226
rect 219430 112170 219498 112226
rect 219554 112170 219622 112226
rect 219678 112170 219774 112226
rect 219154 112102 219774 112170
rect 219154 112046 219250 112102
rect 219306 112046 219374 112102
rect 219430 112046 219498 112102
rect 219554 112046 219622 112102
rect 219678 112046 219774 112102
rect 219154 111978 219774 112046
rect 219154 111922 219250 111978
rect 219306 111922 219374 111978
rect 219430 111922 219498 111978
rect 219554 111922 219622 111978
rect 219678 111922 219774 111978
rect 219154 94350 219774 111922
rect 219154 94294 219250 94350
rect 219306 94294 219374 94350
rect 219430 94294 219498 94350
rect 219554 94294 219622 94350
rect 219678 94294 219774 94350
rect 219154 94226 219774 94294
rect 219154 94170 219250 94226
rect 219306 94170 219374 94226
rect 219430 94170 219498 94226
rect 219554 94170 219622 94226
rect 219678 94170 219774 94226
rect 219154 94102 219774 94170
rect 219154 94046 219250 94102
rect 219306 94046 219374 94102
rect 219430 94046 219498 94102
rect 219554 94046 219622 94102
rect 219678 94046 219774 94102
rect 219154 93978 219774 94046
rect 219154 93922 219250 93978
rect 219306 93922 219374 93978
rect 219430 93922 219498 93978
rect 219554 93922 219622 93978
rect 219678 93922 219774 93978
rect 219154 76350 219774 93922
rect 219154 76294 219250 76350
rect 219306 76294 219374 76350
rect 219430 76294 219498 76350
rect 219554 76294 219622 76350
rect 219678 76294 219774 76350
rect 219154 76226 219774 76294
rect 219154 76170 219250 76226
rect 219306 76170 219374 76226
rect 219430 76170 219498 76226
rect 219554 76170 219622 76226
rect 219678 76170 219774 76226
rect 219154 76102 219774 76170
rect 219154 76046 219250 76102
rect 219306 76046 219374 76102
rect 219430 76046 219498 76102
rect 219554 76046 219622 76102
rect 219678 76046 219774 76102
rect 219154 75978 219774 76046
rect 219154 75922 219250 75978
rect 219306 75922 219374 75978
rect 219430 75922 219498 75978
rect 219554 75922 219622 75978
rect 219678 75922 219774 75978
rect 219154 58350 219774 75922
rect 219154 58294 219250 58350
rect 219306 58294 219374 58350
rect 219430 58294 219498 58350
rect 219554 58294 219622 58350
rect 219678 58294 219774 58350
rect 219154 58226 219774 58294
rect 219154 58170 219250 58226
rect 219306 58170 219374 58226
rect 219430 58170 219498 58226
rect 219554 58170 219622 58226
rect 219678 58170 219774 58226
rect 219154 58102 219774 58170
rect 219154 58046 219250 58102
rect 219306 58046 219374 58102
rect 219430 58046 219498 58102
rect 219554 58046 219622 58102
rect 219678 58046 219774 58102
rect 219154 57978 219774 58046
rect 219154 57922 219250 57978
rect 219306 57922 219374 57978
rect 219430 57922 219498 57978
rect 219554 57922 219622 57978
rect 219678 57922 219774 57978
rect 219154 40350 219774 57922
rect 219154 40294 219250 40350
rect 219306 40294 219374 40350
rect 219430 40294 219498 40350
rect 219554 40294 219622 40350
rect 219678 40294 219774 40350
rect 219154 40226 219774 40294
rect 219154 40170 219250 40226
rect 219306 40170 219374 40226
rect 219430 40170 219498 40226
rect 219554 40170 219622 40226
rect 219678 40170 219774 40226
rect 219154 40102 219774 40170
rect 219154 40046 219250 40102
rect 219306 40046 219374 40102
rect 219430 40046 219498 40102
rect 219554 40046 219622 40102
rect 219678 40046 219774 40102
rect 219154 39978 219774 40046
rect 219154 39922 219250 39978
rect 219306 39922 219374 39978
rect 219430 39922 219498 39978
rect 219554 39922 219622 39978
rect 219678 39922 219774 39978
rect 219154 22350 219774 39922
rect 219154 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 219774 22350
rect 219154 22226 219774 22294
rect 219154 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 219774 22226
rect 219154 22102 219774 22170
rect 219154 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 219774 22102
rect 219154 21978 219774 22046
rect 219154 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 219774 21978
rect 219154 4350 219774 21922
rect 219154 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 219774 4350
rect 219154 4226 219774 4294
rect 219154 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 219774 4226
rect 219154 4102 219774 4170
rect 219154 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 219774 4102
rect 219154 3978 219774 4046
rect 219154 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 219774 3978
rect 219154 -160 219774 3922
rect 219154 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 219774 -160
rect 219154 -284 219774 -216
rect 219154 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 219774 -284
rect 219154 -408 219774 -340
rect 219154 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 219774 -408
rect 219154 -532 219774 -464
rect 219154 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 219774 -532
rect 219154 -1644 219774 -588
rect 222874 190350 223494 207922
rect 222874 190294 222970 190350
rect 223026 190294 223094 190350
rect 223150 190294 223218 190350
rect 223274 190294 223342 190350
rect 223398 190294 223494 190350
rect 222874 190226 223494 190294
rect 222874 190170 222970 190226
rect 223026 190170 223094 190226
rect 223150 190170 223218 190226
rect 223274 190170 223342 190226
rect 223398 190170 223494 190226
rect 222874 190102 223494 190170
rect 222874 190046 222970 190102
rect 223026 190046 223094 190102
rect 223150 190046 223218 190102
rect 223274 190046 223342 190102
rect 223398 190046 223494 190102
rect 222874 189978 223494 190046
rect 222874 189922 222970 189978
rect 223026 189922 223094 189978
rect 223150 189922 223218 189978
rect 223274 189922 223342 189978
rect 223398 189922 223494 189978
rect 222874 172350 223494 189922
rect 222874 172294 222970 172350
rect 223026 172294 223094 172350
rect 223150 172294 223218 172350
rect 223274 172294 223342 172350
rect 223398 172294 223494 172350
rect 222874 172226 223494 172294
rect 222874 172170 222970 172226
rect 223026 172170 223094 172226
rect 223150 172170 223218 172226
rect 223274 172170 223342 172226
rect 223398 172170 223494 172226
rect 222874 172102 223494 172170
rect 222874 172046 222970 172102
rect 223026 172046 223094 172102
rect 223150 172046 223218 172102
rect 223274 172046 223342 172102
rect 223398 172046 223494 172102
rect 222874 171978 223494 172046
rect 222874 171922 222970 171978
rect 223026 171922 223094 171978
rect 223150 171922 223218 171978
rect 223274 171922 223342 171978
rect 223398 171922 223494 171978
rect 222874 154350 223494 171922
rect 222874 154294 222970 154350
rect 223026 154294 223094 154350
rect 223150 154294 223218 154350
rect 223274 154294 223342 154350
rect 223398 154294 223494 154350
rect 222874 154226 223494 154294
rect 222874 154170 222970 154226
rect 223026 154170 223094 154226
rect 223150 154170 223218 154226
rect 223274 154170 223342 154226
rect 223398 154170 223494 154226
rect 222874 154102 223494 154170
rect 222874 154046 222970 154102
rect 223026 154046 223094 154102
rect 223150 154046 223218 154102
rect 223274 154046 223342 154102
rect 223398 154046 223494 154102
rect 222874 153978 223494 154046
rect 222874 153922 222970 153978
rect 223026 153922 223094 153978
rect 223150 153922 223218 153978
rect 223274 153922 223342 153978
rect 223398 153922 223494 153978
rect 222874 136350 223494 153922
rect 222874 136294 222970 136350
rect 223026 136294 223094 136350
rect 223150 136294 223218 136350
rect 223274 136294 223342 136350
rect 223398 136294 223494 136350
rect 222874 136226 223494 136294
rect 222874 136170 222970 136226
rect 223026 136170 223094 136226
rect 223150 136170 223218 136226
rect 223274 136170 223342 136226
rect 223398 136170 223494 136226
rect 222874 136102 223494 136170
rect 222874 136046 222970 136102
rect 223026 136046 223094 136102
rect 223150 136046 223218 136102
rect 223274 136046 223342 136102
rect 223398 136046 223494 136102
rect 222874 135978 223494 136046
rect 222874 135922 222970 135978
rect 223026 135922 223094 135978
rect 223150 135922 223218 135978
rect 223274 135922 223342 135978
rect 223398 135922 223494 135978
rect 222874 118350 223494 135922
rect 222874 118294 222970 118350
rect 223026 118294 223094 118350
rect 223150 118294 223218 118350
rect 223274 118294 223342 118350
rect 223398 118294 223494 118350
rect 222874 118226 223494 118294
rect 222874 118170 222970 118226
rect 223026 118170 223094 118226
rect 223150 118170 223218 118226
rect 223274 118170 223342 118226
rect 223398 118170 223494 118226
rect 222874 118102 223494 118170
rect 222874 118046 222970 118102
rect 223026 118046 223094 118102
rect 223150 118046 223218 118102
rect 223274 118046 223342 118102
rect 223398 118046 223494 118102
rect 222874 117978 223494 118046
rect 222874 117922 222970 117978
rect 223026 117922 223094 117978
rect 223150 117922 223218 117978
rect 223274 117922 223342 117978
rect 223398 117922 223494 117978
rect 222874 100350 223494 117922
rect 222874 100294 222970 100350
rect 223026 100294 223094 100350
rect 223150 100294 223218 100350
rect 223274 100294 223342 100350
rect 223398 100294 223494 100350
rect 222874 100226 223494 100294
rect 222874 100170 222970 100226
rect 223026 100170 223094 100226
rect 223150 100170 223218 100226
rect 223274 100170 223342 100226
rect 223398 100170 223494 100226
rect 222874 100102 223494 100170
rect 222874 100046 222970 100102
rect 223026 100046 223094 100102
rect 223150 100046 223218 100102
rect 223274 100046 223342 100102
rect 223398 100046 223494 100102
rect 222874 99978 223494 100046
rect 222874 99922 222970 99978
rect 223026 99922 223094 99978
rect 223150 99922 223218 99978
rect 223274 99922 223342 99978
rect 223398 99922 223494 99978
rect 222874 82350 223494 99922
rect 222874 82294 222970 82350
rect 223026 82294 223094 82350
rect 223150 82294 223218 82350
rect 223274 82294 223342 82350
rect 223398 82294 223494 82350
rect 222874 82226 223494 82294
rect 222874 82170 222970 82226
rect 223026 82170 223094 82226
rect 223150 82170 223218 82226
rect 223274 82170 223342 82226
rect 223398 82170 223494 82226
rect 222874 82102 223494 82170
rect 222874 82046 222970 82102
rect 223026 82046 223094 82102
rect 223150 82046 223218 82102
rect 223274 82046 223342 82102
rect 223398 82046 223494 82102
rect 222874 81978 223494 82046
rect 222874 81922 222970 81978
rect 223026 81922 223094 81978
rect 223150 81922 223218 81978
rect 223274 81922 223342 81978
rect 223398 81922 223494 81978
rect 222874 64350 223494 81922
rect 222874 64294 222970 64350
rect 223026 64294 223094 64350
rect 223150 64294 223218 64350
rect 223274 64294 223342 64350
rect 223398 64294 223494 64350
rect 222874 64226 223494 64294
rect 222874 64170 222970 64226
rect 223026 64170 223094 64226
rect 223150 64170 223218 64226
rect 223274 64170 223342 64226
rect 223398 64170 223494 64226
rect 222874 64102 223494 64170
rect 222874 64046 222970 64102
rect 223026 64046 223094 64102
rect 223150 64046 223218 64102
rect 223274 64046 223342 64102
rect 223398 64046 223494 64102
rect 222874 63978 223494 64046
rect 222874 63922 222970 63978
rect 223026 63922 223094 63978
rect 223150 63922 223218 63978
rect 223274 63922 223342 63978
rect 223398 63922 223494 63978
rect 222874 46350 223494 63922
rect 222874 46294 222970 46350
rect 223026 46294 223094 46350
rect 223150 46294 223218 46350
rect 223274 46294 223342 46350
rect 223398 46294 223494 46350
rect 222874 46226 223494 46294
rect 222874 46170 222970 46226
rect 223026 46170 223094 46226
rect 223150 46170 223218 46226
rect 223274 46170 223342 46226
rect 223398 46170 223494 46226
rect 222874 46102 223494 46170
rect 222874 46046 222970 46102
rect 223026 46046 223094 46102
rect 223150 46046 223218 46102
rect 223274 46046 223342 46102
rect 223398 46046 223494 46102
rect 222874 45978 223494 46046
rect 222874 45922 222970 45978
rect 223026 45922 223094 45978
rect 223150 45922 223218 45978
rect 223274 45922 223342 45978
rect 223398 45922 223494 45978
rect 222874 28350 223494 45922
rect 222874 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 223494 28350
rect 222874 28226 223494 28294
rect 222874 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 223494 28226
rect 222874 28102 223494 28170
rect 222874 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 223494 28102
rect 222874 27978 223494 28046
rect 222874 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 223494 27978
rect 222874 10350 223494 27922
rect 222874 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 223494 10350
rect 222874 10226 223494 10294
rect 222874 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 223494 10226
rect 222874 10102 223494 10170
rect 222874 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 223494 10102
rect 222874 9978 223494 10046
rect 222874 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 223494 9978
rect 222874 -1120 223494 9922
rect 222874 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 223494 -1120
rect 222874 -1244 223494 -1176
rect 222874 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 223494 -1244
rect 222874 -1368 223494 -1300
rect 222874 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 223494 -1368
rect 222874 -1492 223494 -1424
rect 222874 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 223494 -1492
rect 222874 -1644 223494 -1548
rect 237154 202350 237774 210842
rect 237154 202294 237250 202350
rect 237306 202294 237374 202350
rect 237430 202294 237498 202350
rect 237554 202294 237622 202350
rect 237678 202294 237774 202350
rect 237154 202226 237774 202294
rect 237154 202170 237250 202226
rect 237306 202170 237374 202226
rect 237430 202170 237498 202226
rect 237554 202170 237622 202226
rect 237678 202170 237774 202226
rect 237154 202102 237774 202170
rect 237154 202046 237250 202102
rect 237306 202046 237374 202102
rect 237430 202046 237498 202102
rect 237554 202046 237622 202102
rect 237678 202046 237774 202102
rect 237154 201978 237774 202046
rect 237154 201922 237250 201978
rect 237306 201922 237374 201978
rect 237430 201922 237498 201978
rect 237554 201922 237622 201978
rect 237678 201922 237774 201978
rect 237154 184350 237774 201922
rect 237154 184294 237250 184350
rect 237306 184294 237374 184350
rect 237430 184294 237498 184350
rect 237554 184294 237622 184350
rect 237678 184294 237774 184350
rect 237154 184226 237774 184294
rect 237154 184170 237250 184226
rect 237306 184170 237374 184226
rect 237430 184170 237498 184226
rect 237554 184170 237622 184226
rect 237678 184170 237774 184226
rect 237154 184102 237774 184170
rect 237154 184046 237250 184102
rect 237306 184046 237374 184102
rect 237430 184046 237498 184102
rect 237554 184046 237622 184102
rect 237678 184046 237774 184102
rect 237154 183978 237774 184046
rect 237154 183922 237250 183978
rect 237306 183922 237374 183978
rect 237430 183922 237498 183978
rect 237554 183922 237622 183978
rect 237678 183922 237774 183978
rect 237154 166350 237774 183922
rect 237154 166294 237250 166350
rect 237306 166294 237374 166350
rect 237430 166294 237498 166350
rect 237554 166294 237622 166350
rect 237678 166294 237774 166350
rect 237154 166226 237774 166294
rect 237154 166170 237250 166226
rect 237306 166170 237374 166226
rect 237430 166170 237498 166226
rect 237554 166170 237622 166226
rect 237678 166170 237774 166226
rect 237154 166102 237774 166170
rect 237154 166046 237250 166102
rect 237306 166046 237374 166102
rect 237430 166046 237498 166102
rect 237554 166046 237622 166102
rect 237678 166046 237774 166102
rect 237154 165978 237774 166046
rect 237154 165922 237250 165978
rect 237306 165922 237374 165978
rect 237430 165922 237498 165978
rect 237554 165922 237622 165978
rect 237678 165922 237774 165978
rect 237154 148350 237774 165922
rect 237154 148294 237250 148350
rect 237306 148294 237374 148350
rect 237430 148294 237498 148350
rect 237554 148294 237622 148350
rect 237678 148294 237774 148350
rect 237154 148226 237774 148294
rect 237154 148170 237250 148226
rect 237306 148170 237374 148226
rect 237430 148170 237498 148226
rect 237554 148170 237622 148226
rect 237678 148170 237774 148226
rect 237154 148102 237774 148170
rect 237154 148046 237250 148102
rect 237306 148046 237374 148102
rect 237430 148046 237498 148102
rect 237554 148046 237622 148102
rect 237678 148046 237774 148102
rect 237154 147978 237774 148046
rect 237154 147922 237250 147978
rect 237306 147922 237374 147978
rect 237430 147922 237498 147978
rect 237554 147922 237622 147978
rect 237678 147922 237774 147978
rect 237154 130350 237774 147922
rect 237154 130294 237250 130350
rect 237306 130294 237374 130350
rect 237430 130294 237498 130350
rect 237554 130294 237622 130350
rect 237678 130294 237774 130350
rect 237154 130226 237774 130294
rect 237154 130170 237250 130226
rect 237306 130170 237374 130226
rect 237430 130170 237498 130226
rect 237554 130170 237622 130226
rect 237678 130170 237774 130226
rect 237154 130102 237774 130170
rect 237154 130046 237250 130102
rect 237306 130046 237374 130102
rect 237430 130046 237498 130102
rect 237554 130046 237622 130102
rect 237678 130046 237774 130102
rect 237154 129978 237774 130046
rect 237154 129922 237250 129978
rect 237306 129922 237374 129978
rect 237430 129922 237498 129978
rect 237554 129922 237622 129978
rect 237678 129922 237774 129978
rect 237154 112350 237774 129922
rect 237154 112294 237250 112350
rect 237306 112294 237374 112350
rect 237430 112294 237498 112350
rect 237554 112294 237622 112350
rect 237678 112294 237774 112350
rect 237154 112226 237774 112294
rect 237154 112170 237250 112226
rect 237306 112170 237374 112226
rect 237430 112170 237498 112226
rect 237554 112170 237622 112226
rect 237678 112170 237774 112226
rect 237154 112102 237774 112170
rect 237154 112046 237250 112102
rect 237306 112046 237374 112102
rect 237430 112046 237498 112102
rect 237554 112046 237622 112102
rect 237678 112046 237774 112102
rect 237154 111978 237774 112046
rect 237154 111922 237250 111978
rect 237306 111922 237374 111978
rect 237430 111922 237498 111978
rect 237554 111922 237622 111978
rect 237678 111922 237774 111978
rect 237154 94350 237774 111922
rect 237154 94294 237250 94350
rect 237306 94294 237374 94350
rect 237430 94294 237498 94350
rect 237554 94294 237622 94350
rect 237678 94294 237774 94350
rect 237154 94226 237774 94294
rect 237154 94170 237250 94226
rect 237306 94170 237374 94226
rect 237430 94170 237498 94226
rect 237554 94170 237622 94226
rect 237678 94170 237774 94226
rect 237154 94102 237774 94170
rect 237154 94046 237250 94102
rect 237306 94046 237374 94102
rect 237430 94046 237498 94102
rect 237554 94046 237622 94102
rect 237678 94046 237774 94102
rect 237154 93978 237774 94046
rect 237154 93922 237250 93978
rect 237306 93922 237374 93978
rect 237430 93922 237498 93978
rect 237554 93922 237622 93978
rect 237678 93922 237774 93978
rect 237154 76350 237774 93922
rect 237154 76294 237250 76350
rect 237306 76294 237374 76350
rect 237430 76294 237498 76350
rect 237554 76294 237622 76350
rect 237678 76294 237774 76350
rect 237154 76226 237774 76294
rect 237154 76170 237250 76226
rect 237306 76170 237374 76226
rect 237430 76170 237498 76226
rect 237554 76170 237622 76226
rect 237678 76170 237774 76226
rect 237154 76102 237774 76170
rect 237154 76046 237250 76102
rect 237306 76046 237374 76102
rect 237430 76046 237498 76102
rect 237554 76046 237622 76102
rect 237678 76046 237774 76102
rect 237154 75978 237774 76046
rect 237154 75922 237250 75978
rect 237306 75922 237374 75978
rect 237430 75922 237498 75978
rect 237554 75922 237622 75978
rect 237678 75922 237774 75978
rect 237154 58350 237774 75922
rect 237154 58294 237250 58350
rect 237306 58294 237374 58350
rect 237430 58294 237498 58350
rect 237554 58294 237622 58350
rect 237678 58294 237774 58350
rect 237154 58226 237774 58294
rect 237154 58170 237250 58226
rect 237306 58170 237374 58226
rect 237430 58170 237498 58226
rect 237554 58170 237622 58226
rect 237678 58170 237774 58226
rect 237154 58102 237774 58170
rect 237154 58046 237250 58102
rect 237306 58046 237374 58102
rect 237430 58046 237498 58102
rect 237554 58046 237622 58102
rect 237678 58046 237774 58102
rect 237154 57978 237774 58046
rect 237154 57922 237250 57978
rect 237306 57922 237374 57978
rect 237430 57922 237498 57978
rect 237554 57922 237622 57978
rect 237678 57922 237774 57978
rect 237154 40350 237774 57922
rect 237154 40294 237250 40350
rect 237306 40294 237374 40350
rect 237430 40294 237498 40350
rect 237554 40294 237622 40350
rect 237678 40294 237774 40350
rect 237154 40226 237774 40294
rect 237154 40170 237250 40226
rect 237306 40170 237374 40226
rect 237430 40170 237498 40226
rect 237554 40170 237622 40226
rect 237678 40170 237774 40226
rect 237154 40102 237774 40170
rect 237154 40046 237250 40102
rect 237306 40046 237374 40102
rect 237430 40046 237498 40102
rect 237554 40046 237622 40102
rect 237678 40046 237774 40102
rect 237154 39978 237774 40046
rect 237154 39922 237250 39978
rect 237306 39922 237374 39978
rect 237430 39922 237498 39978
rect 237554 39922 237622 39978
rect 237678 39922 237774 39978
rect 237154 22350 237774 39922
rect 237154 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 237774 22350
rect 237154 22226 237774 22294
rect 237154 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 237774 22226
rect 237154 22102 237774 22170
rect 237154 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 237774 22102
rect 237154 21978 237774 22046
rect 237154 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 237774 21978
rect 237154 4350 237774 21922
rect 237154 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 237774 4350
rect 237154 4226 237774 4294
rect 237154 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 237774 4226
rect 237154 4102 237774 4170
rect 237154 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 237774 4102
rect 237154 3978 237774 4046
rect 237154 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 237774 3978
rect 237154 -160 237774 3922
rect 237154 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 237774 -160
rect 237154 -284 237774 -216
rect 237154 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 237774 -284
rect 237154 -408 237774 -340
rect 237154 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 237774 -408
rect 237154 -532 237774 -464
rect 237154 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 237774 -532
rect 237154 -1644 237774 -588
rect 240874 208350 241494 210842
rect 240874 208294 240970 208350
rect 241026 208294 241094 208350
rect 241150 208294 241218 208350
rect 241274 208294 241342 208350
rect 241398 208294 241494 208350
rect 240874 208226 241494 208294
rect 240874 208170 240970 208226
rect 241026 208170 241094 208226
rect 241150 208170 241218 208226
rect 241274 208170 241342 208226
rect 241398 208170 241494 208226
rect 240874 208102 241494 208170
rect 240874 208046 240970 208102
rect 241026 208046 241094 208102
rect 241150 208046 241218 208102
rect 241274 208046 241342 208102
rect 241398 208046 241494 208102
rect 240874 207978 241494 208046
rect 240874 207922 240970 207978
rect 241026 207922 241094 207978
rect 241150 207922 241218 207978
rect 241274 207922 241342 207978
rect 241398 207922 241494 207978
rect 240874 190350 241494 207922
rect 250528 208350 250848 208384
rect 250528 208294 250598 208350
rect 250654 208294 250722 208350
rect 250778 208294 250848 208350
rect 250528 208226 250848 208294
rect 250528 208170 250598 208226
rect 250654 208170 250722 208226
rect 250778 208170 250848 208226
rect 250528 208102 250848 208170
rect 250528 208046 250598 208102
rect 250654 208046 250722 208102
rect 250778 208046 250848 208102
rect 250528 207978 250848 208046
rect 250528 207922 250598 207978
rect 250654 207922 250722 207978
rect 250778 207922 250848 207978
rect 250528 207888 250848 207922
rect 240874 190294 240970 190350
rect 241026 190294 241094 190350
rect 241150 190294 241218 190350
rect 241274 190294 241342 190350
rect 241398 190294 241494 190350
rect 240874 190226 241494 190294
rect 240874 190170 240970 190226
rect 241026 190170 241094 190226
rect 241150 190170 241218 190226
rect 241274 190170 241342 190226
rect 241398 190170 241494 190226
rect 240874 190102 241494 190170
rect 240874 190046 240970 190102
rect 241026 190046 241094 190102
rect 241150 190046 241218 190102
rect 241274 190046 241342 190102
rect 241398 190046 241494 190102
rect 240874 189978 241494 190046
rect 240874 189922 240970 189978
rect 241026 189922 241094 189978
rect 241150 189922 241218 189978
rect 241274 189922 241342 189978
rect 241398 189922 241494 189978
rect 240874 172350 241494 189922
rect 240874 172294 240970 172350
rect 241026 172294 241094 172350
rect 241150 172294 241218 172350
rect 241274 172294 241342 172350
rect 241398 172294 241494 172350
rect 240874 172226 241494 172294
rect 240874 172170 240970 172226
rect 241026 172170 241094 172226
rect 241150 172170 241218 172226
rect 241274 172170 241342 172226
rect 241398 172170 241494 172226
rect 240874 172102 241494 172170
rect 240874 172046 240970 172102
rect 241026 172046 241094 172102
rect 241150 172046 241218 172102
rect 241274 172046 241342 172102
rect 241398 172046 241494 172102
rect 240874 171978 241494 172046
rect 240874 171922 240970 171978
rect 241026 171922 241094 171978
rect 241150 171922 241218 171978
rect 241274 171922 241342 171978
rect 241398 171922 241494 171978
rect 240874 154350 241494 171922
rect 240874 154294 240970 154350
rect 241026 154294 241094 154350
rect 241150 154294 241218 154350
rect 241274 154294 241342 154350
rect 241398 154294 241494 154350
rect 240874 154226 241494 154294
rect 240874 154170 240970 154226
rect 241026 154170 241094 154226
rect 241150 154170 241218 154226
rect 241274 154170 241342 154226
rect 241398 154170 241494 154226
rect 240874 154102 241494 154170
rect 240874 154046 240970 154102
rect 241026 154046 241094 154102
rect 241150 154046 241218 154102
rect 241274 154046 241342 154102
rect 241398 154046 241494 154102
rect 240874 153978 241494 154046
rect 240874 153922 240970 153978
rect 241026 153922 241094 153978
rect 241150 153922 241218 153978
rect 241274 153922 241342 153978
rect 241398 153922 241494 153978
rect 240874 136350 241494 153922
rect 240874 136294 240970 136350
rect 241026 136294 241094 136350
rect 241150 136294 241218 136350
rect 241274 136294 241342 136350
rect 241398 136294 241494 136350
rect 240874 136226 241494 136294
rect 240874 136170 240970 136226
rect 241026 136170 241094 136226
rect 241150 136170 241218 136226
rect 241274 136170 241342 136226
rect 241398 136170 241494 136226
rect 240874 136102 241494 136170
rect 240874 136046 240970 136102
rect 241026 136046 241094 136102
rect 241150 136046 241218 136102
rect 241274 136046 241342 136102
rect 241398 136046 241494 136102
rect 240874 135978 241494 136046
rect 240874 135922 240970 135978
rect 241026 135922 241094 135978
rect 241150 135922 241218 135978
rect 241274 135922 241342 135978
rect 241398 135922 241494 135978
rect 240874 118350 241494 135922
rect 240874 118294 240970 118350
rect 241026 118294 241094 118350
rect 241150 118294 241218 118350
rect 241274 118294 241342 118350
rect 241398 118294 241494 118350
rect 240874 118226 241494 118294
rect 240874 118170 240970 118226
rect 241026 118170 241094 118226
rect 241150 118170 241218 118226
rect 241274 118170 241342 118226
rect 241398 118170 241494 118226
rect 240874 118102 241494 118170
rect 240874 118046 240970 118102
rect 241026 118046 241094 118102
rect 241150 118046 241218 118102
rect 241274 118046 241342 118102
rect 241398 118046 241494 118102
rect 240874 117978 241494 118046
rect 240874 117922 240970 117978
rect 241026 117922 241094 117978
rect 241150 117922 241218 117978
rect 241274 117922 241342 117978
rect 241398 117922 241494 117978
rect 240874 100350 241494 117922
rect 240874 100294 240970 100350
rect 241026 100294 241094 100350
rect 241150 100294 241218 100350
rect 241274 100294 241342 100350
rect 241398 100294 241494 100350
rect 240874 100226 241494 100294
rect 240874 100170 240970 100226
rect 241026 100170 241094 100226
rect 241150 100170 241218 100226
rect 241274 100170 241342 100226
rect 241398 100170 241494 100226
rect 240874 100102 241494 100170
rect 240874 100046 240970 100102
rect 241026 100046 241094 100102
rect 241150 100046 241218 100102
rect 241274 100046 241342 100102
rect 241398 100046 241494 100102
rect 240874 99978 241494 100046
rect 240874 99922 240970 99978
rect 241026 99922 241094 99978
rect 241150 99922 241218 99978
rect 241274 99922 241342 99978
rect 241398 99922 241494 99978
rect 240874 82350 241494 99922
rect 240874 82294 240970 82350
rect 241026 82294 241094 82350
rect 241150 82294 241218 82350
rect 241274 82294 241342 82350
rect 241398 82294 241494 82350
rect 240874 82226 241494 82294
rect 240874 82170 240970 82226
rect 241026 82170 241094 82226
rect 241150 82170 241218 82226
rect 241274 82170 241342 82226
rect 241398 82170 241494 82226
rect 240874 82102 241494 82170
rect 240874 82046 240970 82102
rect 241026 82046 241094 82102
rect 241150 82046 241218 82102
rect 241274 82046 241342 82102
rect 241398 82046 241494 82102
rect 240874 81978 241494 82046
rect 240874 81922 240970 81978
rect 241026 81922 241094 81978
rect 241150 81922 241218 81978
rect 241274 81922 241342 81978
rect 241398 81922 241494 81978
rect 240874 64350 241494 81922
rect 240874 64294 240970 64350
rect 241026 64294 241094 64350
rect 241150 64294 241218 64350
rect 241274 64294 241342 64350
rect 241398 64294 241494 64350
rect 240874 64226 241494 64294
rect 240874 64170 240970 64226
rect 241026 64170 241094 64226
rect 241150 64170 241218 64226
rect 241274 64170 241342 64226
rect 241398 64170 241494 64226
rect 240874 64102 241494 64170
rect 240874 64046 240970 64102
rect 241026 64046 241094 64102
rect 241150 64046 241218 64102
rect 241274 64046 241342 64102
rect 241398 64046 241494 64102
rect 240874 63978 241494 64046
rect 240874 63922 240970 63978
rect 241026 63922 241094 63978
rect 241150 63922 241218 63978
rect 241274 63922 241342 63978
rect 241398 63922 241494 63978
rect 240874 46350 241494 63922
rect 240874 46294 240970 46350
rect 241026 46294 241094 46350
rect 241150 46294 241218 46350
rect 241274 46294 241342 46350
rect 241398 46294 241494 46350
rect 240874 46226 241494 46294
rect 240874 46170 240970 46226
rect 241026 46170 241094 46226
rect 241150 46170 241218 46226
rect 241274 46170 241342 46226
rect 241398 46170 241494 46226
rect 240874 46102 241494 46170
rect 240874 46046 240970 46102
rect 241026 46046 241094 46102
rect 241150 46046 241218 46102
rect 241274 46046 241342 46102
rect 241398 46046 241494 46102
rect 240874 45978 241494 46046
rect 240874 45922 240970 45978
rect 241026 45922 241094 45978
rect 241150 45922 241218 45978
rect 241274 45922 241342 45978
rect 241398 45922 241494 45978
rect 240874 28350 241494 45922
rect 240874 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 241494 28350
rect 240874 28226 241494 28294
rect 240874 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 241494 28226
rect 240874 28102 241494 28170
rect 240874 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 241494 28102
rect 240874 27978 241494 28046
rect 240874 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 241494 27978
rect 240874 10350 241494 27922
rect 240874 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 241494 10350
rect 240874 10226 241494 10294
rect 240874 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 241494 10226
rect 240874 10102 241494 10170
rect 240874 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 241494 10102
rect 240874 9978 241494 10046
rect 240874 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 241494 9978
rect 240874 -1120 241494 9922
rect 240874 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 241494 -1120
rect 240874 -1244 241494 -1176
rect 240874 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 241494 -1244
rect 240874 -1368 241494 -1300
rect 240874 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 241494 -1368
rect 240874 -1492 241494 -1424
rect 240874 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 241494 -1492
rect 240874 -1644 241494 -1548
rect 255154 202350 255774 210842
rect 255154 202294 255250 202350
rect 255306 202294 255374 202350
rect 255430 202294 255498 202350
rect 255554 202294 255622 202350
rect 255678 202294 255774 202350
rect 255154 202226 255774 202294
rect 255154 202170 255250 202226
rect 255306 202170 255374 202226
rect 255430 202170 255498 202226
rect 255554 202170 255622 202226
rect 255678 202170 255774 202226
rect 255154 202102 255774 202170
rect 255154 202046 255250 202102
rect 255306 202046 255374 202102
rect 255430 202046 255498 202102
rect 255554 202046 255622 202102
rect 255678 202046 255774 202102
rect 255154 201978 255774 202046
rect 255154 201922 255250 201978
rect 255306 201922 255374 201978
rect 255430 201922 255498 201978
rect 255554 201922 255622 201978
rect 255678 201922 255774 201978
rect 255154 184350 255774 201922
rect 255154 184294 255250 184350
rect 255306 184294 255374 184350
rect 255430 184294 255498 184350
rect 255554 184294 255622 184350
rect 255678 184294 255774 184350
rect 255154 184226 255774 184294
rect 255154 184170 255250 184226
rect 255306 184170 255374 184226
rect 255430 184170 255498 184226
rect 255554 184170 255622 184226
rect 255678 184170 255774 184226
rect 255154 184102 255774 184170
rect 255154 184046 255250 184102
rect 255306 184046 255374 184102
rect 255430 184046 255498 184102
rect 255554 184046 255622 184102
rect 255678 184046 255774 184102
rect 255154 183978 255774 184046
rect 255154 183922 255250 183978
rect 255306 183922 255374 183978
rect 255430 183922 255498 183978
rect 255554 183922 255622 183978
rect 255678 183922 255774 183978
rect 255154 166350 255774 183922
rect 255154 166294 255250 166350
rect 255306 166294 255374 166350
rect 255430 166294 255498 166350
rect 255554 166294 255622 166350
rect 255678 166294 255774 166350
rect 255154 166226 255774 166294
rect 255154 166170 255250 166226
rect 255306 166170 255374 166226
rect 255430 166170 255498 166226
rect 255554 166170 255622 166226
rect 255678 166170 255774 166226
rect 255154 166102 255774 166170
rect 255154 166046 255250 166102
rect 255306 166046 255374 166102
rect 255430 166046 255498 166102
rect 255554 166046 255622 166102
rect 255678 166046 255774 166102
rect 255154 165978 255774 166046
rect 255154 165922 255250 165978
rect 255306 165922 255374 165978
rect 255430 165922 255498 165978
rect 255554 165922 255622 165978
rect 255678 165922 255774 165978
rect 255154 148350 255774 165922
rect 255154 148294 255250 148350
rect 255306 148294 255374 148350
rect 255430 148294 255498 148350
rect 255554 148294 255622 148350
rect 255678 148294 255774 148350
rect 255154 148226 255774 148294
rect 255154 148170 255250 148226
rect 255306 148170 255374 148226
rect 255430 148170 255498 148226
rect 255554 148170 255622 148226
rect 255678 148170 255774 148226
rect 255154 148102 255774 148170
rect 255154 148046 255250 148102
rect 255306 148046 255374 148102
rect 255430 148046 255498 148102
rect 255554 148046 255622 148102
rect 255678 148046 255774 148102
rect 255154 147978 255774 148046
rect 255154 147922 255250 147978
rect 255306 147922 255374 147978
rect 255430 147922 255498 147978
rect 255554 147922 255622 147978
rect 255678 147922 255774 147978
rect 255154 130350 255774 147922
rect 255154 130294 255250 130350
rect 255306 130294 255374 130350
rect 255430 130294 255498 130350
rect 255554 130294 255622 130350
rect 255678 130294 255774 130350
rect 255154 130226 255774 130294
rect 255154 130170 255250 130226
rect 255306 130170 255374 130226
rect 255430 130170 255498 130226
rect 255554 130170 255622 130226
rect 255678 130170 255774 130226
rect 255154 130102 255774 130170
rect 255154 130046 255250 130102
rect 255306 130046 255374 130102
rect 255430 130046 255498 130102
rect 255554 130046 255622 130102
rect 255678 130046 255774 130102
rect 255154 129978 255774 130046
rect 255154 129922 255250 129978
rect 255306 129922 255374 129978
rect 255430 129922 255498 129978
rect 255554 129922 255622 129978
rect 255678 129922 255774 129978
rect 255154 112350 255774 129922
rect 255154 112294 255250 112350
rect 255306 112294 255374 112350
rect 255430 112294 255498 112350
rect 255554 112294 255622 112350
rect 255678 112294 255774 112350
rect 255154 112226 255774 112294
rect 255154 112170 255250 112226
rect 255306 112170 255374 112226
rect 255430 112170 255498 112226
rect 255554 112170 255622 112226
rect 255678 112170 255774 112226
rect 255154 112102 255774 112170
rect 255154 112046 255250 112102
rect 255306 112046 255374 112102
rect 255430 112046 255498 112102
rect 255554 112046 255622 112102
rect 255678 112046 255774 112102
rect 255154 111978 255774 112046
rect 255154 111922 255250 111978
rect 255306 111922 255374 111978
rect 255430 111922 255498 111978
rect 255554 111922 255622 111978
rect 255678 111922 255774 111978
rect 255154 94350 255774 111922
rect 255154 94294 255250 94350
rect 255306 94294 255374 94350
rect 255430 94294 255498 94350
rect 255554 94294 255622 94350
rect 255678 94294 255774 94350
rect 255154 94226 255774 94294
rect 255154 94170 255250 94226
rect 255306 94170 255374 94226
rect 255430 94170 255498 94226
rect 255554 94170 255622 94226
rect 255678 94170 255774 94226
rect 255154 94102 255774 94170
rect 255154 94046 255250 94102
rect 255306 94046 255374 94102
rect 255430 94046 255498 94102
rect 255554 94046 255622 94102
rect 255678 94046 255774 94102
rect 255154 93978 255774 94046
rect 255154 93922 255250 93978
rect 255306 93922 255374 93978
rect 255430 93922 255498 93978
rect 255554 93922 255622 93978
rect 255678 93922 255774 93978
rect 255154 76350 255774 93922
rect 255154 76294 255250 76350
rect 255306 76294 255374 76350
rect 255430 76294 255498 76350
rect 255554 76294 255622 76350
rect 255678 76294 255774 76350
rect 255154 76226 255774 76294
rect 255154 76170 255250 76226
rect 255306 76170 255374 76226
rect 255430 76170 255498 76226
rect 255554 76170 255622 76226
rect 255678 76170 255774 76226
rect 255154 76102 255774 76170
rect 255154 76046 255250 76102
rect 255306 76046 255374 76102
rect 255430 76046 255498 76102
rect 255554 76046 255622 76102
rect 255678 76046 255774 76102
rect 255154 75978 255774 76046
rect 255154 75922 255250 75978
rect 255306 75922 255374 75978
rect 255430 75922 255498 75978
rect 255554 75922 255622 75978
rect 255678 75922 255774 75978
rect 255154 58350 255774 75922
rect 255154 58294 255250 58350
rect 255306 58294 255374 58350
rect 255430 58294 255498 58350
rect 255554 58294 255622 58350
rect 255678 58294 255774 58350
rect 255154 58226 255774 58294
rect 255154 58170 255250 58226
rect 255306 58170 255374 58226
rect 255430 58170 255498 58226
rect 255554 58170 255622 58226
rect 255678 58170 255774 58226
rect 255154 58102 255774 58170
rect 255154 58046 255250 58102
rect 255306 58046 255374 58102
rect 255430 58046 255498 58102
rect 255554 58046 255622 58102
rect 255678 58046 255774 58102
rect 255154 57978 255774 58046
rect 255154 57922 255250 57978
rect 255306 57922 255374 57978
rect 255430 57922 255498 57978
rect 255554 57922 255622 57978
rect 255678 57922 255774 57978
rect 255154 40350 255774 57922
rect 255154 40294 255250 40350
rect 255306 40294 255374 40350
rect 255430 40294 255498 40350
rect 255554 40294 255622 40350
rect 255678 40294 255774 40350
rect 255154 40226 255774 40294
rect 255154 40170 255250 40226
rect 255306 40170 255374 40226
rect 255430 40170 255498 40226
rect 255554 40170 255622 40226
rect 255678 40170 255774 40226
rect 255154 40102 255774 40170
rect 255154 40046 255250 40102
rect 255306 40046 255374 40102
rect 255430 40046 255498 40102
rect 255554 40046 255622 40102
rect 255678 40046 255774 40102
rect 255154 39978 255774 40046
rect 255154 39922 255250 39978
rect 255306 39922 255374 39978
rect 255430 39922 255498 39978
rect 255554 39922 255622 39978
rect 255678 39922 255774 39978
rect 255154 22350 255774 39922
rect 255154 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 255774 22350
rect 255154 22226 255774 22294
rect 255154 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 255774 22226
rect 255154 22102 255774 22170
rect 255154 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 255774 22102
rect 255154 21978 255774 22046
rect 255154 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 255774 21978
rect 255154 4350 255774 21922
rect 255154 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 255774 4350
rect 255154 4226 255774 4294
rect 255154 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 255774 4226
rect 255154 4102 255774 4170
rect 255154 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 255774 4102
rect 255154 3978 255774 4046
rect 255154 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 255774 3978
rect 255154 -160 255774 3922
rect 255154 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 255774 -160
rect 255154 -284 255774 -216
rect 255154 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 255774 -284
rect 255154 -408 255774 -340
rect 255154 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 255774 -408
rect 255154 -532 255774 -464
rect 255154 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 255774 -532
rect 255154 -1644 255774 -588
rect 258874 208350 259494 210842
rect 258874 208294 258970 208350
rect 259026 208294 259094 208350
rect 259150 208294 259218 208350
rect 259274 208294 259342 208350
rect 259398 208294 259494 208350
rect 258874 208226 259494 208294
rect 258874 208170 258970 208226
rect 259026 208170 259094 208226
rect 259150 208170 259218 208226
rect 259274 208170 259342 208226
rect 259398 208170 259494 208226
rect 258874 208102 259494 208170
rect 258874 208046 258970 208102
rect 259026 208046 259094 208102
rect 259150 208046 259218 208102
rect 259274 208046 259342 208102
rect 259398 208046 259494 208102
rect 258874 207978 259494 208046
rect 258874 207922 258970 207978
rect 259026 207922 259094 207978
rect 259150 207922 259218 207978
rect 259274 207922 259342 207978
rect 259398 207922 259494 207978
rect 258874 190350 259494 207922
rect 258874 190294 258970 190350
rect 259026 190294 259094 190350
rect 259150 190294 259218 190350
rect 259274 190294 259342 190350
rect 259398 190294 259494 190350
rect 258874 190226 259494 190294
rect 258874 190170 258970 190226
rect 259026 190170 259094 190226
rect 259150 190170 259218 190226
rect 259274 190170 259342 190226
rect 259398 190170 259494 190226
rect 258874 190102 259494 190170
rect 258874 190046 258970 190102
rect 259026 190046 259094 190102
rect 259150 190046 259218 190102
rect 259274 190046 259342 190102
rect 259398 190046 259494 190102
rect 258874 189978 259494 190046
rect 258874 189922 258970 189978
rect 259026 189922 259094 189978
rect 259150 189922 259218 189978
rect 259274 189922 259342 189978
rect 259398 189922 259494 189978
rect 258874 172350 259494 189922
rect 258874 172294 258970 172350
rect 259026 172294 259094 172350
rect 259150 172294 259218 172350
rect 259274 172294 259342 172350
rect 259398 172294 259494 172350
rect 258874 172226 259494 172294
rect 258874 172170 258970 172226
rect 259026 172170 259094 172226
rect 259150 172170 259218 172226
rect 259274 172170 259342 172226
rect 259398 172170 259494 172226
rect 258874 172102 259494 172170
rect 258874 172046 258970 172102
rect 259026 172046 259094 172102
rect 259150 172046 259218 172102
rect 259274 172046 259342 172102
rect 259398 172046 259494 172102
rect 258874 171978 259494 172046
rect 258874 171922 258970 171978
rect 259026 171922 259094 171978
rect 259150 171922 259218 171978
rect 259274 171922 259342 171978
rect 259398 171922 259494 171978
rect 258874 154350 259494 171922
rect 258874 154294 258970 154350
rect 259026 154294 259094 154350
rect 259150 154294 259218 154350
rect 259274 154294 259342 154350
rect 259398 154294 259494 154350
rect 258874 154226 259494 154294
rect 258874 154170 258970 154226
rect 259026 154170 259094 154226
rect 259150 154170 259218 154226
rect 259274 154170 259342 154226
rect 259398 154170 259494 154226
rect 258874 154102 259494 154170
rect 258874 154046 258970 154102
rect 259026 154046 259094 154102
rect 259150 154046 259218 154102
rect 259274 154046 259342 154102
rect 259398 154046 259494 154102
rect 258874 153978 259494 154046
rect 258874 153922 258970 153978
rect 259026 153922 259094 153978
rect 259150 153922 259218 153978
rect 259274 153922 259342 153978
rect 259398 153922 259494 153978
rect 258874 136350 259494 153922
rect 258874 136294 258970 136350
rect 259026 136294 259094 136350
rect 259150 136294 259218 136350
rect 259274 136294 259342 136350
rect 259398 136294 259494 136350
rect 258874 136226 259494 136294
rect 258874 136170 258970 136226
rect 259026 136170 259094 136226
rect 259150 136170 259218 136226
rect 259274 136170 259342 136226
rect 259398 136170 259494 136226
rect 258874 136102 259494 136170
rect 258874 136046 258970 136102
rect 259026 136046 259094 136102
rect 259150 136046 259218 136102
rect 259274 136046 259342 136102
rect 259398 136046 259494 136102
rect 258874 135978 259494 136046
rect 258874 135922 258970 135978
rect 259026 135922 259094 135978
rect 259150 135922 259218 135978
rect 259274 135922 259342 135978
rect 259398 135922 259494 135978
rect 258874 118350 259494 135922
rect 258874 118294 258970 118350
rect 259026 118294 259094 118350
rect 259150 118294 259218 118350
rect 259274 118294 259342 118350
rect 259398 118294 259494 118350
rect 258874 118226 259494 118294
rect 258874 118170 258970 118226
rect 259026 118170 259094 118226
rect 259150 118170 259218 118226
rect 259274 118170 259342 118226
rect 259398 118170 259494 118226
rect 258874 118102 259494 118170
rect 258874 118046 258970 118102
rect 259026 118046 259094 118102
rect 259150 118046 259218 118102
rect 259274 118046 259342 118102
rect 259398 118046 259494 118102
rect 258874 117978 259494 118046
rect 258874 117922 258970 117978
rect 259026 117922 259094 117978
rect 259150 117922 259218 117978
rect 259274 117922 259342 117978
rect 259398 117922 259494 117978
rect 258874 100350 259494 117922
rect 258874 100294 258970 100350
rect 259026 100294 259094 100350
rect 259150 100294 259218 100350
rect 259274 100294 259342 100350
rect 259398 100294 259494 100350
rect 258874 100226 259494 100294
rect 258874 100170 258970 100226
rect 259026 100170 259094 100226
rect 259150 100170 259218 100226
rect 259274 100170 259342 100226
rect 259398 100170 259494 100226
rect 258874 100102 259494 100170
rect 258874 100046 258970 100102
rect 259026 100046 259094 100102
rect 259150 100046 259218 100102
rect 259274 100046 259342 100102
rect 259398 100046 259494 100102
rect 258874 99978 259494 100046
rect 258874 99922 258970 99978
rect 259026 99922 259094 99978
rect 259150 99922 259218 99978
rect 259274 99922 259342 99978
rect 259398 99922 259494 99978
rect 258874 82350 259494 99922
rect 258874 82294 258970 82350
rect 259026 82294 259094 82350
rect 259150 82294 259218 82350
rect 259274 82294 259342 82350
rect 259398 82294 259494 82350
rect 258874 82226 259494 82294
rect 258874 82170 258970 82226
rect 259026 82170 259094 82226
rect 259150 82170 259218 82226
rect 259274 82170 259342 82226
rect 259398 82170 259494 82226
rect 258874 82102 259494 82170
rect 258874 82046 258970 82102
rect 259026 82046 259094 82102
rect 259150 82046 259218 82102
rect 259274 82046 259342 82102
rect 259398 82046 259494 82102
rect 258874 81978 259494 82046
rect 258874 81922 258970 81978
rect 259026 81922 259094 81978
rect 259150 81922 259218 81978
rect 259274 81922 259342 81978
rect 259398 81922 259494 81978
rect 258874 64350 259494 81922
rect 258874 64294 258970 64350
rect 259026 64294 259094 64350
rect 259150 64294 259218 64350
rect 259274 64294 259342 64350
rect 259398 64294 259494 64350
rect 258874 64226 259494 64294
rect 258874 64170 258970 64226
rect 259026 64170 259094 64226
rect 259150 64170 259218 64226
rect 259274 64170 259342 64226
rect 259398 64170 259494 64226
rect 258874 64102 259494 64170
rect 258874 64046 258970 64102
rect 259026 64046 259094 64102
rect 259150 64046 259218 64102
rect 259274 64046 259342 64102
rect 259398 64046 259494 64102
rect 258874 63978 259494 64046
rect 258874 63922 258970 63978
rect 259026 63922 259094 63978
rect 259150 63922 259218 63978
rect 259274 63922 259342 63978
rect 259398 63922 259494 63978
rect 258874 46350 259494 63922
rect 258874 46294 258970 46350
rect 259026 46294 259094 46350
rect 259150 46294 259218 46350
rect 259274 46294 259342 46350
rect 259398 46294 259494 46350
rect 258874 46226 259494 46294
rect 258874 46170 258970 46226
rect 259026 46170 259094 46226
rect 259150 46170 259218 46226
rect 259274 46170 259342 46226
rect 259398 46170 259494 46226
rect 258874 46102 259494 46170
rect 258874 46046 258970 46102
rect 259026 46046 259094 46102
rect 259150 46046 259218 46102
rect 259274 46046 259342 46102
rect 259398 46046 259494 46102
rect 258874 45978 259494 46046
rect 258874 45922 258970 45978
rect 259026 45922 259094 45978
rect 259150 45922 259218 45978
rect 259274 45922 259342 45978
rect 259398 45922 259494 45978
rect 258874 28350 259494 45922
rect 258874 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 259494 28350
rect 258874 28226 259494 28294
rect 258874 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 259494 28226
rect 258874 28102 259494 28170
rect 258874 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 259494 28102
rect 258874 27978 259494 28046
rect 258874 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 259494 27978
rect 258874 10350 259494 27922
rect 258874 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 259494 10350
rect 258874 10226 259494 10294
rect 258874 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 259494 10226
rect 258874 10102 259494 10170
rect 258874 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 259494 10102
rect 258874 9978 259494 10046
rect 258874 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 259494 9978
rect 258874 -1120 259494 9922
rect 258874 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 259494 -1120
rect 258874 -1244 259494 -1176
rect 258874 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 259494 -1244
rect 258874 -1368 259494 -1300
rect 258874 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 259494 -1368
rect 258874 -1492 259494 -1424
rect 258874 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 259494 -1492
rect 258874 -1644 259494 -1548
rect 273154 202350 273774 210842
rect 273154 202294 273250 202350
rect 273306 202294 273374 202350
rect 273430 202294 273498 202350
rect 273554 202294 273622 202350
rect 273678 202294 273774 202350
rect 273154 202226 273774 202294
rect 273154 202170 273250 202226
rect 273306 202170 273374 202226
rect 273430 202170 273498 202226
rect 273554 202170 273622 202226
rect 273678 202170 273774 202226
rect 273154 202102 273774 202170
rect 273154 202046 273250 202102
rect 273306 202046 273374 202102
rect 273430 202046 273498 202102
rect 273554 202046 273622 202102
rect 273678 202046 273774 202102
rect 273154 201978 273774 202046
rect 273154 201922 273250 201978
rect 273306 201922 273374 201978
rect 273430 201922 273498 201978
rect 273554 201922 273622 201978
rect 273678 201922 273774 201978
rect 273154 184350 273774 201922
rect 273154 184294 273250 184350
rect 273306 184294 273374 184350
rect 273430 184294 273498 184350
rect 273554 184294 273622 184350
rect 273678 184294 273774 184350
rect 273154 184226 273774 184294
rect 273154 184170 273250 184226
rect 273306 184170 273374 184226
rect 273430 184170 273498 184226
rect 273554 184170 273622 184226
rect 273678 184170 273774 184226
rect 273154 184102 273774 184170
rect 273154 184046 273250 184102
rect 273306 184046 273374 184102
rect 273430 184046 273498 184102
rect 273554 184046 273622 184102
rect 273678 184046 273774 184102
rect 273154 183978 273774 184046
rect 273154 183922 273250 183978
rect 273306 183922 273374 183978
rect 273430 183922 273498 183978
rect 273554 183922 273622 183978
rect 273678 183922 273774 183978
rect 273154 166350 273774 183922
rect 273154 166294 273250 166350
rect 273306 166294 273374 166350
rect 273430 166294 273498 166350
rect 273554 166294 273622 166350
rect 273678 166294 273774 166350
rect 273154 166226 273774 166294
rect 273154 166170 273250 166226
rect 273306 166170 273374 166226
rect 273430 166170 273498 166226
rect 273554 166170 273622 166226
rect 273678 166170 273774 166226
rect 273154 166102 273774 166170
rect 273154 166046 273250 166102
rect 273306 166046 273374 166102
rect 273430 166046 273498 166102
rect 273554 166046 273622 166102
rect 273678 166046 273774 166102
rect 273154 165978 273774 166046
rect 273154 165922 273250 165978
rect 273306 165922 273374 165978
rect 273430 165922 273498 165978
rect 273554 165922 273622 165978
rect 273678 165922 273774 165978
rect 273154 148350 273774 165922
rect 273154 148294 273250 148350
rect 273306 148294 273374 148350
rect 273430 148294 273498 148350
rect 273554 148294 273622 148350
rect 273678 148294 273774 148350
rect 273154 148226 273774 148294
rect 273154 148170 273250 148226
rect 273306 148170 273374 148226
rect 273430 148170 273498 148226
rect 273554 148170 273622 148226
rect 273678 148170 273774 148226
rect 273154 148102 273774 148170
rect 273154 148046 273250 148102
rect 273306 148046 273374 148102
rect 273430 148046 273498 148102
rect 273554 148046 273622 148102
rect 273678 148046 273774 148102
rect 273154 147978 273774 148046
rect 273154 147922 273250 147978
rect 273306 147922 273374 147978
rect 273430 147922 273498 147978
rect 273554 147922 273622 147978
rect 273678 147922 273774 147978
rect 273154 130350 273774 147922
rect 273154 130294 273250 130350
rect 273306 130294 273374 130350
rect 273430 130294 273498 130350
rect 273554 130294 273622 130350
rect 273678 130294 273774 130350
rect 273154 130226 273774 130294
rect 273154 130170 273250 130226
rect 273306 130170 273374 130226
rect 273430 130170 273498 130226
rect 273554 130170 273622 130226
rect 273678 130170 273774 130226
rect 273154 130102 273774 130170
rect 273154 130046 273250 130102
rect 273306 130046 273374 130102
rect 273430 130046 273498 130102
rect 273554 130046 273622 130102
rect 273678 130046 273774 130102
rect 273154 129978 273774 130046
rect 273154 129922 273250 129978
rect 273306 129922 273374 129978
rect 273430 129922 273498 129978
rect 273554 129922 273622 129978
rect 273678 129922 273774 129978
rect 273154 112350 273774 129922
rect 273154 112294 273250 112350
rect 273306 112294 273374 112350
rect 273430 112294 273498 112350
rect 273554 112294 273622 112350
rect 273678 112294 273774 112350
rect 273154 112226 273774 112294
rect 273154 112170 273250 112226
rect 273306 112170 273374 112226
rect 273430 112170 273498 112226
rect 273554 112170 273622 112226
rect 273678 112170 273774 112226
rect 273154 112102 273774 112170
rect 273154 112046 273250 112102
rect 273306 112046 273374 112102
rect 273430 112046 273498 112102
rect 273554 112046 273622 112102
rect 273678 112046 273774 112102
rect 273154 111978 273774 112046
rect 273154 111922 273250 111978
rect 273306 111922 273374 111978
rect 273430 111922 273498 111978
rect 273554 111922 273622 111978
rect 273678 111922 273774 111978
rect 273154 94350 273774 111922
rect 273154 94294 273250 94350
rect 273306 94294 273374 94350
rect 273430 94294 273498 94350
rect 273554 94294 273622 94350
rect 273678 94294 273774 94350
rect 273154 94226 273774 94294
rect 273154 94170 273250 94226
rect 273306 94170 273374 94226
rect 273430 94170 273498 94226
rect 273554 94170 273622 94226
rect 273678 94170 273774 94226
rect 273154 94102 273774 94170
rect 273154 94046 273250 94102
rect 273306 94046 273374 94102
rect 273430 94046 273498 94102
rect 273554 94046 273622 94102
rect 273678 94046 273774 94102
rect 273154 93978 273774 94046
rect 273154 93922 273250 93978
rect 273306 93922 273374 93978
rect 273430 93922 273498 93978
rect 273554 93922 273622 93978
rect 273678 93922 273774 93978
rect 273154 76350 273774 93922
rect 273154 76294 273250 76350
rect 273306 76294 273374 76350
rect 273430 76294 273498 76350
rect 273554 76294 273622 76350
rect 273678 76294 273774 76350
rect 273154 76226 273774 76294
rect 273154 76170 273250 76226
rect 273306 76170 273374 76226
rect 273430 76170 273498 76226
rect 273554 76170 273622 76226
rect 273678 76170 273774 76226
rect 273154 76102 273774 76170
rect 273154 76046 273250 76102
rect 273306 76046 273374 76102
rect 273430 76046 273498 76102
rect 273554 76046 273622 76102
rect 273678 76046 273774 76102
rect 273154 75978 273774 76046
rect 273154 75922 273250 75978
rect 273306 75922 273374 75978
rect 273430 75922 273498 75978
rect 273554 75922 273622 75978
rect 273678 75922 273774 75978
rect 273154 58350 273774 75922
rect 273154 58294 273250 58350
rect 273306 58294 273374 58350
rect 273430 58294 273498 58350
rect 273554 58294 273622 58350
rect 273678 58294 273774 58350
rect 273154 58226 273774 58294
rect 273154 58170 273250 58226
rect 273306 58170 273374 58226
rect 273430 58170 273498 58226
rect 273554 58170 273622 58226
rect 273678 58170 273774 58226
rect 273154 58102 273774 58170
rect 273154 58046 273250 58102
rect 273306 58046 273374 58102
rect 273430 58046 273498 58102
rect 273554 58046 273622 58102
rect 273678 58046 273774 58102
rect 273154 57978 273774 58046
rect 273154 57922 273250 57978
rect 273306 57922 273374 57978
rect 273430 57922 273498 57978
rect 273554 57922 273622 57978
rect 273678 57922 273774 57978
rect 273154 40350 273774 57922
rect 273154 40294 273250 40350
rect 273306 40294 273374 40350
rect 273430 40294 273498 40350
rect 273554 40294 273622 40350
rect 273678 40294 273774 40350
rect 273154 40226 273774 40294
rect 273154 40170 273250 40226
rect 273306 40170 273374 40226
rect 273430 40170 273498 40226
rect 273554 40170 273622 40226
rect 273678 40170 273774 40226
rect 273154 40102 273774 40170
rect 273154 40046 273250 40102
rect 273306 40046 273374 40102
rect 273430 40046 273498 40102
rect 273554 40046 273622 40102
rect 273678 40046 273774 40102
rect 273154 39978 273774 40046
rect 273154 39922 273250 39978
rect 273306 39922 273374 39978
rect 273430 39922 273498 39978
rect 273554 39922 273622 39978
rect 273678 39922 273774 39978
rect 273154 22350 273774 39922
rect 273154 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 273774 22350
rect 273154 22226 273774 22294
rect 273154 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 273774 22226
rect 273154 22102 273774 22170
rect 273154 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 273774 22102
rect 273154 21978 273774 22046
rect 273154 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 273774 21978
rect 273154 4350 273774 21922
rect 273154 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 273774 4350
rect 273154 4226 273774 4294
rect 273154 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 273774 4226
rect 273154 4102 273774 4170
rect 273154 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 273774 4102
rect 273154 3978 273774 4046
rect 273154 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 273774 3978
rect 273154 -160 273774 3922
rect 273154 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 273774 -160
rect 273154 -284 273774 -216
rect 273154 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 273774 -284
rect 273154 -408 273774 -340
rect 273154 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 273774 -408
rect 273154 -532 273774 -464
rect 273154 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 273774 -532
rect 273154 -1644 273774 -588
rect 276874 208350 277494 210842
rect 276874 208294 276970 208350
rect 277026 208294 277094 208350
rect 277150 208294 277218 208350
rect 277274 208294 277342 208350
rect 277398 208294 277494 208350
rect 276874 208226 277494 208294
rect 276874 208170 276970 208226
rect 277026 208170 277094 208226
rect 277150 208170 277218 208226
rect 277274 208170 277342 208226
rect 277398 208170 277494 208226
rect 276874 208102 277494 208170
rect 276874 208046 276970 208102
rect 277026 208046 277094 208102
rect 277150 208046 277218 208102
rect 277274 208046 277342 208102
rect 277398 208046 277494 208102
rect 276874 207978 277494 208046
rect 276874 207922 276970 207978
rect 277026 207922 277094 207978
rect 277150 207922 277218 207978
rect 277274 207922 277342 207978
rect 277398 207922 277494 207978
rect 276874 190350 277494 207922
rect 281248 208350 281568 208384
rect 281248 208294 281318 208350
rect 281374 208294 281442 208350
rect 281498 208294 281568 208350
rect 281248 208226 281568 208294
rect 281248 208170 281318 208226
rect 281374 208170 281442 208226
rect 281498 208170 281568 208226
rect 281248 208102 281568 208170
rect 281248 208046 281318 208102
rect 281374 208046 281442 208102
rect 281498 208046 281568 208102
rect 281248 207978 281568 208046
rect 281248 207922 281318 207978
rect 281374 207922 281442 207978
rect 281498 207922 281568 207978
rect 281248 207888 281568 207922
rect 276874 190294 276970 190350
rect 277026 190294 277094 190350
rect 277150 190294 277218 190350
rect 277274 190294 277342 190350
rect 277398 190294 277494 190350
rect 276874 190226 277494 190294
rect 276874 190170 276970 190226
rect 277026 190170 277094 190226
rect 277150 190170 277218 190226
rect 277274 190170 277342 190226
rect 277398 190170 277494 190226
rect 276874 190102 277494 190170
rect 276874 190046 276970 190102
rect 277026 190046 277094 190102
rect 277150 190046 277218 190102
rect 277274 190046 277342 190102
rect 277398 190046 277494 190102
rect 276874 189978 277494 190046
rect 276874 189922 276970 189978
rect 277026 189922 277094 189978
rect 277150 189922 277218 189978
rect 277274 189922 277342 189978
rect 277398 189922 277494 189978
rect 276874 172350 277494 189922
rect 276874 172294 276970 172350
rect 277026 172294 277094 172350
rect 277150 172294 277218 172350
rect 277274 172294 277342 172350
rect 277398 172294 277494 172350
rect 276874 172226 277494 172294
rect 276874 172170 276970 172226
rect 277026 172170 277094 172226
rect 277150 172170 277218 172226
rect 277274 172170 277342 172226
rect 277398 172170 277494 172226
rect 276874 172102 277494 172170
rect 276874 172046 276970 172102
rect 277026 172046 277094 172102
rect 277150 172046 277218 172102
rect 277274 172046 277342 172102
rect 277398 172046 277494 172102
rect 276874 171978 277494 172046
rect 276874 171922 276970 171978
rect 277026 171922 277094 171978
rect 277150 171922 277218 171978
rect 277274 171922 277342 171978
rect 277398 171922 277494 171978
rect 276874 154350 277494 171922
rect 276874 154294 276970 154350
rect 277026 154294 277094 154350
rect 277150 154294 277218 154350
rect 277274 154294 277342 154350
rect 277398 154294 277494 154350
rect 276874 154226 277494 154294
rect 276874 154170 276970 154226
rect 277026 154170 277094 154226
rect 277150 154170 277218 154226
rect 277274 154170 277342 154226
rect 277398 154170 277494 154226
rect 276874 154102 277494 154170
rect 276874 154046 276970 154102
rect 277026 154046 277094 154102
rect 277150 154046 277218 154102
rect 277274 154046 277342 154102
rect 277398 154046 277494 154102
rect 276874 153978 277494 154046
rect 276874 153922 276970 153978
rect 277026 153922 277094 153978
rect 277150 153922 277218 153978
rect 277274 153922 277342 153978
rect 277398 153922 277494 153978
rect 276874 136350 277494 153922
rect 276874 136294 276970 136350
rect 277026 136294 277094 136350
rect 277150 136294 277218 136350
rect 277274 136294 277342 136350
rect 277398 136294 277494 136350
rect 276874 136226 277494 136294
rect 276874 136170 276970 136226
rect 277026 136170 277094 136226
rect 277150 136170 277218 136226
rect 277274 136170 277342 136226
rect 277398 136170 277494 136226
rect 276874 136102 277494 136170
rect 276874 136046 276970 136102
rect 277026 136046 277094 136102
rect 277150 136046 277218 136102
rect 277274 136046 277342 136102
rect 277398 136046 277494 136102
rect 276874 135978 277494 136046
rect 276874 135922 276970 135978
rect 277026 135922 277094 135978
rect 277150 135922 277218 135978
rect 277274 135922 277342 135978
rect 277398 135922 277494 135978
rect 276874 118350 277494 135922
rect 276874 118294 276970 118350
rect 277026 118294 277094 118350
rect 277150 118294 277218 118350
rect 277274 118294 277342 118350
rect 277398 118294 277494 118350
rect 276874 118226 277494 118294
rect 276874 118170 276970 118226
rect 277026 118170 277094 118226
rect 277150 118170 277218 118226
rect 277274 118170 277342 118226
rect 277398 118170 277494 118226
rect 276874 118102 277494 118170
rect 276874 118046 276970 118102
rect 277026 118046 277094 118102
rect 277150 118046 277218 118102
rect 277274 118046 277342 118102
rect 277398 118046 277494 118102
rect 276874 117978 277494 118046
rect 276874 117922 276970 117978
rect 277026 117922 277094 117978
rect 277150 117922 277218 117978
rect 277274 117922 277342 117978
rect 277398 117922 277494 117978
rect 276874 100350 277494 117922
rect 276874 100294 276970 100350
rect 277026 100294 277094 100350
rect 277150 100294 277218 100350
rect 277274 100294 277342 100350
rect 277398 100294 277494 100350
rect 276874 100226 277494 100294
rect 276874 100170 276970 100226
rect 277026 100170 277094 100226
rect 277150 100170 277218 100226
rect 277274 100170 277342 100226
rect 277398 100170 277494 100226
rect 276874 100102 277494 100170
rect 276874 100046 276970 100102
rect 277026 100046 277094 100102
rect 277150 100046 277218 100102
rect 277274 100046 277342 100102
rect 277398 100046 277494 100102
rect 276874 99978 277494 100046
rect 276874 99922 276970 99978
rect 277026 99922 277094 99978
rect 277150 99922 277218 99978
rect 277274 99922 277342 99978
rect 277398 99922 277494 99978
rect 276874 82350 277494 99922
rect 276874 82294 276970 82350
rect 277026 82294 277094 82350
rect 277150 82294 277218 82350
rect 277274 82294 277342 82350
rect 277398 82294 277494 82350
rect 276874 82226 277494 82294
rect 276874 82170 276970 82226
rect 277026 82170 277094 82226
rect 277150 82170 277218 82226
rect 277274 82170 277342 82226
rect 277398 82170 277494 82226
rect 276874 82102 277494 82170
rect 276874 82046 276970 82102
rect 277026 82046 277094 82102
rect 277150 82046 277218 82102
rect 277274 82046 277342 82102
rect 277398 82046 277494 82102
rect 276874 81978 277494 82046
rect 276874 81922 276970 81978
rect 277026 81922 277094 81978
rect 277150 81922 277218 81978
rect 277274 81922 277342 81978
rect 277398 81922 277494 81978
rect 276874 64350 277494 81922
rect 276874 64294 276970 64350
rect 277026 64294 277094 64350
rect 277150 64294 277218 64350
rect 277274 64294 277342 64350
rect 277398 64294 277494 64350
rect 276874 64226 277494 64294
rect 276874 64170 276970 64226
rect 277026 64170 277094 64226
rect 277150 64170 277218 64226
rect 277274 64170 277342 64226
rect 277398 64170 277494 64226
rect 276874 64102 277494 64170
rect 276874 64046 276970 64102
rect 277026 64046 277094 64102
rect 277150 64046 277218 64102
rect 277274 64046 277342 64102
rect 277398 64046 277494 64102
rect 276874 63978 277494 64046
rect 276874 63922 276970 63978
rect 277026 63922 277094 63978
rect 277150 63922 277218 63978
rect 277274 63922 277342 63978
rect 277398 63922 277494 63978
rect 276874 46350 277494 63922
rect 276874 46294 276970 46350
rect 277026 46294 277094 46350
rect 277150 46294 277218 46350
rect 277274 46294 277342 46350
rect 277398 46294 277494 46350
rect 276874 46226 277494 46294
rect 276874 46170 276970 46226
rect 277026 46170 277094 46226
rect 277150 46170 277218 46226
rect 277274 46170 277342 46226
rect 277398 46170 277494 46226
rect 276874 46102 277494 46170
rect 276874 46046 276970 46102
rect 277026 46046 277094 46102
rect 277150 46046 277218 46102
rect 277274 46046 277342 46102
rect 277398 46046 277494 46102
rect 276874 45978 277494 46046
rect 276874 45922 276970 45978
rect 277026 45922 277094 45978
rect 277150 45922 277218 45978
rect 277274 45922 277342 45978
rect 277398 45922 277494 45978
rect 276874 28350 277494 45922
rect 276874 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 277494 28350
rect 276874 28226 277494 28294
rect 276874 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 277494 28226
rect 276874 28102 277494 28170
rect 276874 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 277494 28102
rect 276874 27978 277494 28046
rect 276874 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 277494 27978
rect 276874 10350 277494 27922
rect 276874 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 277494 10350
rect 276874 10226 277494 10294
rect 276874 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 277494 10226
rect 276874 10102 277494 10170
rect 276874 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 277494 10102
rect 276874 9978 277494 10046
rect 276874 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 277494 9978
rect 276874 -1120 277494 9922
rect 276874 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 277494 -1120
rect 276874 -1244 277494 -1176
rect 276874 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 277494 -1244
rect 276874 -1368 277494 -1300
rect 276874 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 277494 -1368
rect 276874 -1492 277494 -1424
rect 276874 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 277494 -1492
rect 276874 -1644 277494 -1548
rect 291154 202350 291774 210842
rect 291154 202294 291250 202350
rect 291306 202294 291374 202350
rect 291430 202294 291498 202350
rect 291554 202294 291622 202350
rect 291678 202294 291774 202350
rect 291154 202226 291774 202294
rect 291154 202170 291250 202226
rect 291306 202170 291374 202226
rect 291430 202170 291498 202226
rect 291554 202170 291622 202226
rect 291678 202170 291774 202226
rect 291154 202102 291774 202170
rect 291154 202046 291250 202102
rect 291306 202046 291374 202102
rect 291430 202046 291498 202102
rect 291554 202046 291622 202102
rect 291678 202046 291774 202102
rect 291154 201978 291774 202046
rect 291154 201922 291250 201978
rect 291306 201922 291374 201978
rect 291430 201922 291498 201978
rect 291554 201922 291622 201978
rect 291678 201922 291774 201978
rect 291154 184350 291774 201922
rect 291154 184294 291250 184350
rect 291306 184294 291374 184350
rect 291430 184294 291498 184350
rect 291554 184294 291622 184350
rect 291678 184294 291774 184350
rect 291154 184226 291774 184294
rect 291154 184170 291250 184226
rect 291306 184170 291374 184226
rect 291430 184170 291498 184226
rect 291554 184170 291622 184226
rect 291678 184170 291774 184226
rect 291154 184102 291774 184170
rect 291154 184046 291250 184102
rect 291306 184046 291374 184102
rect 291430 184046 291498 184102
rect 291554 184046 291622 184102
rect 291678 184046 291774 184102
rect 291154 183978 291774 184046
rect 291154 183922 291250 183978
rect 291306 183922 291374 183978
rect 291430 183922 291498 183978
rect 291554 183922 291622 183978
rect 291678 183922 291774 183978
rect 291154 166350 291774 183922
rect 291154 166294 291250 166350
rect 291306 166294 291374 166350
rect 291430 166294 291498 166350
rect 291554 166294 291622 166350
rect 291678 166294 291774 166350
rect 291154 166226 291774 166294
rect 291154 166170 291250 166226
rect 291306 166170 291374 166226
rect 291430 166170 291498 166226
rect 291554 166170 291622 166226
rect 291678 166170 291774 166226
rect 291154 166102 291774 166170
rect 291154 166046 291250 166102
rect 291306 166046 291374 166102
rect 291430 166046 291498 166102
rect 291554 166046 291622 166102
rect 291678 166046 291774 166102
rect 291154 165978 291774 166046
rect 291154 165922 291250 165978
rect 291306 165922 291374 165978
rect 291430 165922 291498 165978
rect 291554 165922 291622 165978
rect 291678 165922 291774 165978
rect 291154 148350 291774 165922
rect 291154 148294 291250 148350
rect 291306 148294 291374 148350
rect 291430 148294 291498 148350
rect 291554 148294 291622 148350
rect 291678 148294 291774 148350
rect 291154 148226 291774 148294
rect 291154 148170 291250 148226
rect 291306 148170 291374 148226
rect 291430 148170 291498 148226
rect 291554 148170 291622 148226
rect 291678 148170 291774 148226
rect 291154 148102 291774 148170
rect 291154 148046 291250 148102
rect 291306 148046 291374 148102
rect 291430 148046 291498 148102
rect 291554 148046 291622 148102
rect 291678 148046 291774 148102
rect 291154 147978 291774 148046
rect 291154 147922 291250 147978
rect 291306 147922 291374 147978
rect 291430 147922 291498 147978
rect 291554 147922 291622 147978
rect 291678 147922 291774 147978
rect 291154 130350 291774 147922
rect 291154 130294 291250 130350
rect 291306 130294 291374 130350
rect 291430 130294 291498 130350
rect 291554 130294 291622 130350
rect 291678 130294 291774 130350
rect 291154 130226 291774 130294
rect 291154 130170 291250 130226
rect 291306 130170 291374 130226
rect 291430 130170 291498 130226
rect 291554 130170 291622 130226
rect 291678 130170 291774 130226
rect 291154 130102 291774 130170
rect 291154 130046 291250 130102
rect 291306 130046 291374 130102
rect 291430 130046 291498 130102
rect 291554 130046 291622 130102
rect 291678 130046 291774 130102
rect 291154 129978 291774 130046
rect 291154 129922 291250 129978
rect 291306 129922 291374 129978
rect 291430 129922 291498 129978
rect 291554 129922 291622 129978
rect 291678 129922 291774 129978
rect 291154 112350 291774 129922
rect 291154 112294 291250 112350
rect 291306 112294 291374 112350
rect 291430 112294 291498 112350
rect 291554 112294 291622 112350
rect 291678 112294 291774 112350
rect 291154 112226 291774 112294
rect 291154 112170 291250 112226
rect 291306 112170 291374 112226
rect 291430 112170 291498 112226
rect 291554 112170 291622 112226
rect 291678 112170 291774 112226
rect 291154 112102 291774 112170
rect 291154 112046 291250 112102
rect 291306 112046 291374 112102
rect 291430 112046 291498 112102
rect 291554 112046 291622 112102
rect 291678 112046 291774 112102
rect 291154 111978 291774 112046
rect 291154 111922 291250 111978
rect 291306 111922 291374 111978
rect 291430 111922 291498 111978
rect 291554 111922 291622 111978
rect 291678 111922 291774 111978
rect 291154 94350 291774 111922
rect 291154 94294 291250 94350
rect 291306 94294 291374 94350
rect 291430 94294 291498 94350
rect 291554 94294 291622 94350
rect 291678 94294 291774 94350
rect 291154 94226 291774 94294
rect 291154 94170 291250 94226
rect 291306 94170 291374 94226
rect 291430 94170 291498 94226
rect 291554 94170 291622 94226
rect 291678 94170 291774 94226
rect 291154 94102 291774 94170
rect 291154 94046 291250 94102
rect 291306 94046 291374 94102
rect 291430 94046 291498 94102
rect 291554 94046 291622 94102
rect 291678 94046 291774 94102
rect 291154 93978 291774 94046
rect 291154 93922 291250 93978
rect 291306 93922 291374 93978
rect 291430 93922 291498 93978
rect 291554 93922 291622 93978
rect 291678 93922 291774 93978
rect 291154 76350 291774 93922
rect 291154 76294 291250 76350
rect 291306 76294 291374 76350
rect 291430 76294 291498 76350
rect 291554 76294 291622 76350
rect 291678 76294 291774 76350
rect 291154 76226 291774 76294
rect 291154 76170 291250 76226
rect 291306 76170 291374 76226
rect 291430 76170 291498 76226
rect 291554 76170 291622 76226
rect 291678 76170 291774 76226
rect 291154 76102 291774 76170
rect 291154 76046 291250 76102
rect 291306 76046 291374 76102
rect 291430 76046 291498 76102
rect 291554 76046 291622 76102
rect 291678 76046 291774 76102
rect 291154 75978 291774 76046
rect 291154 75922 291250 75978
rect 291306 75922 291374 75978
rect 291430 75922 291498 75978
rect 291554 75922 291622 75978
rect 291678 75922 291774 75978
rect 291154 58350 291774 75922
rect 291154 58294 291250 58350
rect 291306 58294 291374 58350
rect 291430 58294 291498 58350
rect 291554 58294 291622 58350
rect 291678 58294 291774 58350
rect 291154 58226 291774 58294
rect 291154 58170 291250 58226
rect 291306 58170 291374 58226
rect 291430 58170 291498 58226
rect 291554 58170 291622 58226
rect 291678 58170 291774 58226
rect 291154 58102 291774 58170
rect 291154 58046 291250 58102
rect 291306 58046 291374 58102
rect 291430 58046 291498 58102
rect 291554 58046 291622 58102
rect 291678 58046 291774 58102
rect 291154 57978 291774 58046
rect 291154 57922 291250 57978
rect 291306 57922 291374 57978
rect 291430 57922 291498 57978
rect 291554 57922 291622 57978
rect 291678 57922 291774 57978
rect 291154 40350 291774 57922
rect 291154 40294 291250 40350
rect 291306 40294 291374 40350
rect 291430 40294 291498 40350
rect 291554 40294 291622 40350
rect 291678 40294 291774 40350
rect 291154 40226 291774 40294
rect 291154 40170 291250 40226
rect 291306 40170 291374 40226
rect 291430 40170 291498 40226
rect 291554 40170 291622 40226
rect 291678 40170 291774 40226
rect 291154 40102 291774 40170
rect 291154 40046 291250 40102
rect 291306 40046 291374 40102
rect 291430 40046 291498 40102
rect 291554 40046 291622 40102
rect 291678 40046 291774 40102
rect 291154 39978 291774 40046
rect 291154 39922 291250 39978
rect 291306 39922 291374 39978
rect 291430 39922 291498 39978
rect 291554 39922 291622 39978
rect 291678 39922 291774 39978
rect 291154 22350 291774 39922
rect 291154 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 291774 22350
rect 291154 22226 291774 22294
rect 291154 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 291774 22226
rect 291154 22102 291774 22170
rect 291154 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 291774 22102
rect 291154 21978 291774 22046
rect 291154 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 291774 21978
rect 291154 4350 291774 21922
rect 291154 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 291774 4350
rect 291154 4226 291774 4294
rect 291154 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 291774 4226
rect 291154 4102 291774 4170
rect 291154 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 291774 4102
rect 291154 3978 291774 4046
rect 291154 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 291774 3978
rect 291154 -160 291774 3922
rect 291154 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 291774 -160
rect 291154 -284 291774 -216
rect 291154 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 291774 -284
rect 291154 -408 291774 -340
rect 291154 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 291774 -408
rect 291154 -532 291774 -464
rect 291154 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 291774 -532
rect 291154 -1644 291774 -588
rect 294874 208350 295494 210842
rect 294874 208294 294970 208350
rect 295026 208294 295094 208350
rect 295150 208294 295218 208350
rect 295274 208294 295342 208350
rect 295398 208294 295494 208350
rect 294874 208226 295494 208294
rect 294874 208170 294970 208226
rect 295026 208170 295094 208226
rect 295150 208170 295218 208226
rect 295274 208170 295342 208226
rect 295398 208170 295494 208226
rect 294874 208102 295494 208170
rect 294874 208046 294970 208102
rect 295026 208046 295094 208102
rect 295150 208046 295218 208102
rect 295274 208046 295342 208102
rect 295398 208046 295494 208102
rect 294874 207978 295494 208046
rect 294874 207922 294970 207978
rect 295026 207922 295094 207978
rect 295150 207922 295218 207978
rect 295274 207922 295342 207978
rect 295398 207922 295494 207978
rect 294874 190350 295494 207922
rect 294874 190294 294970 190350
rect 295026 190294 295094 190350
rect 295150 190294 295218 190350
rect 295274 190294 295342 190350
rect 295398 190294 295494 190350
rect 294874 190226 295494 190294
rect 294874 190170 294970 190226
rect 295026 190170 295094 190226
rect 295150 190170 295218 190226
rect 295274 190170 295342 190226
rect 295398 190170 295494 190226
rect 294874 190102 295494 190170
rect 294874 190046 294970 190102
rect 295026 190046 295094 190102
rect 295150 190046 295218 190102
rect 295274 190046 295342 190102
rect 295398 190046 295494 190102
rect 294874 189978 295494 190046
rect 294874 189922 294970 189978
rect 295026 189922 295094 189978
rect 295150 189922 295218 189978
rect 295274 189922 295342 189978
rect 295398 189922 295494 189978
rect 294874 172350 295494 189922
rect 294874 172294 294970 172350
rect 295026 172294 295094 172350
rect 295150 172294 295218 172350
rect 295274 172294 295342 172350
rect 295398 172294 295494 172350
rect 294874 172226 295494 172294
rect 294874 172170 294970 172226
rect 295026 172170 295094 172226
rect 295150 172170 295218 172226
rect 295274 172170 295342 172226
rect 295398 172170 295494 172226
rect 294874 172102 295494 172170
rect 294874 172046 294970 172102
rect 295026 172046 295094 172102
rect 295150 172046 295218 172102
rect 295274 172046 295342 172102
rect 295398 172046 295494 172102
rect 294874 171978 295494 172046
rect 294874 171922 294970 171978
rect 295026 171922 295094 171978
rect 295150 171922 295218 171978
rect 295274 171922 295342 171978
rect 295398 171922 295494 171978
rect 294874 154350 295494 171922
rect 294874 154294 294970 154350
rect 295026 154294 295094 154350
rect 295150 154294 295218 154350
rect 295274 154294 295342 154350
rect 295398 154294 295494 154350
rect 294874 154226 295494 154294
rect 294874 154170 294970 154226
rect 295026 154170 295094 154226
rect 295150 154170 295218 154226
rect 295274 154170 295342 154226
rect 295398 154170 295494 154226
rect 294874 154102 295494 154170
rect 294874 154046 294970 154102
rect 295026 154046 295094 154102
rect 295150 154046 295218 154102
rect 295274 154046 295342 154102
rect 295398 154046 295494 154102
rect 294874 153978 295494 154046
rect 294874 153922 294970 153978
rect 295026 153922 295094 153978
rect 295150 153922 295218 153978
rect 295274 153922 295342 153978
rect 295398 153922 295494 153978
rect 294874 136350 295494 153922
rect 294874 136294 294970 136350
rect 295026 136294 295094 136350
rect 295150 136294 295218 136350
rect 295274 136294 295342 136350
rect 295398 136294 295494 136350
rect 294874 136226 295494 136294
rect 294874 136170 294970 136226
rect 295026 136170 295094 136226
rect 295150 136170 295218 136226
rect 295274 136170 295342 136226
rect 295398 136170 295494 136226
rect 294874 136102 295494 136170
rect 294874 136046 294970 136102
rect 295026 136046 295094 136102
rect 295150 136046 295218 136102
rect 295274 136046 295342 136102
rect 295398 136046 295494 136102
rect 294874 135978 295494 136046
rect 294874 135922 294970 135978
rect 295026 135922 295094 135978
rect 295150 135922 295218 135978
rect 295274 135922 295342 135978
rect 295398 135922 295494 135978
rect 294874 118350 295494 135922
rect 294874 118294 294970 118350
rect 295026 118294 295094 118350
rect 295150 118294 295218 118350
rect 295274 118294 295342 118350
rect 295398 118294 295494 118350
rect 294874 118226 295494 118294
rect 294874 118170 294970 118226
rect 295026 118170 295094 118226
rect 295150 118170 295218 118226
rect 295274 118170 295342 118226
rect 295398 118170 295494 118226
rect 294874 118102 295494 118170
rect 294874 118046 294970 118102
rect 295026 118046 295094 118102
rect 295150 118046 295218 118102
rect 295274 118046 295342 118102
rect 295398 118046 295494 118102
rect 294874 117978 295494 118046
rect 294874 117922 294970 117978
rect 295026 117922 295094 117978
rect 295150 117922 295218 117978
rect 295274 117922 295342 117978
rect 295398 117922 295494 117978
rect 294874 100350 295494 117922
rect 294874 100294 294970 100350
rect 295026 100294 295094 100350
rect 295150 100294 295218 100350
rect 295274 100294 295342 100350
rect 295398 100294 295494 100350
rect 294874 100226 295494 100294
rect 294874 100170 294970 100226
rect 295026 100170 295094 100226
rect 295150 100170 295218 100226
rect 295274 100170 295342 100226
rect 295398 100170 295494 100226
rect 294874 100102 295494 100170
rect 294874 100046 294970 100102
rect 295026 100046 295094 100102
rect 295150 100046 295218 100102
rect 295274 100046 295342 100102
rect 295398 100046 295494 100102
rect 294874 99978 295494 100046
rect 294874 99922 294970 99978
rect 295026 99922 295094 99978
rect 295150 99922 295218 99978
rect 295274 99922 295342 99978
rect 295398 99922 295494 99978
rect 294874 82350 295494 99922
rect 294874 82294 294970 82350
rect 295026 82294 295094 82350
rect 295150 82294 295218 82350
rect 295274 82294 295342 82350
rect 295398 82294 295494 82350
rect 294874 82226 295494 82294
rect 294874 82170 294970 82226
rect 295026 82170 295094 82226
rect 295150 82170 295218 82226
rect 295274 82170 295342 82226
rect 295398 82170 295494 82226
rect 294874 82102 295494 82170
rect 294874 82046 294970 82102
rect 295026 82046 295094 82102
rect 295150 82046 295218 82102
rect 295274 82046 295342 82102
rect 295398 82046 295494 82102
rect 294874 81978 295494 82046
rect 294874 81922 294970 81978
rect 295026 81922 295094 81978
rect 295150 81922 295218 81978
rect 295274 81922 295342 81978
rect 295398 81922 295494 81978
rect 294874 64350 295494 81922
rect 294874 64294 294970 64350
rect 295026 64294 295094 64350
rect 295150 64294 295218 64350
rect 295274 64294 295342 64350
rect 295398 64294 295494 64350
rect 294874 64226 295494 64294
rect 294874 64170 294970 64226
rect 295026 64170 295094 64226
rect 295150 64170 295218 64226
rect 295274 64170 295342 64226
rect 295398 64170 295494 64226
rect 294874 64102 295494 64170
rect 294874 64046 294970 64102
rect 295026 64046 295094 64102
rect 295150 64046 295218 64102
rect 295274 64046 295342 64102
rect 295398 64046 295494 64102
rect 294874 63978 295494 64046
rect 294874 63922 294970 63978
rect 295026 63922 295094 63978
rect 295150 63922 295218 63978
rect 295274 63922 295342 63978
rect 295398 63922 295494 63978
rect 294874 46350 295494 63922
rect 294874 46294 294970 46350
rect 295026 46294 295094 46350
rect 295150 46294 295218 46350
rect 295274 46294 295342 46350
rect 295398 46294 295494 46350
rect 294874 46226 295494 46294
rect 294874 46170 294970 46226
rect 295026 46170 295094 46226
rect 295150 46170 295218 46226
rect 295274 46170 295342 46226
rect 295398 46170 295494 46226
rect 294874 46102 295494 46170
rect 294874 46046 294970 46102
rect 295026 46046 295094 46102
rect 295150 46046 295218 46102
rect 295274 46046 295342 46102
rect 295398 46046 295494 46102
rect 294874 45978 295494 46046
rect 294874 45922 294970 45978
rect 295026 45922 295094 45978
rect 295150 45922 295218 45978
rect 295274 45922 295342 45978
rect 295398 45922 295494 45978
rect 294874 28350 295494 45922
rect 294874 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 295494 28350
rect 294874 28226 295494 28294
rect 294874 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 295494 28226
rect 294874 28102 295494 28170
rect 294874 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 295494 28102
rect 294874 27978 295494 28046
rect 294874 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 295494 27978
rect 294874 10350 295494 27922
rect 294874 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 295494 10350
rect 294874 10226 295494 10294
rect 294874 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 295494 10226
rect 294874 10102 295494 10170
rect 294874 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 295494 10102
rect 294874 9978 295494 10046
rect 294874 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 295494 9978
rect 294874 -1120 295494 9922
rect 294874 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 295494 -1120
rect 294874 -1244 295494 -1176
rect 294874 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 295494 -1244
rect 294874 -1368 295494 -1300
rect 294874 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 295494 -1368
rect 294874 -1492 295494 -1424
rect 294874 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 295494 -1492
rect 294874 -1644 295494 -1548
rect 309154 202350 309774 210842
rect 311968 208350 312288 208384
rect 311968 208294 312038 208350
rect 312094 208294 312162 208350
rect 312218 208294 312288 208350
rect 311968 208226 312288 208294
rect 311968 208170 312038 208226
rect 312094 208170 312162 208226
rect 312218 208170 312288 208226
rect 311968 208102 312288 208170
rect 311968 208046 312038 208102
rect 312094 208046 312162 208102
rect 312218 208046 312288 208102
rect 311968 207978 312288 208046
rect 311968 207922 312038 207978
rect 312094 207922 312162 207978
rect 312218 207922 312288 207978
rect 311968 207888 312288 207922
rect 312874 208350 313494 210842
rect 312874 208294 312970 208350
rect 313026 208294 313094 208350
rect 313150 208294 313218 208350
rect 313274 208294 313342 208350
rect 313398 208294 313494 208350
rect 312874 208226 313494 208294
rect 312874 208170 312970 208226
rect 313026 208170 313094 208226
rect 313150 208170 313218 208226
rect 313274 208170 313342 208226
rect 313398 208170 313494 208226
rect 312874 208102 313494 208170
rect 312874 208046 312970 208102
rect 313026 208046 313094 208102
rect 313150 208046 313218 208102
rect 313274 208046 313342 208102
rect 313398 208046 313494 208102
rect 312874 207978 313494 208046
rect 312874 207922 312970 207978
rect 313026 207922 313094 207978
rect 313150 207922 313218 207978
rect 313274 207922 313342 207978
rect 313398 207922 313494 207978
rect 309154 202294 309250 202350
rect 309306 202294 309374 202350
rect 309430 202294 309498 202350
rect 309554 202294 309622 202350
rect 309678 202294 309774 202350
rect 309154 202226 309774 202294
rect 309154 202170 309250 202226
rect 309306 202170 309374 202226
rect 309430 202170 309498 202226
rect 309554 202170 309622 202226
rect 309678 202170 309774 202226
rect 309154 202102 309774 202170
rect 309154 202046 309250 202102
rect 309306 202046 309374 202102
rect 309430 202046 309498 202102
rect 309554 202046 309622 202102
rect 309678 202046 309774 202102
rect 309154 201978 309774 202046
rect 309154 201922 309250 201978
rect 309306 201922 309374 201978
rect 309430 201922 309498 201978
rect 309554 201922 309622 201978
rect 309678 201922 309774 201978
rect 309154 184350 309774 201922
rect 309154 184294 309250 184350
rect 309306 184294 309374 184350
rect 309430 184294 309498 184350
rect 309554 184294 309622 184350
rect 309678 184294 309774 184350
rect 309154 184226 309774 184294
rect 309154 184170 309250 184226
rect 309306 184170 309374 184226
rect 309430 184170 309498 184226
rect 309554 184170 309622 184226
rect 309678 184170 309774 184226
rect 309154 184102 309774 184170
rect 309154 184046 309250 184102
rect 309306 184046 309374 184102
rect 309430 184046 309498 184102
rect 309554 184046 309622 184102
rect 309678 184046 309774 184102
rect 309154 183978 309774 184046
rect 309154 183922 309250 183978
rect 309306 183922 309374 183978
rect 309430 183922 309498 183978
rect 309554 183922 309622 183978
rect 309678 183922 309774 183978
rect 309154 166350 309774 183922
rect 309154 166294 309250 166350
rect 309306 166294 309374 166350
rect 309430 166294 309498 166350
rect 309554 166294 309622 166350
rect 309678 166294 309774 166350
rect 309154 166226 309774 166294
rect 309154 166170 309250 166226
rect 309306 166170 309374 166226
rect 309430 166170 309498 166226
rect 309554 166170 309622 166226
rect 309678 166170 309774 166226
rect 309154 166102 309774 166170
rect 309154 166046 309250 166102
rect 309306 166046 309374 166102
rect 309430 166046 309498 166102
rect 309554 166046 309622 166102
rect 309678 166046 309774 166102
rect 309154 165978 309774 166046
rect 309154 165922 309250 165978
rect 309306 165922 309374 165978
rect 309430 165922 309498 165978
rect 309554 165922 309622 165978
rect 309678 165922 309774 165978
rect 309154 148350 309774 165922
rect 309154 148294 309250 148350
rect 309306 148294 309374 148350
rect 309430 148294 309498 148350
rect 309554 148294 309622 148350
rect 309678 148294 309774 148350
rect 309154 148226 309774 148294
rect 309154 148170 309250 148226
rect 309306 148170 309374 148226
rect 309430 148170 309498 148226
rect 309554 148170 309622 148226
rect 309678 148170 309774 148226
rect 309154 148102 309774 148170
rect 309154 148046 309250 148102
rect 309306 148046 309374 148102
rect 309430 148046 309498 148102
rect 309554 148046 309622 148102
rect 309678 148046 309774 148102
rect 309154 147978 309774 148046
rect 309154 147922 309250 147978
rect 309306 147922 309374 147978
rect 309430 147922 309498 147978
rect 309554 147922 309622 147978
rect 309678 147922 309774 147978
rect 309154 130350 309774 147922
rect 309154 130294 309250 130350
rect 309306 130294 309374 130350
rect 309430 130294 309498 130350
rect 309554 130294 309622 130350
rect 309678 130294 309774 130350
rect 309154 130226 309774 130294
rect 309154 130170 309250 130226
rect 309306 130170 309374 130226
rect 309430 130170 309498 130226
rect 309554 130170 309622 130226
rect 309678 130170 309774 130226
rect 309154 130102 309774 130170
rect 309154 130046 309250 130102
rect 309306 130046 309374 130102
rect 309430 130046 309498 130102
rect 309554 130046 309622 130102
rect 309678 130046 309774 130102
rect 309154 129978 309774 130046
rect 309154 129922 309250 129978
rect 309306 129922 309374 129978
rect 309430 129922 309498 129978
rect 309554 129922 309622 129978
rect 309678 129922 309774 129978
rect 309154 112350 309774 129922
rect 309154 112294 309250 112350
rect 309306 112294 309374 112350
rect 309430 112294 309498 112350
rect 309554 112294 309622 112350
rect 309678 112294 309774 112350
rect 309154 112226 309774 112294
rect 309154 112170 309250 112226
rect 309306 112170 309374 112226
rect 309430 112170 309498 112226
rect 309554 112170 309622 112226
rect 309678 112170 309774 112226
rect 309154 112102 309774 112170
rect 309154 112046 309250 112102
rect 309306 112046 309374 112102
rect 309430 112046 309498 112102
rect 309554 112046 309622 112102
rect 309678 112046 309774 112102
rect 309154 111978 309774 112046
rect 309154 111922 309250 111978
rect 309306 111922 309374 111978
rect 309430 111922 309498 111978
rect 309554 111922 309622 111978
rect 309678 111922 309774 111978
rect 309154 94350 309774 111922
rect 309154 94294 309250 94350
rect 309306 94294 309374 94350
rect 309430 94294 309498 94350
rect 309554 94294 309622 94350
rect 309678 94294 309774 94350
rect 309154 94226 309774 94294
rect 309154 94170 309250 94226
rect 309306 94170 309374 94226
rect 309430 94170 309498 94226
rect 309554 94170 309622 94226
rect 309678 94170 309774 94226
rect 309154 94102 309774 94170
rect 309154 94046 309250 94102
rect 309306 94046 309374 94102
rect 309430 94046 309498 94102
rect 309554 94046 309622 94102
rect 309678 94046 309774 94102
rect 309154 93978 309774 94046
rect 309154 93922 309250 93978
rect 309306 93922 309374 93978
rect 309430 93922 309498 93978
rect 309554 93922 309622 93978
rect 309678 93922 309774 93978
rect 309154 76350 309774 93922
rect 309154 76294 309250 76350
rect 309306 76294 309374 76350
rect 309430 76294 309498 76350
rect 309554 76294 309622 76350
rect 309678 76294 309774 76350
rect 309154 76226 309774 76294
rect 309154 76170 309250 76226
rect 309306 76170 309374 76226
rect 309430 76170 309498 76226
rect 309554 76170 309622 76226
rect 309678 76170 309774 76226
rect 309154 76102 309774 76170
rect 309154 76046 309250 76102
rect 309306 76046 309374 76102
rect 309430 76046 309498 76102
rect 309554 76046 309622 76102
rect 309678 76046 309774 76102
rect 309154 75978 309774 76046
rect 309154 75922 309250 75978
rect 309306 75922 309374 75978
rect 309430 75922 309498 75978
rect 309554 75922 309622 75978
rect 309678 75922 309774 75978
rect 309154 58350 309774 75922
rect 309154 58294 309250 58350
rect 309306 58294 309374 58350
rect 309430 58294 309498 58350
rect 309554 58294 309622 58350
rect 309678 58294 309774 58350
rect 309154 58226 309774 58294
rect 309154 58170 309250 58226
rect 309306 58170 309374 58226
rect 309430 58170 309498 58226
rect 309554 58170 309622 58226
rect 309678 58170 309774 58226
rect 309154 58102 309774 58170
rect 309154 58046 309250 58102
rect 309306 58046 309374 58102
rect 309430 58046 309498 58102
rect 309554 58046 309622 58102
rect 309678 58046 309774 58102
rect 309154 57978 309774 58046
rect 309154 57922 309250 57978
rect 309306 57922 309374 57978
rect 309430 57922 309498 57978
rect 309554 57922 309622 57978
rect 309678 57922 309774 57978
rect 309154 40350 309774 57922
rect 309154 40294 309250 40350
rect 309306 40294 309374 40350
rect 309430 40294 309498 40350
rect 309554 40294 309622 40350
rect 309678 40294 309774 40350
rect 309154 40226 309774 40294
rect 309154 40170 309250 40226
rect 309306 40170 309374 40226
rect 309430 40170 309498 40226
rect 309554 40170 309622 40226
rect 309678 40170 309774 40226
rect 309154 40102 309774 40170
rect 309154 40046 309250 40102
rect 309306 40046 309374 40102
rect 309430 40046 309498 40102
rect 309554 40046 309622 40102
rect 309678 40046 309774 40102
rect 309154 39978 309774 40046
rect 309154 39922 309250 39978
rect 309306 39922 309374 39978
rect 309430 39922 309498 39978
rect 309554 39922 309622 39978
rect 309678 39922 309774 39978
rect 309154 22350 309774 39922
rect 309154 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 309774 22350
rect 309154 22226 309774 22294
rect 309154 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 309774 22226
rect 309154 22102 309774 22170
rect 309154 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 309774 22102
rect 309154 21978 309774 22046
rect 309154 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 309774 21978
rect 309154 4350 309774 21922
rect 309154 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 309774 4350
rect 309154 4226 309774 4294
rect 309154 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 309774 4226
rect 309154 4102 309774 4170
rect 309154 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 309774 4102
rect 309154 3978 309774 4046
rect 309154 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 309774 3978
rect 309154 -160 309774 3922
rect 309154 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 309774 -160
rect 309154 -284 309774 -216
rect 309154 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 309774 -284
rect 309154 -408 309774 -340
rect 309154 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 309774 -408
rect 309154 -532 309774 -464
rect 309154 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 309774 -532
rect 309154 -1644 309774 -588
rect 312874 190350 313494 207922
rect 330874 208350 331494 210842
rect 330874 208294 330970 208350
rect 331026 208294 331094 208350
rect 331150 208294 331218 208350
rect 331274 208294 331342 208350
rect 331398 208294 331494 208350
rect 330874 208226 331494 208294
rect 330874 208170 330970 208226
rect 331026 208170 331094 208226
rect 331150 208170 331218 208226
rect 331274 208170 331342 208226
rect 331398 208170 331494 208226
rect 330874 208102 331494 208170
rect 330874 208046 330970 208102
rect 331026 208046 331094 208102
rect 331150 208046 331218 208102
rect 331274 208046 331342 208102
rect 331398 208046 331494 208102
rect 330874 207978 331494 208046
rect 330874 207922 330970 207978
rect 331026 207922 331094 207978
rect 331150 207922 331218 207978
rect 331274 207922 331342 207978
rect 331398 207922 331494 207978
rect 312874 190294 312970 190350
rect 313026 190294 313094 190350
rect 313150 190294 313218 190350
rect 313274 190294 313342 190350
rect 313398 190294 313494 190350
rect 312874 190226 313494 190294
rect 312874 190170 312970 190226
rect 313026 190170 313094 190226
rect 313150 190170 313218 190226
rect 313274 190170 313342 190226
rect 313398 190170 313494 190226
rect 312874 190102 313494 190170
rect 312874 190046 312970 190102
rect 313026 190046 313094 190102
rect 313150 190046 313218 190102
rect 313274 190046 313342 190102
rect 313398 190046 313494 190102
rect 312874 189978 313494 190046
rect 312874 189922 312970 189978
rect 313026 189922 313094 189978
rect 313150 189922 313218 189978
rect 313274 189922 313342 189978
rect 313398 189922 313494 189978
rect 312874 172350 313494 189922
rect 312874 172294 312970 172350
rect 313026 172294 313094 172350
rect 313150 172294 313218 172350
rect 313274 172294 313342 172350
rect 313398 172294 313494 172350
rect 312874 172226 313494 172294
rect 312874 172170 312970 172226
rect 313026 172170 313094 172226
rect 313150 172170 313218 172226
rect 313274 172170 313342 172226
rect 313398 172170 313494 172226
rect 312874 172102 313494 172170
rect 312874 172046 312970 172102
rect 313026 172046 313094 172102
rect 313150 172046 313218 172102
rect 313274 172046 313342 172102
rect 313398 172046 313494 172102
rect 312874 171978 313494 172046
rect 312874 171922 312970 171978
rect 313026 171922 313094 171978
rect 313150 171922 313218 171978
rect 313274 171922 313342 171978
rect 313398 171922 313494 171978
rect 312874 154350 313494 171922
rect 312874 154294 312970 154350
rect 313026 154294 313094 154350
rect 313150 154294 313218 154350
rect 313274 154294 313342 154350
rect 313398 154294 313494 154350
rect 312874 154226 313494 154294
rect 312874 154170 312970 154226
rect 313026 154170 313094 154226
rect 313150 154170 313218 154226
rect 313274 154170 313342 154226
rect 313398 154170 313494 154226
rect 312874 154102 313494 154170
rect 312874 154046 312970 154102
rect 313026 154046 313094 154102
rect 313150 154046 313218 154102
rect 313274 154046 313342 154102
rect 313398 154046 313494 154102
rect 312874 153978 313494 154046
rect 312874 153922 312970 153978
rect 313026 153922 313094 153978
rect 313150 153922 313218 153978
rect 313274 153922 313342 153978
rect 313398 153922 313494 153978
rect 312874 136350 313494 153922
rect 312874 136294 312970 136350
rect 313026 136294 313094 136350
rect 313150 136294 313218 136350
rect 313274 136294 313342 136350
rect 313398 136294 313494 136350
rect 312874 136226 313494 136294
rect 312874 136170 312970 136226
rect 313026 136170 313094 136226
rect 313150 136170 313218 136226
rect 313274 136170 313342 136226
rect 313398 136170 313494 136226
rect 312874 136102 313494 136170
rect 312874 136046 312970 136102
rect 313026 136046 313094 136102
rect 313150 136046 313218 136102
rect 313274 136046 313342 136102
rect 313398 136046 313494 136102
rect 312874 135978 313494 136046
rect 312874 135922 312970 135978
rect 313026 135922 313094 135978
rect 313150 135922 313218 135978
rect 313274 135922 313342 135978
rect 313398 135922 313494 135978
rect 312874 118350 313494 135922
rect 312874 118294 312970 118350
rect 313026 118294 313094 118350
rect 313150 118294 313218 118350
rect 313274 118294 313342 118350
rect 313398 118294 313494 118350
rect 312874 118226 313494 118294
rect 312874 118170 312970 118226
rect 313026 118170 313094 118226
rect 313150 118170 313218 118226
rect 313274 118170 313342 118226
rect 313398 118170 313494 118226
rect 312874 118102 313494 118170
rect 312874 118046 312970 118102
rect 313026 118046 313094 118102
rect 313150 118046 313218 118102
rect 313274 118046 313342 118102
rect 313398 118046 313494 118102
rect 312874 117978 313494 118046
rect 312874 117922 312970 117978
rect 313026 117922 313094 117978
rect 313150 117922 313218 117978
rect 313274 117922 313342 117978
rect 313398 117922 313494 117978
rect 312874 100350 313494 117922
rect 312874 100294 312970 100350
rect 313026 100294 313094 100350
rect 313150 100294 313218 100350
rect 313274 100294 313342 100350
rect 313398 100294 313494 100350
rect 312874 100226 313494 100294
rect 312874 100170 312970 100226
rect 313026 100170 313094 100226
rect 313150 100170 313218 100226
rect 313274 100170 313342 100226
rect 313398 100170 313494 100226
rect 312874 100102 313494 100170
rect 312874 100046 312970 100102
rect 313026 100046 313094 100102
rect 313150 100046 313218 100102
rect 313274 100046 313342 100102
rect 313398 100046 313494 100102
rect 312874 99978 313494 100046
rect 312874 99922 312970 99978
rect 313026 99922 313094 99978
rect 313150 99922 313218 99978
rect 313274 99922 313342 99978
rect 313398 99922 313494 99978
rect 312874 82350 313494 99922
rect 312874 82294 312970 82350
rect 313026 82294 313094 82350
rect 313150 82294 313218 82350
rect 313274 82294 313342 82350
rect 313398 82294 313494 82350
rect 312874 82226 313494 82294
rect 312874 82170 312970 82226
rect 313026 82170 313094 82226
rect 313150 82170 313218 82226
rect 313274 82170 313342 82226
rect 313398 82170 313494 82226
rect 312874 82102 313494 82170
rect 312874 82046 312970 82102
rect 313026 82046 313094 82102
rect 313150 82046 313218 82102
rect 313274 82046 313342 82102
rect 313398 82046 313494 82102
rect 312874 81978 313494 82046
rect 312874 81922 312970 81978
rect 313026 81922 313094 81978
rect 313150 81922 313218 81978
rect 313274 81922 313342 81978
rect 313398 81922 313494 81978
rect 312874 64350 313494 81922
rect 312874 64294 312970 64350
rect 313026 64294 313094 64350
rect 313150 64294 313218 64350
rect 313274 64294 313342 64350
rect 313398 64294 313494 64350
rect 312874 64226 313494 64294
rect 312874 64170 312970 64226
rect 313026 64170 313094 64226
rect 313150 64170 313218 64226
rect 313274 64170 313342 64226
rect 313398 64170 313494 64226
rect 312874 64102 313494 64170
rect 312874 64046 312970 64102
rect 313026 64046 313094 64102
rect 313150 64046 313218 64102
rect 313274 64046 313342 64102
rect 313398 64046 313494 64102
rect 312874 63978 313494 64046
rect 312874 63922 312970 63978
rect 313026 63922 313094 63978
rect 313150 63922 313218 63978
rect 313274 63922 313342 63978
rect 313398 63922 313494 63978
rect 312874 46350 313494 63922
rect 312874 46294 312970 46350
rect 313026 46294 313094 46350
rect 313150 46294 313218 46350
rect 313274 46294 313342 46350
rect 313398 46294 313494 46350
rect 312874 46226 313494 46294
rect 312874 46170 312970 46226
rect 313026 46170 313094 46226
rect 313150 46170 313218 46226
rect 313274 46170 313342 46226
rect 313398 46170 313494 46226
rect 312874 46102 313494 46170
rect 312874 46046 312970 46102
rect 313026 46046 313094 46102
rect 313150 46046 313218 46102
rect 313274 46046 313342 46102
rect 313398 46046 313494 46102
rect 312874 45978 313494 46046
rect 312874 45922 312970 45978
rect 313026 45922 313094 45978
rect 313150 45922 313218 45978
rect 313274 45922 313342 45978
rect 313398 45922 313494 45978
rect 312874 28350 313494 45922
rect 312874 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 313494 28350
rect 312874 28226 313494 28294
rect 312874 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 313494 28226
rect 312874 28102 313494 28170
rect 312874 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 313494 28102
rect 312874 27978 313494 28046
rect 312874 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 313494 27978
rect 312874 10350 313494 27922
rect 312874 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 313494 10350
rect 312874 10226 313494 10294
rect 312874 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 313494 10226
rect 312874 10102 313494 10170
rect 312874 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 313494 10102
rect 312874 9978 313494 10046
rect 312874 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 313494 9978
rect 312874 -1120 313494 9922
rect 312874 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 313494 -1120
rect 312874 -1244 313494 -1176
rect 312874 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 313494 -1244
rect 312874 -1368 313494 -1300
rect 312874 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 313494 -1368
rect 312874 -1492 313494 -1424
rect 312874 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 313494 -1492
rect 312874 -1644 313494 -1548
rect 327154 184350 327774 201020
rect 327154 184294 327250 184350
rect 327306 184294 327374 184350
rect 327430 184294 327498 184350
rect 327554 184294 327622 184350
rect 327678 184294 327774 184350
rect 327154 184226 327774 184294
rect 327154 184170 327250 184226
rect 327306 184170 327374 184226
rect 327430 184170 327498 184226
rect 327554 184170 327622 184226
rect 327678 184170 327774 184226
rect 327154 184102 327774 184170
rect 327154 184046 327250 184102
rect 327306 184046 327374 184102
rect 327430 184046 327498 184102
rect 327554 184046 327622 184102
rect 327678 184046 327774 184102
rect 327154 183978 327774 184046
rect 327154 183922 327250 183978
rect 327306 183922 327374 183978
rect 327430 183922 327498 183978
rect 327554 183922 327622 183978
rect 327678 183922 327774 183978
rect 327154 166350 327774 183922
rect 327154 166294 327250 166350
rect 327306 166294 327374 166350
rect 327430 166294 327498 166350
rect 327554 166294 327622 166350
rect 327678 166294 327774 166350
rect 327154 166226 327774 166294
rect 327154 166170 327250 166226
rect 327306 166170 327374 166226
rect 327430 166170 327498 166226
rect 327554 166170 327622 166226
rect 327678 166170 327774 166226
rect 327154 166102 327774 166170
rect 327154 166046 327250 166102
rect 327306 166046 327374 166102
rect 327430 166046 327498 166102
rect 327554 166046 327622 166102
rect 327678 166046 327774 166102
rect 327154 165978 327774 166046
rect 327154 165922 327250 165978
rect 327306 165922 327374 165978
rect 327430 165922 327498 165978
rect 327554 165922 327622 165978
rect 327678 165922 327774 165978
rect 327154 148350 327774 165922
rect 327154 148294 327250 148350
rect 327306 148294 327374 148350
rect 327430 148294 327498 148350
rect 327554 148294 327622 148350
rect 327678 148294 327774 148350
rect 327154 148226 327774 148294
rect 327154 148170 327250 148226
rect 327306 148170 327374 148226
rect 327430 148170 327498 148226
rect 327554 148170 327622 148226
rect 327678 148170 327774 148226
rect 327154 148102 327774 148170
rect 327154 148046 327250 148102
rect 327306 148046 327374 148102
rect 327430 148046 327498 148102
rect 327554 148046 327622 148102
rect 327678 148046 327774 148102
rect 327154 147978 327774 148046
rect 327154 147922 327250 147978
rect 327306 147922 327374 147978
rect 327430 147922 327498 147978
rect 327554 147922 327622 147978
rect 327678 147922 327774 147978
rect 327154 130350 327774 147922
rect 327154 130294 327250 130350
rect 327306 130294 327374 130350
rect 327430 130294 327498 130350
rect 327554 130294 327622 130350
rect 327678 130294 327774 130350
rect 327154 130226 327774 130294
rect 327154 130170 327250 130226
rect 327306 130170 327374 130226
rect 327430 130170 327498 130226
rect 327554 130170 327622 130226
rect 327678 130170 327774 130226
rect 327154 130102 327774 130170
rect 327154 130046 327250 130102
rect 327306 130046 327374 130102
rect 327430 130046 327498 130102
rect 327554 130046 327622 130102
rect 327678 130046 327774 130102
rect 327154 129978 327774 130046
rect 327154 129922 327250 129978
rect 327306 129922 327374 129978
rect 327430 129922 327498 129978
rect 327554 129922 327622 129978
rect 327678 129922 327774 129978
rect 327154 112350 327774 129922
rect 327154 112294 327250 112350
rect 327306 112294 327374 112350
rect 327430 112294 327498 112350
rect 327554 112294 327622 112350
rect 327678 112294 327774 112350
rect 327154 112226 327774 112294
rect 327154 112170 327250 112226
rect 327306 112170 327374 112226
rect 327430 112170 327498 112226
rect 327554 112170 327622 112226
rect 327678 112170 327774 112226
rect 327154 112102 327774 112170
rect 327154 112046 327250 112102
rect 327306 112046 327374 112102
rect 327430 112046 327498 112102
rect 327554 112046 327622 112102
rect 327678 112046 327774 112102
rect 327154 111978 327774 112046
rect 327154 111922 327250 111978
rect 327306 111922 327374 111978
rect 327430 111922 327498 111978
rect 327554 111922 327622 111978
rect 327678 111922 327774 111978
rect 327154 94350 327774 111922
rect 327154 94294 327250 94350
rect 327306 94294 327374 94350
rect 327430 94294 327498 94350
rect 327554 94294 327622 94350
rect 327678 94294 327774 94350
rect 327154 94226 327774 94294
rect 327154 94170 327250 94226
rect 327306 94170 327374 94226
rect 327430 94170 327498 94226
rect 327554 94170 327622 94226
rect 327678 94170 327774 94226
rect 327154 94102 327774 94170
rect 327154 94046 327250 94102
rect 327306 94046 327374 94102
rect 327430 94046 327498 94102
rect 327554 94046 327622 94102
rect 327678 94046 327774 94102
rect 327154 93978 327774 94046
rect 327154 93922 327250 93978
rect 327306 93922 327374 93978
rect 327430 93922 327498 93978
rect 327554 93922 327622 93978
rect 327678 93922 327774 93978
rect 327154 76350 327774 93922
rect 327154 76294 327250 76350
rect 327306 76294 327374 76350
rect 327430 76294 327498 76350
rect 327554 76294 327622 76350
rect 327678 76294 327774 76350
rect 327154 76226 327774 76294
rect 327154 76170 327250 76226
rect 327306 76170 327374 76226
rect 327430 76170 327498 76226
rect 327554 76170 327622 76226
rect 327678 76170 327774 76226
rect 327154 76102 327774 76170
rect 327154 76046 327250 76102
rect 327306 76046 327374 76102
rect 327430 76046 327498 76102
rect 327554 76046 327622 76102
rect 327678 76046 327774 76102
rect 327154 75978 327774 76046
rect 327154 75922 327250 75978
rect 327306 75922 327374 75978
rect 327430 75922 327498 75978
rect 327554 75922 327622 75978
rect 327678 75922 327774 75978
rect 327154 58350 327774 75922
rect 327154 58294 327250 58350
rect 327306 58294 327374 58350
rect 327430 58294 327498 58350
rect 327554 58294 327622 58350
rect 327678 58294 327774 58350
rect 327154 58226 327774 58294
rect 327154 58170 327250 58226
rect 327306 58170 327374 58226
rect 327430 58170 327498 58226
rect 327554 58170 327622 58226
rect 327678 58170 327774 58226
rect 327154 58102 327774 58170
rect 327154 58046 327250 58102
rect 327306 58046 327374 58102
rect 327430 58046 327498 58102
rect 327554 58046 327622 58102
rect 327678 58046 327774 58102
rect 327154 57978 327774 58046
rect 327154 57922 327250 57978
rect 327306 57922 327374 57978
rect 327430 57922 327498 57978
rect 327554 57922 327622 57978
rect 327678 57922 327774 57978
rect 327154 40350 327774 57922
rect 327154 40294 327250 40350
rect 327306 40294 327374 40350
rect 327430 40294 327498 40350
rect 327554 40294 327622 40350
rect 327678 40294 327774 40350
rect 327154 40226 327774 40294
rect 327154 40170 327250 40226
rect 327306 40170 327374 40226
rect 327430 40170 327498 40226
rect 327554 40170 327622 40226
rect 327678 40170 327774 40226
rect 327154 40102 327774 40170
rect 327154 40046 327250 40102
rect 327306 40046 327374 40102
rect 327430 40046 327498 40102
rect 327554 40046 327622 40102
rect 327678 40046 327774 40102
rect 327154 39978 327774 40046
rect 327154 39922 327250 39978
rect 327306 39922 327374 39978
rect 327430 39922 327498 39978
rect 327554 39922 327622 39978
rect 327678 39922 327774 39978
rect 327154 22350 327774 39922
rect 327154 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 327774 22350
rect 327154 22226 327774 22294
rect 327154 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 327774 22226
rect 327154 22102 327774 22170
rect 327154 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 327774 22102
rect 327154 21978 327774 22046
rect 327154 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 327774 21978
rect 327154 4350 327774 21922
rect 327154 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 327774 4350
rect 327154 4226 327774 4294
rect 327154 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 327774 4226
rect 327154 4102 327774 4170
rect 327154 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 327774 4102
rect 327154 3978 327774 4046
rect 327154 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 327774 3978
rect 327154 -160 327774 3922
rect 327154 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 327774 -160
rect 327154 -284 327774 -216
rect 327154 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 327774 -284
rect 327154 -408 327774 -340
rect 327154 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 327774 -408
rect 327154 -532 327774 -464
rect 327154 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 327774 -532
rect 327154 -1644 327774 -588
rect 330874 190350 331494 207922
rect 342688 208350 343008 208384
rect 342688 208294 342758 208350
rect 342814 208294 342882 208350
rect 342938 208294 343008 208350
rect 342688 208226 343008 208294
rect 342688 208170 342758 208226
rect 342814 208170 342882 208226
rect 342938 208170 343008 208226
rect 342688 208102 343008 208170
rect 342688 208046 342758 208102
rect 342814 208046 342882 208102
rect 342938 208046 343008 208102
rect 342688 207978 343008 208046
rect 342688 207922 342758 207978
rect 342814 207922 342882 207978
rect 342938 207922 343008 207978
rect 342688 207888 343008 207922
rect 330874 190294 330970 190350
rect 331026 190294 331094 190350
rect 331150 190294 331218 190350
rect 331274 190294 331342 190350
rect 331398 190294 331494 190350
rect 330874 190226 331494 190294
rect 330874 190170 330970 190226
rect 331026 190170 331094 190226
rect 331150 190170 331218 190226
rect 331274 190170 331342 190226
rect 331398 190170 331494 190226
rect 330874 190102 331494 190170
rect 330874 190046 330970 190102
rect 331026 190046 331094 190102
rect 331150 190046 331218 190102
rect 331274 190046 331342 190102
rect 331398 190046 331494 190102
rect 330874 189978 331494 190046
rect 330874 189922 330970 189978
rect 331026 189922 331094 189978
rect 331150 189922 331218 189978
rect 331274 189922 331342 189978
rect 331398 189922 331494 189978
rect 330874 172350 331494 189922
rect 330874 172294 330970 172350
rect 331026 172294 331094 172350
rect 331150 172294 331218 172350
rect 331274 172294 331342 172350
rect 331398 172294 331494 172350
rect 330874 172226 331494 172294
rect 330874 172170 330970 172226
rect 331026 172170 331094 172226
rect 331150 172170 331218 172226
rect 331274 172170 331342 172226
rect 331398 172170 331494 172226
rect 330874 172102 331494 172170
rect 330874 172046 330970 172102
rect 331026 172046 331094 172102
rect 331150 172046 331218 172102
rect 331274 172046 331342 172102
rect 331398 172046 331494 172102
rect 330874 171978 331494 172046
rect 330874 171922 330970 171978
rect 331026 171922 331094 171978
rect 331150 171922 331218 171978
rect 331274 171922 331342 171978
rect 331398 171922 331494 171978
rect 330874 154350 331494 171922
rect 330874 154294 330970 154350
rect 331026 154294 331094 154350
rect 331150 154294 331218 154350
rect 331274 154294 331342 154350
rect 331398 154294 331494 154350
rect 330874 154226 331494 154294
rect 330874 154170 330970 154226
rect 331026 154170 331094 154226
rect 331150 154170 331218 154226
rect 331274 154170 331342 154226
rect 331398 154170 331494 154226
rect 330874 154102 331494 154170
rect 330874 154046 330970 154102
rect 331026 154046 331094 154102
rect 331150 154046 331218 154102
rect 331274 154046 331342 154102
rect 331398 154046 331494 154102
rect 330874 153978 331494 154046
rect 330874 153922 330970 153978
rect 331026 153922 331094 153978
rect 331150 153922 331218 153978
rect 331274 153922 331342 153978
rect 331398 153922 331494 153978
rect 330874 136350 331494 153922
rect 330874 136294 330970 136350
rect 331026 136294 331094 136350
rect 331150 136294 331218 136350
rect 331274 136294 331342 136350
rect 331398 136294 331494 136350
rect 330874 136226 331494 136294
rect 330874 136170 330970 136226
rect 331026 136170 331094 136226
rect 331150 136170 331218 136226
rect 331274 136170 331342 136226
rect 331398 136170 331494 136226
rect 330874 136102 331494 136170
rect 330874 136046 330970 136102
rect 331026 136046 331094 136102
rect 331150 136046 331218 136102
rect 331274 136046 331342 136102
rect 331398 136046 331494 136102
rect 330874 135978 331494 136046
rect 330874 135922 330970 135978
rect 331026 135922 331094 135978
rect 331150 135922 331218 135978
rect 331274 135922 331342 135978
rect 331398 135922 331494 135978
rect 330874 118350 331494 135922
rect 330874 118294 330970 118350
rect 331026 118294 331094 118350
rect 331150 118294 331218 118350
rect 331274 118294 331342 118350
rect 331398 118294 331494 118350
rect 330874 118226 331494 118294
rect 330874 118170 330970 118226
rect 331026 118170 331094 118226
rect 331150 118170 331218 118226
rect 331274 118170 331342 118226
rect 331398 118170 331494 118226
rect 330874 118102 331494 118170
rect 330874 118046 330970 118102
rect 331026 118046 331094 118102
rect 331150 118046 331218 118102
rect 331274 118046 331342 118102
rect 331398 118046 331494 118102
rect 330874 117978 331494 118046
rect 330874 117922 330970 117978
rect 331026 117922 331094 117978
rect 331150 117922 331218 117978
rect 331274 117922 331342 117978
rect 331398 117922 331494 117978
rect 330874 100350 331494 117922
rect 330874 100294 330970 100350
rect 331026 100294 331094 100350
rect 331150 100294 331218 100350
rect 331274 100294 331342 100350
rect 331398 100294 331494 100350
rect 330874 100226 331494 100294
rect 330874 100170 330970 100226
rect 331026 100170 331094 100226
rect 331150 100170 331218 100226
rect 331274 100170 331342 100226
rect 331398 100170 331494 100226
rect 330874 100102 331494 100170
rect 330874 100046 330970 100102
rect 331026 100046 331094 100102
rect 331150 100046 331218 100102
rect 331274 100046 331342 100102
rect 331398 100046 331494 100102
rect 330874 99978 331494 100046
rect 330874 99922 330970 99978
rect 331026 99922 331094 99978
rect 331150 99922 331218 99978
rect 331274 99922 331342 99978
rect 331398 99922 331494 99978
rect 330874 82350 331494 99922
rect 330874 82294 330970 82350
rect 331026 82294 331094 82350
rect 331150 82294 331218 82350
rect 331274 82294 331342 82350
rect 331398 82294 331494 82350
rect 330874 82226 331494 82294
rect 330874 82170 330970 82226
rect 331026 82170 331094 82226
rect 331150 82170 331218 82226
rect 331274 82170 331342 82226
rect 331398 82170 331494 82226
rect 330874 82102 331494 82170
rect 330874 82046 330970 82102
rect 331026 82046 331094 82102
rect 331150 82046 331218 82102
rect 331274 82046 331342 82102
rect 331398 82046 331494 82102
rect 330874 81978 331494 82046
rect 330874 81922 330970 81978
rect 331026 81922 331094 81978
rect 331150 81922 331218 81978
rect 331274 81922 331342 81978
rect 331398 81922 331494 81978
rect 330874 64350 331494 81922
rect 330874 64294 330970 64350
rect 331026 64294 331094 64350
rect 331150 64294 331218 64350
rect 331274 64294 331342 64350
rect 331398 64294 331494 64350
rect 330874 64226 331494 64294
rect 330874 64170 330970 64226
rect 331026 64170 331094 64226
rect 331150 64170 331218 64226
rect 331274 64170 331342 64226
rect 331398 64170 331494 64226
rect 330874 64102 331494 64170
rect 330874 64046 330970 64102
rect 331026 64046 331094 64102
rect 331150 64046 331218 64102
rect 331274 64046 331342 64102
rect 331398 64046 331494 64102
rect 330874 63978 331494 64046
rect 330874 63922 330970 63978
rect 331026 63922 331094 63978
rect 331150 63922 331218 63978
rect 331274 63922 331342 63978
rect 331398 63922 331494 63978
rect 330874 46350 331494 63922
rect 330874 46294 330970 46350
rect 331026 46294 331094 46350
rect 331150 46294 331218 46350
rect 331274 46294 331342 46350
rect 331398 46294 331494 46350
rect 330874 46226 331494 46294
rect 330874 46170 330970 46226
rect 331026 46170 331094 46226
rect 331150 46170 331218 46226
rect 331274 46170 331342 46226
rect 331398 46170 331494 46226
rect 330874 46102 331494 46170
rect 330874 46046 330970 46102
rect 331026 46046 331094 46102
rect 331150 46046 331218 46102
rect 331274 46046 331342 46102
rect 331398 46046 331494 46102
rect 330874 45978 331494 46046
rect 330874 45922 330970 45978
rect 331026 45922 331094 45978
rect 331150 45922 331218 45978
rect 331274 45922 331342 45978
rect 331398 45922 331494 45978
rect 330874 28350 331494 45922
rect 330874 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 331494 28350
rect 330874 28226 331494 28294
rect 330874 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 331494 28226
rect 330874 28102 331494 28170
rect 330874 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 331494 28102
rect 330874 27978 331494 28046
rect 330874 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 331494 27978
rect 330874 10350 331494 27922
rect 330874 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 331494 10350
rect 330874 10226 331494 10294
rect 330874 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 331494 10226
rect 330874 10102 331494 10170
rect 330874 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 331494 10102
rect 330874 9978 331494 10046
rect 330874 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 331494 9978
rect 330874 -1120 331494 9922
rect 330874 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 331494 -1120
rect 330874 -1244 331494 -1176
rect 330874 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 331494 -1244
rect 330874 -1368 331494 -1300
rect 330874 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 331494 -1368
rect 330874 -1492 331494 -1424
rect 330874 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 331494 -1492
rect 330874 -1644 331494 -1548
rect 345154 202350 345774 210842
rect 345154 202294 345250 202350
rect 345306 202294 345374 202350
rect 345430 202294 345498 202350
rect 345554 202294 345622 202350
rect 345678 202294 345774 202350
rect 345154 202226 345774 202294
rect 345154 202170 345250 202226
rect 345306 202170 345374 202226
rect 345430 202170 345498 202226
rect 345554 202170 345622 202226
rect 345678 202170 345774 202226
rect 345154 202102 345774 202170
rect 345154 202046 345250 202102
rect 345306 202046 345374 202102
rect 345430 202046 345498 202102
rect 345554 202046 345622 202102
rect 345678 202046 345774 202102
rect 345154 201978 345774 202046
rect 345154 201922 345250 201978
rect 345306 201922 345374 201978
rect 345430 201922 345498 201978
rect 345554 201922 345622 201978
rect 345678 201922 345774 201978
rect 345154 184350 345774 201922
rect 345154 184294 345250 184350
rect 345306 184294 345374 184350
rect 345430 184294 345498 184350
rect 345554 184294 345622 184350
rect 345678 184294 345774 184350
rect 345154 184226 345774 184294
rect 345154 184170 345250 184226
rect 345306 184170 345374 184226
rect 345430 184170 345498 184226
rect 345554 184170 345622 184226
rect 345678 184170 345774 184226
rect 345154 184102 345774 184170
rect 345154 184046 345250 184102
rect 345306 184046 345374 184102
rect 345430 184046 345498 184102
rect 345554 184046 345622 184102
rect 345678 184046 345774 184102
rect 345154 183978 345774 184046
rect 345154 183922 345250 183978
rect 345306 183922 345374 183978
rect 345430 183922 345498 183978
rect 345554 183922 345622 183978
rect 345678 183922 345774 183978
rect 345154 166350 345774 183922
rect 345154 166294 345250 166350
rect 345306 166294 345374 166350
rect 345430 166294 345498 166350
rect 345554 166294 345622 166350
rect 345678 166294 345774 166350
rect 345154 166226 345774 166294
rect 345154 166170 345250 166226
rect 345306 166170 345374 166226
rect 345430 166170 345498 166226
rect 345554 166170 345622 166226
rect 345678 166170 345774 166226
rect 345154 166102 345774 166170
rect 345154 166046 345250 166102
rect 345306 166046 345374 166102
rect 345430 166046 345498 166102
rect 345554 166046 345622 166102
rect 345678 166046 345774 166102
rect 345154 165978 345774 166046
rect 345154 165922 345250 165978
rect 345306 165922 345374 165978
rect 345430 165922 345498 165978
rect 345554 165922 345622 165978
rect 345678 165922 345774 165978
rect 345154 148350 345774 165922
rect 345154 148294 345250 148350
rect 345306 148294 345374 148350
rect 345430 148294 345498 148350
rect 345554 148294 345622 148350
rect 345678 148294 345774 148350
rect 345154 148226 345774 148294
rect 345154 148170 345250 148226
rect 345306 148170 345374 148226
rect 345430 148170 345498 148226
rect 345554 148170 345622 148226
rect 345678 148170 345774 148226
rect 345154 148102 345774 148170
rect 345154 148046 345250 148102
rect 345306 148046 345374 148102
rect 345430 148046 345498 148102
rect 345554 148046 345622 148102
rect 345678 148046 345774 148102
rect 345154 147978 345774 148046
rect 345154 147922 345250 147978
rect 345306 147922 345374 147978
rect 345430 147922 345498 147978
rect 345554 147922 345622 147978
rect 345678 147922 345774 147978
rect 345154 130350 345774 147922
rect 345154 130294 345250 130350
rect 345306 130294 345374 130350
rect 345430 130294 345498 130350
rect 345554 130294 345622 130350
rect 345678 130294 345774 130350
rect 345154 130226 345774 130294
rect 345154 130170 345250 130226
rect 345306 130170 345374 130226
rect 345430 130170 345498 130226
rect 345554 130170 345622 130226
rect 345678 130170 345774 130226
rect 345154 130102 345774 130170
rect 345154 130046 345250 130102
rect 345306 130046 345374 130102
rect 345430 130046 345498 130102
rect 345554 130046 345622 130102
rect 345678 130046 345774 130102
rect 345154 129978 345774 130046
rect 345154 129922 345250 129978
rect 345306 129922 345374 129978
rect 345430 129922 345498 129978
rect 345554 129922 345622 129978
rect 345678 129922 345774 129978
rect 345154 112350 345774 129922
rect 345154 112294 345250 112350
rect 345306 112294 345374 112350
rect 345430 112294 345498 112350
rect 345554 112294 345622 112350
rect 345678 112294 345774 112350
rect 345154 112226 345774 112294
rect 345154 112170 345250 112226
rect 345306 112170 345374 112226
rect 345430 112170 345498 112226
rect 345554 112170 345622 112226
rect 345678 112170 345774 112226
rect 345154 112102 345774 112170
rect 345154 112046 345250 112102
rect 345306 112046 345374 112102
rect 345430 112046 345498 112102
rect 345554 112046 345622 112102
rect 345678 112046 345774 112102
rect 345154 111978 345774 112046
rect 345154 111922 345250 111978
rect 345306 111922 345374 111978
rect 345430 111922 345498 111978
rect 345554 111922 345622 111978
rect 345678 111922 345774 111978
rect 345154 94350 345774 111922
rect 345154 94294 345250 94350
rect 345306 94294 345374 94350
rect 345430 94294 345498 94350
rect 345554 94294 345622 94350
rect 345678 94294 345774 94350
rect 345154 94226 345774 94294
rect 345154 94170 345250 94226
rect 345306 94170 345374 94226
rect 345430 94170 345498 94226
rect 345554 94170 345622 94226
rect 345678 94170 345774 94226
rect 345154 94102 345774 94170
rect 345154 94046 345250 94102
rect 345306 94046 345374 94102
rect 345430 94046 345498 94102
rect 345554 94046 345622 94102
rect 345678 94046 345774 94102
rect 345154 93978 345774 94046
rect 345154 93922 345250 93978
rect 345306 93922 345374 93978
rect 345430 93922 345498 93978
rect 345554 93922 345622 93978
rect 345678 93922 345774 93978
rect 345154 76350 345774 93922
rect 345154 76294 345250 76350
rect 345306 76294 345374 76350
rect 345430 76294 345498 76350
rect 345554 76294 345622 76350
rect 345678 76294 345774 76350
rect 345154 76226 345774 76294
rect 345154 76170 345250 76226
rect 345306 76170 345374 76226
rect 345430 76170 345498 76226
rect 345554 76170 345622 76226
rect 345678 76170 345774 76226
rect 345154 76102 345774 76170
rect 345154 76046 345250 76102
rect 345306 76046 345374 76102
rect 345430 76046 345498 76102
rect 345554 76046 345622 76102
rect 345678 76046 345774 76102
rect 345154 75978 345774 76046
rect 345154 75922 345250 75978
rect 345306 75922 345374 75978
rect 345430 75922 345498 75978
rect 345554 75922 345622 75978
rect 345678 75922 345774 75978
rect 345154 58350 345774 75922
rect 345154 58294 345250 58350
rect 345306 58294 345374 58350
rect 345430 58294 345498 58350
rect 345554 58294 345622 58350
rect 345678 58294 345774 58350
rect 345154 58226 345774 58294
rect 345154 58170 345250 58226
rect 345306 58170 345374 58226
rect 345430 58170 345498 58226
rect 345554 58170 345622 58226
rect 345678 58170 345774 58226
rect 345154 58102 345774 58170
rect 345154 58046 345250 58102
rect 345306 58046 345374 58102
rect 345430 58046 345498 58102
rect 345554 58046 345622 58102
rect 345678 58046 345774 58102
rect 345154 57978 345774 58046
rect 345154 57922 345250 57978
rect 345306 57922 345374 57978
rect 345430 57922 345498 57978
rect 345554 57922 345622 57978
rect 345678 57922 345774 57978
rect 345154 40350 345774 57922
rect 345154 40294 345250 40350
rect 345306 40294 345374 40350
rect 345430 40294 345498 40350
rect 345554 40294 345622 40350
rect 345678 40294 345774 40350
rect 345154 40226 345774 40294
rect 345154 40170 345250 40226
rect 345306 40170 345374 40226
rect 345430 40170 345498 40226
rect 345554 40170 345622 40226
rect 345678 40170 345774 40226
rect 345154 40102 345774 40170
rect 345154 40046 345250 40102
rect 345306 40046 345374 40102
rect 345430 40046 345498 40102
rect 345554 40046 345622 40102
rect 345678 40046 345774 40102
rect 345154 39978 345774 40046
rect 345154 39922 345250 39978
rect 345306 39922 345374 39978
rect 345430 39922 345498 39978
rect 345554 39922 345622 39978
rect 345678 39922 345774 39978
rect 345154 22350 345774 39922
rect 345154 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 345774 22350
rect 345154 22226 345774 22294
rect 345154 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 345774 22226
rect 345154 22102 345774 22170
rect 345154 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 345774 22102
rect 345154 21978 345774 22046
rect 345154 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 345774 21978
rect 345154 4350 345774 21922
rect 345154 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 345774 4350
rect 345154 4226 345774 4294
rect 345154 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 345774 4226
rect 345154 4102 345774 4170
rect 345154 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 345774 4102
rect 345154 3978 345774 4046
rect 345154 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 345774 3978
rect 345154 -160 345774 3922
rect 345154 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 345774 -160
rect 345154 -284 345774 -216
rect 345154 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 345774 -284
rect 345154 -408 345774 -340
rect 345154 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 345774 -408
rect 345154 -532 345774 -464
rect 345154 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 345774 -532
rect 345154 -1644 345774 -588
rect 348874 208350 349494 210842
rect 348874 208294 348970 208350
rect 349026 208294 349094 208350
rect 349150 208294 349218 208350
rect 349274 208294 349342 208350
rect 349398 208294 349494 208350
rect 348874 208226 349494 208294
rect 348874 208170 348970 208226
rect 349026 208170 349094 208226
rect 349150 208170 349218 208226
rect 349274 208170 349342 208226
rect 349398 208170 349494 208226
rect 348874 208102 349494 208170
rect 348874 208046 348970 208102
rect 349026 208046 349094 208102
rect 349150 208046 349218 208102
rect 349274 208046 349342 208102
rect 349398 208046 349494 208102
rect 348874 207978 349494 208046
rect 348874 207922 348970 207978
rect 349026 207922 349094 207978
rect 349150 207922 349218 207978
rect 349274 207922 349342 207978
rect 349398 207922 349494 207978
rect 348874 190350 349494 207922
rect 348874 190294 348970 190350
rect 349026 190294 349094 190350
rect 349150 190294 349218 190350
rect 349274 190294 349342 190350
rect 349398 190294 349494 190350
rect 348874 190226 349494 190294
rect 348874 190170 348970 190226
rect 349026 190170 349094 190226
rect 349150 190170 349218 190226
rect 349274 190170 349342 190226
rect 349398 190170 349494 190226
rect 348874 190102 349494 190170
rect 348874 190046 348970 190102
rect 349026 190046 349094 190102
rect 349150 190046 349218 190102
rect 349274 190046 349342 190102
rect 349398 190046 349494 190102
rect 348874 189978 349494 190046
rect 348874 189922 348970 189978
rect 349026 189922 349094 189978
rect 349150 189922 349218 189978
rect 349274 189922 349342 189978
rect 349398 189922 349494 189978
rect 348874 172350 349494 189922
rect 348874 172294 348970 172350
rect 349026 172294 349094 172350
rect 349150 172294 349218 172350
rect 349274 172294 349342 172350
rect 349398 172294 349494 172350
rect 348874 172226 349494 172294
rect 348874 172170 348970 172226
rect 349026 172170 349094 172226
rect 349150 172170 349218 172226
rect 349274 172170 349342 172226
rect 349398 172170 349494 172226
rect 348874 172102 349494 172170
rect 348874 172046 348970 172102
rect 349026 172046 349094 172102
rect 349150 172046 349218 172102
rect 349274 172046 349342 172102
rect 349398 172046 349494 172102
rect 348874 171978 349494 172046
rect 348874 171922 348970 171978
rect 349026 171922 349094 171978
rect 349150 171922 349218 171978
rect 349274 171922 349342 171978
rect 349398 171922 349494 171978
rect 348874 154350 349494 171922
rect 348874 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 349494 154350
rect 348874 154226 349494 154294
rect 348874 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 349494 154226
rect 348874 154102 349494 154170
rect 348874 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 349494 154102
rect 348874 153978 349494 154046
rect 348874 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 349494 153978
rect 348874 136350 349494 153922
rect 348874 136294 348970 136350
rect 349026 136294 349094 136350
rect 349150 136294 349218 136350
rect 349274 136294 349342 136350
rect 349398 136294 349494 136350
rect 348874 136226 349494 136294
rect 348874 136170 348970 136226
rect 349026 136170 349094 136226
rect 349150 136170 349218 136226
rect 349274 136170 349342 136226
rect 349398 136170 349494 136226
rect 348874 136102 349494 136170
rect 348874 136046 348970 136102
rect 349026 136046 349094 136102
rect 349150 136046 349218 136102
rect 349274 136046 349342 136102
rect 349398 136046 349494 136102
rect 348874 135978 349494 136046
rect 348874 135922 348970 135978
rect 349026 135922 349094 135978
rect 349150 135922 349218 135978
rect 349274 135922 349342 135978
rect 349398 135922 349494 135978
rect 348874 118350 349494 135922
rect 348874 118294 348970 118350
rect 349026 118294 349094 118350
rect 349150 118294 349218 118350
rect 349274 118294 349342 118350
rect 349398 118294 349494 118350
rect 348874 118226 349494 118294
rect 348874 118170 348970 118226
rect 349026 118170 349094 118226
rect 349150 118170 349218 118226
rect 349274 118170 349342 118226
rect 349398 118170 349494 118226
rect 348874 118102 349494 118170
rect 348874 118046 348970 118102
rect 349026 118046 349094 118102
rect 349150 118046 349218 118102
rect 349274 118046 349342 118102
rect 349398 118046 349494 118102
rect 348874 117978 349494 118046
rect 348874 117922 348970 117978
rect 349026 117922 349094 117978
rect 349150 117922 349218 117978
rect 349274 117922 349342 117978
rect 349398 117922 349494 117978
rect 348874 100350 349494 117922
rect 348874 100294 348970 100350
rect 349026 100294 349094 100350
rect 349150 100294 349218 100350
rect 349274 100294 349342 100350
rect 349398 100294 349494 100350
rect 348874 100226 349494 100294
rect 348874 100170 348970 100226
rect 349026 100170 349094 100226
rect 349150 100170 349218 100226
rect 349274 100170 349342 100226
rect 349398 100170 349494 100226
rect 348874 100102 349494 100170
rect 348874 100046 348970 100102
rect 349026 100046 349094 100102
rect 349150 100046 349218 100102
rect 349274 100046 349342 100102
rect 349398 100046 349494 100102
rect 348874 99978 349494 100046
rect 348874 99922 348970 99978
rect 349026 99922 349094 99978
rect 349150 99922 349218 99978
rect 349274 99922 349342 99978
rect 349398 99922 349494 99978
rect 348874 82350 349494 99922
rect 348874 82294 348970 82350
rect 349026 82294 349094 82350
rect 349150 82294 349218 82350
rect 349274 82294 349342 82350
rect 349398 82294 349494 82350
rect 348874 82226 349494 82294
rect 348874 82170 348970 82226
rect 349026 82170 349094 82226
rect 349150 82170 349218 82226
rect 349274 82170 349342 82226
rect 349398 82170 349494 82226
rect 348874 82102 349494 82170
rect 348874 82046 348970 82102
rect 349026 82046 349094 82102
rect 349150 82046 349218 82102
rect 349274 82046 349342 82102
rect 349398 82046 349494 82102
rect 348874 81978 349494 82046
rect 348874 81922 348970 81978
rect 349026 81922 349094 81978
rect 349150 81922 349218 81978
rect 349274 81922 349342 81978
rect 349398 81922 349494 81978
rect 348874 64350 349494 81922
rect 348874 64294 348970 64350
rect 349026 64294 349094 64350
rect 349150 64294 349218 64350
rect 349274 64294 349342 64350
rect 349398 64294 349494 64350
rect 348874 64226 349494 64294
rect 348874 64170 348970 64226
rect 349026 64170 349094 64226
rect 349150 64170 349218 64226
rect 349274 64170 349342 64226
rect 349398 64170 349494 64226
rect 348874 64102 349494 64170
rect 348874 64046 348970 64102
rect 349026 64046 349094 64102
rect 349150 64046 349218 64102
rect 349274 64046 349342 64102
rect 349398 64046 349494 64102
rect 348874 63978 349494 64046
rect 348874 63922 348970 63978
rect 349026 63922 349094 63978
rect 349150 63922 349218 63978
rect 349274 63922 349342 63978
rect 349398 63922 349494 63978
rect 348874 46350 349494 63922
rect 348874 46294 348970 46350
rect 349026 46294 349094 46350
rect 349150 46294 349218 46350
rect 349274 46294 349342 46350
rect 349398 46294 349494 46350
rect 348874 46226 349494 46294
rect 348874 46170 348970 46226
rect 349026 46170 349094 46226
rect 349150 46170 349218 46226
rect 349274 46170 349342 46226
rect 349398 46170 349494 46226
rect 348874 46102 349494 46170
rect 348874 46046 348970 46102
rect 349026 46046 349094 46102
rect 349150 46046 349218 46102
rect 349274 46046 349342 46102
rect 349398 46046 349494 46102
rect 348874 45978 349494 46046
rect 348874 45922 348970 45978
rect 349026 45922 349094 45978
rect 349150 45922 349218 45978
rect 349274 45922 349342 45978
rect 349398 45922 349494 45978
rect 348874 28350 349494 45922
rect 348874 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 349494 28350
rect 348874 28226 349494 28294
rect 348874 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 349494 28226
rect 348874 28102 349494 28170
rect 348874 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 349494 28102
rect 348874 27978 349494 28046
rect 348874 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 349494 27978
rect 348874 10350 349494 27922
rect 348874 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 349494 10350
rect 348874 10226 349494 10294
rect 348874 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 349494 10226
rect 348874 10102 349494 10170
rect 348874 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 349494 10102
rect 348874 9978 349494 10046
rect 348874 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 349494 9978
rect 348874 -1120 349494 9922
rect 348874 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 349494 -1120
rect 348874 -1244 349494 -1176
rect 348874 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 349494 -1244
rect 348874 -1368 349494 -1300
rect 348874 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 349494 -1368
rect 348874 -1492 349494 -1424
rect 348874 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 349494 -1492
rect 348874 -1644 349494 -1548
rect 363154 202350 363774 210842
rect 363154 202294 363250 202350
rect 363306 202294 363374 202350
rect 363430 202294 363498 202350
rect 363554 202294 363622 202350
rect 363678 202294 363774 202350
rect 363154 202226 363774 202294
rect 363154 202170 363250 202226
rect 363306 202170 363374 202226
rect 363430 202170 363498 202226
rect 363554 202170 363622 202226
rect 363678 202170 363774 202226
rect 363154 202102 363774 202170
rect 363154 202046 363250 202102
rect 363306 202046 363374 202102
rect 363430 202046 363498 202102
rect 363554 202046 363622 202102
rect 363678 202046 363774 202102
rect 363154 201978 363774 202046
rect 363154 201922 363250 201978
rect 363306 201922 363374 201978
rect 363430 201922 363498 201978
rect 363554 201922 363622 201978
rect 363678 201922 363774 201978
rect 363154 184350 363774 201922
rect 363154 184294 363250 184350
rect 363306 184294 363374 184350
rect 363430 184294 363498 184350
rect 363554 184294 363622 184350
rect 363678 184294 363774 184350
rect 363154 184226 363774 184294
rect 363154 184170 363250 184226
rect 363306 184170 363374 184226
rect 363430 184170 363498 184226
rect 363554 184170 363622 184226
rect 363678 184170 363774 184226
rect 363154 184102 363774 184170
rect 363154 184046 363250 184102
rect 363306 184046 363374 184102
rect 363430 184046 363498 184102
rect 363554 184046 363622 184102
rect 363678 184046 363774 184102
rect 363154 183978 363774 184046
rect 363154 183922 363250 183978
rect 363306 183922 363374 183978
rect 363430 183922 363498 183978
rect 363554 183922 363622 183978
rect 363678 183922 363774 183978
rect 363154 166350 363774 183922
rect 363154 166294 363250 166350
rect 363306 166294 363374 166350
rect 363430 166294 363498 166350
rect 363554 166294 363622 166350
rect 363678 166294 363774 166350
rect 363154 166226 363774 166294
rect 363154 166170 363250 166226
rect 363306 166170 363374 166226
rect 363430 166170 363498 166226
rect 363554 166170 363622 166226
rect 363678 166170 363774 166226
rect 363154 166102 363774 166170
rect 363154 166046 363250 166102
rect 363306 166046 363374 166102
rect 363430 166046 363498 166102
rect 363554 166046 363622 166102
rect 363678 166046 363774 166102
rect 363154 165978 363774 166046
rect 363154 165922 363250 165978
rect 363306 165922 363374 165978
rect 363430 165922 363498 165978
rect 363554 165922 363622 165978
rect 363678 165922 363774 165978
rect 363154 148350 363774 165922
rect 363154 148294 363250 148350
rect 363306 148294 363374 148350
rect 363430 148294 363498 148350
rect 363554 148294 363622 148350
rect 363678 148294 363774 148350
rect 363154 148226 363774 148294
rect 363154 148170 363250 148226
rect 363306 148170 363374 148226
rect 363430 148170 363498 148226
rect 363554 148170 363622 148226
rect 363678 148170 363774 148226
rect 363154 148102 363774 148170
rect 363154 148046 363250 148102
rect 363306 148046 363374 148102
rect 363430 148046 363498 148102
rect 363554 148046 363622 148102
rect 363678 148046 363774 148102
rect 363154 147978 363774 148046
rect 363154 147922 363250 147978
rect 363306 147922 363374 147978
rect 363430 147922 363498 147978
rect 363554 147922 363622 147978
rect 363678 147922 363774 147978
rect 363154 130350 363774 147922
rect 363154 130294 363250 130350
rect 363306 130294 363374 130350
rect 363430 130294 363498 130350
rect 363554 130294 363622 130350
rect 363678 130294 363774 130350
rect 363154 130226 363774 130294
rect 363154 130170 363250 130226
rect 363306 130170 363374 130226
rect 363430 130170 363498 130226
rect 363554 130170 363622 130226
rect 363678 130170 363774 130226
rect 363154 130102 363774 130170
rect 363154 130046 363250 130102
rect 363306 130046 363374 130102
rect 363430 130046 363498 130102
rect 363554 130046 363622 130102
rect 363678 130046 363774 130102
rect 363154 129978 363774 130046
rect 363154 129922 363250 129978
rect 363306 129922 363374 129978
rect 363430 129922 363498 129978
rect 363554 129922 363622 129978
rect 363678 129922 363774 129978
rect 363154 112350 363774 129922
rect 363154 112294 363250 112350
rect 363306 112294 363374 112350
rect 363430 112294 363498 112350
rect 363554 112294 363622 112350
rect 363678 112294 363774 112350
rect 363154 112226 363774 112294
rect 363154 112170 363250 112226
rect 363306 112170 363374 112226
rect 363430 112170 363498 112226
rect 363554 112170 363622 112226
rect 363678 112170 363774 112226
rect 363154 112102 363774 112170
rect 363154 112046 363250 112102
rect 363306 112046 363374 112102
rect 363430 112046 363498 112102
rect 363554 112046 363622 112102
rect 363678 112046 363774 112102
rect 363154 111978 363774 112046
rect 363154 111922 363250 111978
rect 363306 111922 363374 111978
rect 363430 111922 363498 111978
rect 363554 111922 363622 111978
rect 363678 111922 363774 111978
rect 363154 94350 363774 111922
rect 363154 94294 363250 94350
rect 363306 94294 363374 94350
rect 363430 94294 363498 94350
rect 363554 94294 363622 94350
rect 363678 94294 363774 94350
rect 363154 94226 363774 94294
rect 363154 94170 363250 94226
rect 363306 94170 363374 94226
rect 363430 94170 363498 94226
rect 363554 94170 363622 94226
rect 363678 94170 363774 94226
rect 363154 94102 363774 94170
rect 363154 94046 363250 94102
rect 363306 94046 363374 94102
rect 363430 94046 363498 94102
rect 363554 94046 363622 94102
rect 363678 94046 363774 94102
rect 363154 93978 363774 94046
rect 363154 93922 363250 93978
rect 363306 93922 363374 93978
rect 363430 93922 363498 93978
rect 363554 93922 363622 93978
rect 363678 93922 363774 93978
rect 363154 76350 363774 93922
rect 363154 76294 363250 76350
rect 363306 76294 363374 76350
rect 363430 76294 363498 76350
rect 363554 76294 363622 76350
rect 363678 76294 363774 76350
rect 363154 76226 363774 76294
rect 363154 76170 363250 76226
rect 363306 76170 363374 76226
rect 363430 76170 363498 76226
rect 363554 76170 363622 76226
rect 363678 76170 363774 76226
rect 363154 76102 363774 76170
rect 363154 76046 363250 76102
rect 363306 76046 363374 76102
rect 363430 76046 363498 76102
rect 363554 76046 363622 76102
rect 363678 76046 363774 76102
rect 363154 75978 363774 76046
rect 363154 75922 363250 75978
rect 363306 75922 363374 75978
rect 363430 75922 363498 75978
rect 363554 75922 363622 75978
rect 363678 75922 363774 75978
rect 363154 58350 363774 75922
rect 363154 58294 363250 58350
rect 363306 58294 363374 58350
rect 363430 58294 363498 58350
rect 363554 58294 363622 58350
rect 363678 58294 363774 58350
rect 363154 58226 363774 58294
rect 363154 58170 363250 58226
rect 363306 58170 363374 58226
rect 363430 58170 363498 58226
rect 363554 58170 363622 58226
rect 363678 58170 363774 58226
rect 363154 58102 363774 58170
rect 363154 58046 363250 58102
rect 363306 58046 363374 58102
rect 363430 58046 363498 58102
rect 363554 58046 363622 58102
rect 363678 58046 363774 58102
rect 363154 57978 363774 58046
rect 363154 57922 363250 57978
rect 363306 57922 363374 57978
rect 363430 57922 363498 57978
rect 363554 57922 363622 57978
rect 363678 57922 363774 57978
rect 363154 40350 363774 57922
rect 363154 40294 363250 40350
rect 363306 40294 363374 40350
rect 363430 40294 363498 40350
rect 363554 40294 363622 40350
rect 363678 40294 363774 40350
rect 363154 40226 363774 40294
rect 363154 40170 363250 40226
rect 363306 40170 363374 40226
rect 363430 40170 363498 40226
rect 363554 40170 363622 40226
rect 363678 40170 363774 40226
rect 363154 40102 363774 40170
rect 363154 40046 363250 40102
rect 363306 40046 363374 40102
rect 363430 40046 363498 40102
rect 363554 40046 363622 40102
rect 363678 40046 363774 40102
rect 363154 39978 363774 40046
rect 363154 39922 363250 39978
rect 363306 39922 363374 39978
rect 363430 39922 363498 39978
rect 363554 39922 363622 39978
rect 363678 39922 363774 39978
rect 363154 22350 363774 39922
rect 363154 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 363774 22350
rect 363154 22226 363774 22294
rect 363154 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 363774 22226
rect 363154 22102 363774 22170
rect 363154 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 363774 22102
rect 363154 21978 363774 22046
rect 363154 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 363774 21978
rect 363154 4350 363774 21922
rect 363154 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 363774 4350
rect 363154 4226 363774 4294
rect 363154 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 363774 4226
rect 363154 4102 363774 4170
rect 363154 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 363774 4102
rect 363154 3978 363774 4046
rect 363154 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 363774 3978
rect 363154 -160 363774 3922
rect 363154 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 363774 -160
rect 363154 -284 363774 -216
rect 363154 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 363774 -284
rect 363154 -408 363774 -340
rect 363154 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 363774 -408
rect 363154 -532 363774 -464
rect 363154 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 363774 -532
rect 363154 -1644 363774 -588
rect 366874 208350 367494 210842
rect 366874 208294 366970 208350
rect 367026 208294 367094 208350
rect 367150 208294 367218 208350
rect 367274 208294 367342 208350
rect 367398 208294 367494 208350
rect 366874 208226 367494 208294
rect 366874 208170 366970 208226
rect 367026 208170 367094 208226
rect 367150 208170 367218 208226
rect 367274 208170 367342 208226
rect 367398 208170 367494 208226
rect 366874 208102 367494 208170
rect 366874 208046 366970 208102
rect 367026 208046 367094 208102
rect 367150 208046 367218 208102
rect 367274 208046 367342 208102
rect 367398 208046 367494 208102
rect 366874 207978 367494 208046
rect 366874 207922 366970 207978
rect 367026 207922 367094 207978
rect 367150 207922 367218 207978
rect 367274 207922 367342 207978
rect 367398 207922 367494 207978
rect 366874 190350 367494 207922
rect 373408 208350 373728 208384
rect 373408 208294 373478 208350
rect 373534 208294 373602 208350
rect 373658 208294 373728 208350
rect 373408 208226 373728 208294
rect 373408 208170 373478 208226
rect 373534 208170 373602 208226
rect 373658 208170 373728 208226
rect 373408 208102 373728 208170
rect 373408 208046 373478 208102
rect 373534 208046 373602 208102
rect 373658 208046 373728 208102
rect 373408 207978 373728 208046
rect 373408 207922 373478 207978
rect 373534 207922 373602 207978
rect 373658 207922 373728 207978
rect 373408 207888 373728 207922
rect 366874 190294 366970 190350
rect 367026 190294 367094 190350
rect 367150 190294 367218 190350
rect 367274 190294 367342 190350
rect 367398 190294 367494 190350
rect 366874 190226 367494 190294
rect 366874 190170 366970 190226
rect 367026 190170 367094 190226
rect 367150 190170 367218 190226
rect 367274 190170 367342 190226
rect 367398 190170 367494 190226
rect 366874 190102 367494 190170
rect 366874 190046 366970 190102
rect 367026 190046 367094 190102
rect 367150 190046 367218 190102
rect 367274 190046 367342 190102
rect 367398 190046 367494 190102
rect 366874 189978 367494 190046
rect 366874 189922 366970 189978
rect 367026 189922 367094 189978
rect 367150 189922 367218 189978
rect 367274 189922 367342 189978
rect 367398 189922 367494 189978
rect 366874 172350 367494 189922
rect 366874 172294 366970 172350
rect 367026 172294 367094 172350
rect 367150 172294 367218 172350
rect 367274 172294 367342 172350
rect 367398 172294 367494 172350
rect 366874 172226 367494 172294
rect 366874 172170 366970 172226
rect 367026 172170 367094 172226
rect 367150 172170 367218 172226
rect 367274 172170 367342 172226
rect 367398 172170 367494 172226
rect 366874 172102 367494 172170
rect 366874 172046 366970 172102
rect 367026 172046 367094 172102
rect 367150 172046 367218 172102
rect 367274 172046 367342 172102
rect 367398 172046 367494 172102
rect 366874 171978 367494 172046
rect 366874 171922 366970 171978
rect 367026 171922 367094 171978
rect 367150 171922 367218 171978
rect 367274 171922 367342 171978
rect 367398 171922 367494 171978
rect 366874 154350 367494 171922
rect 366874 154294 366970 154350
rect 367026 154294 367094 154350
rect 367150 154294 367218 154350
rect 367274 154294 367342 154350
rect 367398 154294 367494 154350
rect 366874 154226 367494 154294
rect 366874 154170 366970 154226
rect 367026 154170 367094 154226
rect 367150 154170 367218 154226
rect 367274 154170 367342 154226
rect 367398 154170 367494 154226
rect 366874 154102 367494 154170
rect 366874 154046 366970 154102
rect 367026 154046 367094 154102
rect 367150 154046 367218 154102
rect 367274 154046 367342 154102
rect 367398 154046 367494 154102
rect 366874 153978 367494 154046
rect 366874 153922 366970 153978
rect 367026 153922 367094 153978
rect 367150 153922 367218 153978
rect 367274 153922 367342 153978
rect 367398 153922 367494 153978
rect 366874 136350 367494 153922
rect 366874 136294 366970 136350
rect 367026 136294 367094 136350
rect 367150 136294 367218 136350
rect 367274 136294 367342 136350
rect 367398 136294 367494 136350
rect 366874 136226 367494 136294
rect 366874 136170 366970 136226
rect 367026 136170 367094 136226
rect 367150 136170 367218 136226
rect 367274 136170 367342 136226
rect 367398 136170 367494 136226
rect 366874 136102 367494 136170
rect 366874 136046 366970 136102
rect 367026 136046 367094 136102
rect 367150 136046 367218 136102
rect 367274 136046 367342 136102
rect 367398 136046 367494 136102
rect 366874 135978 367494 136046
rect 366874 135922 366970 135978
rect 367026 135922 367094 135978
rect 367150 135922 367218 135978
rect 367274 135922 367342 135978
rect 367398 135922 367494 135978
rect 366874 118350 367494 135922
rect 366874 118294 366970 118350
rect 367026 118294 367094 118350
rect 367150 118294 367218 118350
rect 367274 118294 367342 118350
rect 367398 118294 367494 118350
rect 366874 118226 367494 118294
rect 366874 118170 366970 118226
rect 367026 118170 367094 118226
rect 367150 118170 367218 118226
rect 367274 118170 367342 118226
rect 367398 118170 367494 118226
rect 366874 118102 367494 118170
rect 366874 118046 366970 118102
rect 367026 118046 367094 118102
rect 367150 118046 367218 118102
rect 367274 118046 367342 118102
rect 367398 118046 367494 118102
rect 366874 117978 367494 118046
rect 366874 117922 366970 117978
rect 367026 117922 367094 117978
rect 367150 117922 367218 117978
rect 367274 117922 367342 117978
rect 367398 117922 367494 117978
rect 366874 100350 367494 117922
rect 366874 100294 366970 100350
rect 367026 100294 367094 100350
rect 367150 100294 367218 100350
rect 367274 100294 367342 100350
rect 367398 100294 367494 100350
rect 366874 100226 367494 100294
rect 366874 100170 366970 100226
rect 367026 100170 367094 100226
rect 367150 100170 367218 100226
rect 367274 100170 367342 100226
rect 367398 100170 367494 100226
rect 366874 100102 367494 100170
rect 366874 100046 366970 100102
rect 367026 100046 367094 100102
rect 367150 100046 367218 100102
rect 367274 100046 367342 100102
rect 367398 100046 367494 100102
rect 366874 99978 367494 100046
rect 366874 99922 366970 99978
rect 367026 99922 367094 99978
rect 367150 99922 367218 99978
rect 367274 99922 367342 99978
rect 367398 99922 367494 99978
rect 366874 82350 367494 99922
rect 366874 82294 366970 82350
rect 367026 82294 367094 82350
rect 367150 82294 367218 82350
rect 367274 82294 367342 82350
rect 367398 82294 367494 82350
rect 366874 82226 367494 82294
rect 366874 82170 366970 82226
rect 367026 82170 367094 82226
rect 367150 82170 367218 82226
rect 367274 82170 367342 82226
rect 367398 82170 367494 82226
rect 366874 82102 367494 82170
rect 366874 82046 366970 82102
rect 367026 82046 367094 82102
rect 367150 82046 367218 82102
rect 367274 82046 367342 82102
rect 367398 82046 367494 82102
rect 366874 81978 367494 82046
rect 366874 81922 366970 81978
rect 367026 81922 367094 81978
rect 367150 81922 367218 81978
rect 367274 81922 367342 81978
rect 367398 81922 367494 81978
rect 366874 64350 367494 81922
rect 366874 64294 366970 64350
rect 367026 64294 367094 64350
rect 367150 64294 367218 64350
rect 367274 64294 367342 64350
rect 367398 64294 367494 64350
rect 366874 64226 367494 64294
rect 366874 64170 366970 64226
rect 367026 64170 367094 64226
rect 367150 64170 367218 64226
rect 367274 64170 367342 64226
rect 367398 64170 367494 64226
rect 366874 64102 367494 64170
rect 366874 64046 366970 64102
rect 367026 64046 367094 64102
rect 367150 64046 367218 64102
rect 367274 64046 367342 64102
rect 367398 64046 367494 64102
rect 366874 63978 367494 64046
rect 366874 63922 366970 63978
rect 367026 63922 367094 63978
rect 367150 63922 367218 63978
rect 367274 63922 367342 63978
rect 367398 63922 367494 63978
rect 366874 46350 367494 63922
rect 366874 46294 366970 46350
rect 367026 46294 367094 46350
rect 367150 46294 367218 46350
rect 367274 46294 367342 46350
rect 367398 46294 367494 46350
rect 366874 46226 367494 46294
rect 366874 46170 366970 46226
rect 367026 46170 367094 46226
rect 367150 46170 367218 46226
rect 367274 46170 367342 46226
rect 367398 46170 367494 46226
rect 366874 46102 367494 46170
rect 366874 46046 366970 46102
rect 367026 46046 367094 46102
rect 367150 46046 367218 46102
rect 367274 46046 367342 46102
rect 367398 46046 367494 46102
rect 366874 45978 367494 46046
rect 366874 45922 366970 45978
rect 367026 45922 367094 45978
rect 367150 45922 367218 45978
rect 367274 45922 367342 45978
rect 367398 45922 367494 45978
rect 366874 28350 367494 45922
rect 366874 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 367494 28350
rect 366874 28226 367494 28294
rect 366874 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 367494 28226
rect 366874 28102 367494 28170
rect 366874 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 367494 28102
rect 366874 27978 367494 28046
rect 366874 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 367494 27978
rect 366874 10350 367494 27922
rect 366874 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 367494 10350
rect 366874 10226 367494 10294
rect 366874 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 367494 10226
rect 366874 10102 367494 10170
rect 366874 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 367494 10102
rect 366874 9978 367494 10046
rect 366874 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 367494 9978
rect 366874 -1120 367494 9922
rect 366874 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 367494 -1120
rect 366874 -1244 367494 -1176
rect 366874 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 367494 -1244
rect 366874 -1368 367494 -1300
rect 366874 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 367494 -1368
rect 366874 -1492 367494 -1424
rect 366874 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 367494 -1492
rect 366874 -1644 367494 -1548
rect 381154 202350 381774 210842
rect 381154 202294 381250 202350
rect 381306 202294 381374 202350
rect 381430 202294 381498 202350
rect 381554 202294 381622 202350
rect 381678 202294 381774 202350
rect 381154 202226 381774 202294
rect 381154 202170 381250 202226
rect 381306 202170 381374 202226
rect 381430 202170 381498 202226
rect 381554 202170 381622 202226
rect 381678 202170 381774 202226
rect 381154 202102 381774 202170
rect 381154 202046 381250 202102
rect 381306 202046 381374 202102
rect 381430 202046 381498 202102
rect 381554 202046 381622 202102
rect 381678 202046 381774 202102
rect 381154 201978 381774 202046
rect 381154 201922 381250 201978
rect 381306 201922 381374 201978
rect 381430 201922 381498 201978
rect 381554 201922 381622 201978
rect 381678 201922 381774 201978
rect 381154 184350 381774 201922
rect 381154 184294 381250 184350
rect 381306 184294 381374 184350
rect 381430 184294 381498 184350
rect 381554 184294 381622 184350
rect 381678 184294 381774 184350
rect 381154 184226 381774 184294
rect 381154 184170 381250 184226
rect 381306 184170 381374 184226
rect 381430 184170 381498 184226
rect 381554 184170 381622 184226
rect 381678 184170 381774 184226
rect 381154 184102 381774 184170
rect 381154 184046 381250 184102
rect 381306 184046 381374 184102
rect 381430 184046 381498 184102
rect 381554 184046 381622 184102
rect 381678 184046 381774 184102
rect 381154 183978 381774 184046
rect 381154 183922 381250 183978
rect 381306 183922 381374 183978
rect 381430 183922 381498 183978
rect 381554 183922 381622 183978
rect 381678 183922 381774 183978
rect 381154 166350 381774 183922
rect 381154 166294 381250 166350
rect 381306 166294 381374 166350
rect 381430 166294 381498 166350
rect 381554 166294 381622 166350
rect 381678 166294 381774 166350
rect 381154 166226 381774 166294
rect 381154 166170 381250 166226
rect 381306 166170 381374 166226
rect 381430 166170 381498 166226
rect 381554 166170 381622 166226
rect 381678 166170 381774 166226
rect 381154 166102 381774 166170
rect 381154 166046 381250 166102
rect 381306 166046 381374 166102
rect 381430 166046 381498 166102
rect 381554 166046 381622 166102
rect 381678 166046 381774 166102
rect 381154 165978 381774 166046
rect 381154 165922 381250 165978
rect 381306 165922 381374 165978
rect 381430 165922 381498 165978
rect 381554 165922 381622 165978
rect 381678 165922 381774 165978
rect 381154 148350 381774 165922
rect 381154 148294 381250 148350
rect 381306 148294 381374 148350
rect 381430 148294 381498 148350
rect 381554 148294 381622 148350
rect 381678 148294 381774 148350
rect 381154 148226 381774 148294
rect 381154 148170 381250 148226
rect 381306 148170 381374 148226
rect 381430 148170 381498 148226
rect 381554 148170 381622 148226
rect 381678 148170 381774 148226
rect 381154 148102 381774 148170
rect 381154 148046 381250 148102
rect 381306 148046 381374 148102
rect 381430 148046 381498 148102
rect 381554 148046 381622 148102
rect 381678 148046 381774 148102
rect 381154 147978 381774 148046
rect 381154 147922 381250 147978
rect 381306 147922 381374 147978
rect 381430 147922 381498 147978
rect 381554 147922 381622 147978
rect 381678 147922 381774 147978
rect 381154 130350 381774 147922
rect 381154 130294 381250 130350
rect 381306 130294 381374 130350
rect 381430 130294 381498 130350
rect 381554 130294 381622 130350
rect 381678 130294 381774 130350
rect 381154 130226 381774 130294
rect 381154 130170 381250 130226
rect 381306 130170 381374 130226
rect 381430 130170 381498 130226
rect 381554 130170 381622 130226
rect 381678 130170 381774 130226
rect 381154 130102 381774 130170
rect 381154 130046 381250 130102
rect 381306 130046 381374 130102
rect 381430 130046 381498 130102
rect 381554 130046 381622 130102
rect 381678 130046 381774 130102
rect 381154 129978 381774 130046
rect 381154 129922 381250 129978
rect 381306 129922 381374 129978
rect 381430 129922 381498 129978
rect 381554 129922 381622 129978
rect 381678 129922 381774 129978
rect 381154 112350 381774 129922
rect 381154 112294 381250 112350
rect 381306 112294 381374 112350
rect 381430 112294 381498 112350
rect 381554 112294 381622 112350
rect 381678 112294 381774 112350
rect 381154 112226 381774 112294
rect 381154 112170 381250 112226
rect 381306 112170 381374 112226
rect 381430 112170 381498 112226
rect 381554 112170 381622 112226
rect 381678 112170 381774 112226
rect 381154 112102 381774 112170
rect 381154 112046 381250 112102
rect 381306 112046 381374 112102
rect 381430 112046 381498 112102
rect 381554 112046 381622 112102
rect 381678 112046 381774 112102
rect 381154 111978 381774 112046
rect 381154 111922 381250 111978
rect 381306 111922 381374 111978
rect 381430 111922 381498 111978
rect 381554 111922 381622 111978
rect 381678 111922 381774 111978
rect 381154 94350 381774 111922
rect 381154 94294 381250 94350
rect 381306 94294 381374 94350
rect 381430 94294 381498 94350
rect 381554 94294 381622 94350
rect 381678 94294 381774 94350
rect 381154 94226 381774 94294
rect 381154 94170 381250 94226
rect 381306 94170 381374 94226
rect 381430 94170 381498 94226
rect 381554 94170 381622 94226
rect 381678 94170 381774 94226
rect 381154 94102 381774 94170
rect 381154 94046 381250 94102
rect 381306 94046 381374 94102
rect 381430 94046 381498 94102
rect 381554 94046 381622 94102
rect 381678 94046 381774 94102
rect 381154 93978 381774 94046
rect 381154 93922 381250 93978
rect 381306 93922 381374 93978
rect 381430 93922 381498 93978
rect 381554 93922 381622 93978
rect 381678 93922 381774 93978
rect 381154 76350 381774 93922
rect 381154 76294 381250 76350
rect 381306 76294 381374 76350
rect 381430 76294 381498 76350
rect 381554 76294 381622 76350
rect 381678 76294 381774 76350
rect 381154 76226 381774 76294
rect 381154 76170 381250 76226
rect 381306 76170 381374 76226
rect 381430 76170 381498 76226
rect 381554 76170 381622 76226
rect 381678 76170 381774 76226
rect 381154 76102 381774 76170
rect 381154 76046 381250 76102
rect 381306 76046 381374 76102
rect 381430 76046 381498 76102
rect 381554 76046 381622 76102
rect 381678 76046 381774 76102
rect 381154 75978 381774 76046
rect 381154 75922 381250 75978
rect 381306 75922 381374 75978
rect 381430 75922 381498 75978
rect 381554 75922 381622 75978
rect 381678 75922 381774 75978
rect 381154 58350 381774 75922
rect 381154 58294 381250 58350
rect 381306 58294 381374 58350
rect 381430 58294 381498 58350
rect 381554 58294 381622 58350
rect 381678 58294 381774 58350
rect 381154 58226 381774 58294
rect 381154 58170 381250 58226
rect 381306 58170 381374 58226
rect 381430 58170 381498 58226
rect 381554 58170 381622 58226
rect 381678 58170 381774 58226
rect 381154 58102 381774 58170
rect 381154 58046 381250 58102
rect 381306 58046 381374 58102
rect 381430 58046 381498 58102
rect 381554 58046 381622 58102
rect 381678 58046 381774 58102
rect 381154 57978 381774 58046
rect 381154 57922 381250 57978
rect 381306 57922 381374 57978
rect 381430 57922 381498 57978
rect 381554 57922 381622 57978
rect 381678 57922 381774 57978
rect 381154 40350 381774 57922
rect 381154 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 381774 40350
rect 381154 40226 381774 40294
rect 381154 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 381774 40226
rect 381154 40102 381774 40170
rect 381154 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 381774 40102
rect 381154 39978 381774 40046
rect 381154 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 381774 39978
rect 381154 22350 381774 39922
rect 381154 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 381774 22350
rect 381154 22226 381774 22294
rect 381154 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 381774 22226
rect 381154 22102 381774 22170
rect 381154 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 381774 22102
rect 381154 21978 381774 22046
rect 381154 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 381774 21978
rect 381154 4350 381774 21922
rect 381154 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 381774 4350
rect 381154 4226 381774 4294
rect 381154 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 381774 4226
rect 381154 4102 381774 4170
rect 381154 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 381774 4102
rect 381154 3978 381774 4046
rect 381154 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 381774 3978
rect 381154 -160 381774 3922
rect 381154 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 381774 -160
rect 381154 -284 381774 -216
rect 381154 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 381774 -284
rect 381154 -408 381774 -340
rect 381154 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 381774 -408
rect 381154 -532 381774 -464
rect 381154 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 381774 -532
rect 381154 -1644 381774 -588
rect 384874 208350 385494 210842
rect 384874 208294 384970 208350
rect 385026 208294 385094 208350
rect 385150 208294 385218 208350
rect 385274 208294 385342 208350
rect 385398 208294 385494 208350
rect 384874 208226 385494 208294
rect 384874 208170 384970 208226
rect 385026 208170 385094 208226
rect 385150 208170 385218 208226
rect 385274 208170 385342 208226
rect 385398 208170 385494 208226
rect 384874 208102 385494 208170
rect 384874 208046 384970 208102
rect 385026 208046 385094 208102
rect 385150 208046 385218 208102
rect 385274 208046 385342 208102
rect 385398 208046 385494 208102
rect 384874 207978 385494 208046
rect 384874 207922 384970 207978
rect 385026 207922 385094 207978
rect 385150 207922 385218 207978
rect 385274 207922 385342 207978
rect 385398 207922 385494 207978
rect 384874 190350 385494 207922
rect 384874 190294 384970 190350
rect 385026 190294 385094 190350
rect 385150 190294 385218 190350
rect 385274 190294 385342 190350
rect 385398 190294 385494 190350
rect 384874 190226 385494 190294
rect 384874 190170 384970 190226
rect 385026 190170 385094 190226
rect 385150 190170 385218 190226
rect 385274 190170 385342 190226
rect 385398 190170 385494 190226
rect 384874 190102 385494 190170
rect 384874 190046 384970 190102
rect 385026 190046 385094 190102
rect 385150 190046 385218 190102
rect 385274 190046 385342 190102
rect 385398 190046 385494 190102
rect 384874 189978 385494 190046
rect 384874 189922 384970 189978
rect 385026 189922 385094 189978
rect 385150 189922 385218 189978
rect 385274 189922 385342 189978
rect 385398 189922 385494 189978
rect 384874 172350 385494 189922
rect 384874 172294 384970 172350
rect 385026 172294 385094 172350
rect 385150 172294 385218 172350
rect 385274 172294 385342 172350
rect 385398 172294 385494 172350
rect 384874 172226 385494 172294
rect 384874 172170 384970 172226
rect 385026 172170 385094 172226
rect 385150 172170 385218 172226
rect 385274 172170 385342 172226
rect 385398 172170 385494 172226
rect 384874 172102 385494 172170
rect 384874 172046 384970 172102
rect 385026 172046 385094 172102
rect 385150 172046 385218 172102
rect 385274 172046 385342 172102
rect 385398 172046 385494 172102
rect 384874 171978 385494 172046
rect 384874 171922 384970 171978
rect 385026 171922 385094 171978
rect 385150 171922 385218 171978
rect 385274 171922 385342 171978
rect 385398 171922 385494 171978
rect 384874 154350 385494 171922
rect 384874 154294 384970 154350
rect 385026 154294 385094 154350
rect 385150 154294 385218 154350
rect 385274 154294 385342 154350
rect 385398 154294 385494 154350
rect 384874 154226 385494 154294
rect 384874 154170 384970 154226
rect 385026 154170 385094 154226
rect 385150 154170 385218 154226
rect 385274 154170 385342 154226
rect 385398 154170 385494 154226
rect 384874 154102 385494 154170
rect 384874 154046 384970 154102
rect 385026 154046 385094 154102
rect 385150 154046 385218 154102
rect 385274 154046 385342 154102
rect 385398 154046 385494 154102
rect 384874 153978 385494 154046
rect 384874 153922 384970 153978
rect 385026 153922 385094 153978
rect 385150 153922 385218 153978
rect 385274 153922 385342 153978
rect 385398 153922 385494 153978
rect 384874 136350 385494 153922
rect 384874 136294 384970 136350
rect 385026 136294 385094 136350
rect 385150 136294 385218 136350
rect 385274 136294 385342 136350
rect 385398 136294 385494 136350
rect 384874 136226 385494 136294
rect 384874 136170 384970 136226
rect 385026 136170 385094 136226
rect 385150 136170 385218 136226
rect 385274 136170 385342 136226
rect 385398 136170 385494 136226
rect 384874 136102 385494 136170
rect 384874 136046 384970 136102
rect 385026 136046 385094 136102
rect 385150 136046 385218 136102
rect 385274 136046 385342 136102
rect 385398 136046 385494 136102
rect 384874 135978 385494 136046
rect 384874 135922 384970 135978
rect 385026 135922 385094 135978
rect 385150 135922 385218 135978
rect 385274 135922 385342 135978
rect 385398 135922 385494 135978
rect 384874 118350 385494 135922
rect 384874 118294 384970 118350
rect 385026 118294 385094 118350
rect 385150 118294 385218 118350
rect 385274 118294 385342 118350
rect 385398 118294 385494 118350
rect 384874 118226 385494 118294
rect 384874 118170 384970 118226
rect 385026 118170 385094 118226
rect 385150 118170 385218 118226
rect 385274 118170 385342 118226
rect 385398 118170 385494 118226
rect 384874 118102 385494 118170
rect 384874 118046 384970 118102
rect 385026 118046 385094 118102
rect 385150 118046 385218 118102
rect 385274 118046 385342 118102
rect 385398 118046 385494 118102
rect 384874 117978 385494 118046
rect 384874 117922 384970 117978
rect 385026 117922 385094 117978
rect 385150 117922 385218 117978
rect 385274 117922 385342 117978
rect 385398 117922 385494 117978
rect 384874 100350 385494 117922
rect 384874 100294 384970 100350
rect 385026 100294 385094 100350
rect 385150 100294 385218 100350
rect 385274 100294 385342 100350
rect 385398 100294 385494 100350
rect 384874 100226 385494 100294
rect 384874 100170 384970 100226
rect 385026 100170 385094 100226
rect 385150 100170 385218 100226
rect 385274 100170 385342 100226
rect 385398 100170 385494 100226
rect 384874 100102 385494 100170
rect 384874 100046 384970 100102
rect 385026 100046 385094 100102
rect 385150 100046 385218 100102
rect 385274 100046 385342 100102
rect 385398 100046 385494 100102
rect 384874 99978 385494 100046
rect 384874 99922 384970 99978
rect 385026 99922 385094 99978
rect 385150 99922 385218 99978
rect 385274 99922 385342 99978
rect 385398 99922 385494 99978
rect 384874 82350 385494 99922
rect 384874 82294 384970 82350
rect 385026 82294 385094 82350
rect 385150 82294 385218 82350
rect 385274 82294 385342 82350
rect 385398 82294 385494 82350
rect 384874 82226 385494 82294
rect 384874 82170 384970 82226
rect 385026 82170 385094 82226
rect 385150 82170 385218 82226
rect 385274 82170 385342 82226
rect 385398 82170 385494 82226
rect 384874 82102 385494 82170
rect 384874 82046 384970 82102
rect 385026 82046 385094 82102
rect 385150 82046 385218 82102
rect 385274 82046 385342 82102
rect 385398 82046 385494 82102
rect 384874 81978 385494 82046
rect 384874 81922 384970 81978
rect 385026 81922 385094 81978
rect 385150 81922 385218 81978
rect 385274 81922 385342 81978
rect 385398 81922 385494 81978
rect 384874 64350 385494 81922
rect 384874 64294 384970 64350
rect 385026 64294 385094 64350
rect 385150 64294 385218 64350
rect 385274 64294 385342 64350
rect 385398 64294 385494 64350
rect 384874 64226 385494 64294
rect 384874 64170 384970 64226
rect 385026 64170 385094 64226
rect 385150 64170 385218 64226
rect 385274 64170 385342 64226
rect 385398 64170 385494 64226
rect 384874 64102 385494 64170
rect 384874 64046 384970 64102
rect 385026 64046 385094 64102
rect 385150 64046 385218 64102
rect 385274 64046 385342 64102
rect 385398 64046 385494 64102
rect 384874 63978 385494 64046
rect 384874 63922 384970 63978
rect 385026 63922 385094 63978
rect 385150 63922 385218 63978
rect 385274 63922 385342 63978
rect 385398 63922 385494 63978
rect 384874 46350 385494 63922
rect 384874 46294 384970 46350
rect 385026 46294 385094 46350
rect 385150 46294 385218 46350
rect 385274 46294 385342 46350
rect 385398 46294 385494 46350
rect 384874 46226 385494 46294
rect 384874 46170 384970 46226
rect 385026 46170 385094 46226
rect 385150 46170 385218 46226
rect 385274 46170 385342 46226
rect 385398 46170 385494 46226
rect 384874 46102 385494 46170
rect 384874 46046 384970 46102
rect 385026 46046 385094 46102
rect 385150 46046 385218 46102
rect 385274 46046 385342 46102
rect 385398 46046 385494 46102
rect 384874 45978 385494 46046
rect 384874 45922 384970 45978
rect 385026 45922 385094 45978
rect 385150 45922 385218 45978
rect 385274 45922 385342 45978
rect 385398 45922 385494 45978
rect 384874 28350 385494 45922
rect 384874 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 385494 28350
rect 384874 28226 385494 28294
rect 384874 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 385494 28226
rect 384874 28102 385494 28170
rect 384874 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 385494 28102
rect 384874 27978 385494 28046
rect 384874 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 385494 27978
rect 384874 10350 385494 27922
rect 384874 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 385494 10350
rect 384874 10226 385494 10294
rect 384874 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 385494 10226
rect 384874 10102 385494 10170
rect 384874 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 385494 10102
rect 384874 9978 385494 10046
rect 384874 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 385494 9978
rect 384874 -1120 385494 9922
rect 384874 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 385494 -1120
rect 384874 -1244 385494 -1176
rect 384874 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 385494 -1244
rect 384874 -1368 385494 -1300
rect 384874 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 385494 -1368
rect 384874 -1492 385494 -1424
rect 384874 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 385494 -1492
rect 384874 -1644 385494 -1548
rect 399154 202350 399774 210842
rect 399154 202294 399250 202350
rect 399306 202294 399374 202350
rect 399430 202294 399498 202350
rect 399554 202294 399622 202350
rect 399678 202294 399774 202350
rect 399154 202226 399774 202294
rect 399154 202170 399250 202226
rect 399306 202170 399374 202226
rect 399430 202170 399498 202226
rect 399554 202170 399622 202226
rect 399678 202170 399774 202226
rect 399154 202102 399774 202170
rect 399154 202046 399250 202102
rect 399306 202046 399374 202102
rect 399430 202046 399498 202102
rect 399554 202046 399622 202102
rect 399678 202046 399774 202102
rect 399154 201978 399774 202046
rect 399154 201922 399250 201978
rect 399306 201922 399374 201978
rect 399430 201922 399498 201978
rect 399554 201922 399622 201978
rect 399678 201922 399774 201978
rect 399154 184350 399774 201922
rect 399154 184294 399250 184350
rect 399306 184294 399374 184350
rect 399430 184294 399498 184350
rect 399554 184294 399622 184350
rect 399678 184294 399774 184350
rect 399154 184226 399774 184294
rect 399154 184170 399250 184226
rect 399306 184170 399374 184226
rect 399430 184170 399498 184226
rect 399554 184170 399622 184226
rect 399678 184170 399774 184226
rect 399154 184102 399774 184170
rect 399154 184046 399250 184102
rect 399306 184046 399374 184102
rect 399430 184046 399498 184102
rect 399554 184046 399622 184102
rect 399678 184046 399774 184102
rect 399154 183978 399774 184046
rect 399154 183922 399250 183978
rect 399306 183922 399374 183978
rect 399430 183922 399498 183978
rect 399554 183922 399622 183978
rect 399678 183922 399774 183978
rect 399154 166350 399774 183922
rect 399154 166294 399250 166350
rect 399306 166294 399374 166350
rect 399430 166294 399498 166350
rect 399554 166294 399622 166350
rect 399678 166294 399774 166350
rect 399154 166226 399774 166294
rect 399154 166170 399250 166226
rect 399306 166170 399374 166226
rect 399430 166170 399498 166226
rect 399554 166170 399622 166226
rect 399678 166170 399774 166226
rect 399154 166102 399774 166170
rect 399154 166046 399250 166102
rect 399306 166046 399374 166102
rect 399430 166046 399498 166102
rect 399554 166046 399622 166102
rect 399678 166046 399774 166102
rect 399154 165978 399774 166046
rect 399154 165922 399250 165978
rect 399306 165922 399374 165978
rect 399430 165922 399498 165978
rect 399554 165922 399622 165978
rect 399678 165922 399774 165978
rect 399154 148350 399774 165922
rect 399154 148294 399250 148350
rect 399306 148294 399374 148350
rect 399430 148294 399498 148350
rect 399554 148294 399622 148350
rect 399678 148294 399774 148350
rect 399154 148226 399774 148294
rect 399154 148170 399250 148226
rect 399306 148170 399374 148226
rect 399430 148170 399498 148226
rect 399554 148170 399622 148226
rect 399678 148170 399774 148226
rect 399154 148102 399774 148170
rect 399154 148046 399250 148102
rect 399306 148046 399374 148102
rect 399430 148046 399498 148102
rect 399554 148046 399622 148102
rect 399678 148046 399774 148102
rect 399154 147978 399774 148046
rect 399154 147922 399250 147978
rect 399306 147922 399374 147978
rect 399430 147922 399498 147978
rect 399554 147922 399622 147978
rect 399678 147922 399774 147978
rect 399154 130350 399774 147922
rect 399154 130294 399250 130350
rect 399306 130294 399374 130350
rect 399430 130294 399498 130350
rect 399554 130294 399622 130350
rect 399678 130294 399774 130350
rect 399154 130226 399774 130294
rect 399154 130170 399250 130226
rect 399306 130170 399374 130226
rect 399430 130170 399498 130226
rect 399554 130170 399622 130226
rect 399678 130170 399774 130226
rect 399154 130102 399774 130170
rect 399154 130046 399250 130102
rect 399306 130046 399374 130102
rect 399430 130046 399498 130102
rect 399554 130046 399622 130102
rect 399678 130046 399774 130102
rect 399154 129978 399774 130046
rect 399154 129922 399250 129978
rect 399306 129922 399374 129978
rect 399430 129922 399498 129978
rect 399554 129922 399622 129978
rect 399678 129922 399774 129978
rect 399154 112350 399774 129922
rect 399154 112294 399250 112350
rect 399306 112294 399374 112350
rect 399430 112294 399498 112350
rect 399554 112294 399622 112350
rect 399678 112294 399774 112350
rect 399154 112226 399774 112294
rect 399154 112170 399250 112226
rect 399306 112170 399374 112226
rect 399430 112170 399498 112226
rect 399554 112170 399622 112226
rect 399678 112170 399774 112226
rect 399154 112102 399774 112170
rect 399154 112046 399250 112102
rect 399306 112046 399374 112102
rect 399430 112046 399498 112102
rect 399554 112046 399622 112102
rect 399678 112046 399774 112102
rect 399154 111978 399774 112046
rect 399154 111922 399250 111978
rect 399306 111922 399374 111978
rect 399430 111922 399498 111978
rect 399554 111922 399622 111978
rect 399678 111922 399774 111978
rect 399154 94350 399774 111922
rect 399154 94294 399250 94350
rect 399306 94294 399374 94350
rect 399430 94294 399498 94350
rect 399554 94294 399622 94350
rect 399678 94294 399774 94350
rect 399154 94226 399774 94294
rect 399154 94170 399250 94226
rect 399306 94170 399374 94226
rect 399430 94170 399498 94226
rect 399554 94170 399622 94226
rect 399678 94170 399774 94226
rect 399154 94102 399774 94170
rect 399154 94046 399250 94102
rect 399306 94046 399374 94102
rect 399430 94046 399498 94102
rect 399554 94046 399622 94102
rect 399678 94046 399774 94102
rect 399154 93978 399774 94046
rect 399154 93922 399250 93978
rect 399306 93922 399374 93978
rect 399430 93922 399498 93978
rect 399554 93922 399622 93978
rect 399678 93922 399774 93978
rect 399154 76350 399774 93922
rect 399154 76294 399250 76350
rect 399306 76294 399374 76350
rect 399430 76294 399498 76350
rect 399554 76294 399622 76350
rect 399678 76294 399774 76350
rect 399154 76226 399774 76294
rect 399154 76170 399250 76226
rect 399306 76170 399374 76226
rect 399430 76170 399498 76226
rect 399554 76170 399622 76226
rect 399678 76170 399774 76226
rect 399154 76102 399774 76170
rect 399154 76046 399250 76102
rect 399306 76046 399374 76102
rect 399430 76046 399498 76102
rect 399554 76046 399622 76102
rect 399678 76046 399774 76102
rect 399154 75978 399774 76046
rect 399154 75922 399250 75978
rect 399306 75922 399374 75978
rect 399430 75922 399498 75978
rect 399554 75922 399622 75978
rect 399678 75922 399774 75978
rect 399154 58350 399774 75922
rect 399154 58294 399250 58350
rect 399306 58294 399374 58350
rect 399430 58294 399498 58350
rect 399554 58294 399622 58350
rect 399678 58294 399774 58350
rect 399154 58226 399774 58294
rect 399154 58170 399250 58226
rect 399306 58170 399374 58226
rect 399430 58170 399498 58226
rect 399554 58170 399622 58226
rect 399678 58170 399774 58226
rect 399154 58102 399774 58170
rect 399154 58046 399250 58102
rect 399306 58046 399374 58102
rect 399430 58046 399498 58102
rect 399554 58046 399622 58102
rect 399678 58046 399774 58102
rect 399154 57978 399774 58046
rect 399154 57922 399250 57978
rect 399306 57922 399374 57978
rect 399430 57922 399498 57978
rect 399554 57922 399622 57978
rect 399678 57922 399774 57978
rect 399154 40350 399774 57922
rect 399154 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 399774 40350
rect 399154 40226 399774 40294
rect 399154 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 399774 40226
rect 399154 40102 399774 40170
rect 399154 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 399774 40102
rect 399154 39978 399774 40046
rect 399154 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 399774 39978
rect 399154 22350 399774 39922
rect 399154 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 399774 22350
rect 399154 22226 399774 22294
rect 399154 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 399774 22226
rect 399154 22102 399774 22170
rect 399154 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 399774 22102
rect 399154 21978 399774 22046
rect 399154 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 399774 21978
rect 399154 4350 399774 21922
rect 399154 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 399774 4350
rect 399154 4226 399774 4294
rect 399154 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 399774 4226
rect 399154 4102 399774 4170
rect 399154 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 399774 4102
rect 399154 3978 399774 4046
rect 399154 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 399774 3978
rect 399154 -160 399774 3922
rect 399154 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 399774 -160
rect 399154 -284 399774 -216
rect 399154 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 399774 -284
rect 399154 -408 399774 -340
rect 399154 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 399774 -408
rect 399154 -532 399774 -464
rect 399154 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 399774 -532
rect 399154 -1644 399774 -588
rect 402874 208350 403494 210842
rect 402874 208294 402970 208350
rect 403026 208294 403094 208350
rect 403150 208294 403218 208350
rect 403274 208294 403342 208350
rect 403398 208294 403494 208350
rect 402874 208226 403494 208294
rect 402874 208170 402970 208226
rect 403026 208170 403094 208226
rect 403150 208170 403218 208226
rect 403274 208170 403342 208226
rect 403398 208170 403494 208226
rect 402874 208102 403494 208170
rect 402874 208046 402970 208102
rect 403026 208046 403094 208102
rect 403150 208046 403218 208102
rect 403274 208046 403342 208102
rect 403398 208046 403494 208102
rect 402874 207978 403494 208046
rect 402874 207922 402970 207978
rect 403026 207922 403094 207978
rect 403150 207922 403218 207978
rect 403274 207922 403342 207978
rect 403398 207922 403494 207978
rect 402874 190350 403494 207922
rect 404128 208350 404448 208384
rect 404128 208294 404198 208350
rect 404254 208294 404322 208350
rect 404378 208294 404448 208350
rect 404128 208226 404448 208294
rect 404128 208170 404198 208226
rect 404254 208170 404322 208226
rect 404378 208170 404448 208226
rect 404128 208102 404448 208170
rect 404128 208046 404198 208102
rect 404254 208046 404322 208102
rect 404378 208046 404448 208102
rect 404128 207978 404448 208046
rect 404128 207922 404198 207978
rect 404254 207922 404322 207978
rect 404378 207922 404448 207978
rect 404128 207888 404448 207922
rect 402874 190294 402970 190350
rect 403026 190294 403094 190350
rect 403150 190294 403218 190350
rect 403274 190294 403342 190350
rect 403398 190294 403494 190350
rect 402874 190226 403494 190294
rect 402874 190170 402970 190226
rect 403026 190170 403094 190226
rect 403150 190170 403218 190226
rect 403274 190170 403342 190226
rect 403398 190170 403494 190226
rect 402874 190102 403494 190170
rect 402874 190046 402970 190102
rect 403026 190046 403094 190102
rect 403150 190046 403218 190102
rect 403274 190046 403342 190102
rect 403398 190046 403494 190102
rect 402874 189978 403494 190046
rect 402874 189922 402970 189978
rect 403026 189922 403094 189978
rect 403150 189922 403218 189978
rect 403274 189922 403342 189978
rect 403398 189922 403494 189978
rect 402874 172350 403494 189922
rect 402874 172294 402970 172350
rect 403026 172294 403094 172350
rect 403150 172294 403218 172350
rect 403274 172294 403342 172350
rect 403398 172294 403494 172350
rect 402874 172226 403494 172294
rect 402874 172170 402970 172226
rect 403026 172170 403094 172226
rect 403150 172170 403218 172226
rect 403274 172170 403342 172226
rect 403398 172170 403494 172226
rect 402874 172102 403494 172170
rect 402874 172046 402970 172102
rect 403026 172046 403094 172102
rect 403150 172046 403218 172102
rect 403274 172046 403342 172102
rect 403398 172046 403494 172102
rect 402874 171978 403494 172046
rect 402874 171922 402970 171978
rect 403026 171922 403094 171978
rect 403150 171922 403218 171978
rect 403274 171922 403342 171978
rect 403398 171922 403494 171978
rect 402874 154350 403494 171922
rect 402874 154294 402970 154350
rect 403026 154294 403094 154350
rect 403150 154294 403218 154350
rect 403274 154294 403342 154350
rect 403398 154294 403494 154350
rect 402874 154226 403494 154294
rect 402874 154170 402970 154226
rect 403026 154170 403094 154226
rect 403150 154170 403218 154226
rect 403274 154170 403342 154226
rect 403398 154170 403494 154226
rect 402874 154102 403494 154170
rect 402874 154046 402970 154102
rect 403026 154046 403094 154102
rect 403150 154046 403218 154102
rect 403274 154046 403342 154102
rect 403398 154046 403494 154102
rect 402874 153978 403494 154046
rect 402874 153922 402970 153978
rect 403026 153922 403094 153978
rect 403150 153922 403218 153978
rect 403274 153922 403342 153978
rect 403398 153922 403494 153978
rect 402874 136350 403494 153922
rect 402874 136294 402970 136350
rect 403026 136294 403094 136350
rect 403150 136294 403218 136350
rect 403274 136294 403342 136350
rect 403398 136294 403494 136350
rect 402874 136226 403494 136294
rect 402874 136170 402970 136226
rect 403026 136170 403094 136226
rect 403150 136170 403218 136226
rect 403274 136170 403342 136226
rect 403398 136170 403494 136226
rect 402874 136102 403494 136170
rect 402874 136046 402970 136102
rect 403026 136046 403094 136102
rect 403150 136046 403218 136102
rect 403274 136046 403342 136102
rect 403398 136046 403494 136102
rect 402874 135978 403494 136046
rect 402874 135922 402970 135978
rect 403026 135922 403094 135978
rect 403150 135922 403218 135978
rect 403274 135922 403342 135978
rect 403398 135922 403494 135978
rect 402874 118350 403494 135922
rect 402874 118294 402970 118350
rect 403026 118294 403094 118350
rect 403150 118294 403218 118350
rect 403274 118294 403342 118350
rect 403398 118294 403494 118350
rect 402874 118226 403494 118294
rect 402874 118170 402970 118226
rect 403026 118170 403094 118226
rect 403150 118170 403218 118226
rect 403274 118170 403342 118226
rect 403398 118170 403494 118226
rect 402874 118102 403494 118170
rect 402874 118046 402970 118102
rect 403026 118046 403094 118102
rect 403150 118046 403218 118102
rect 403274 118046 403342 118102
rect 403398 118046 403494 118102
rect 402874 117978 403494 118046
rect 402874 117922 402970 117978
rect 403026 117922 403094 117978
rect 403150 117922 403218 117978
rect 403274 117922 403342 117978
rect 403398 117922 403494 117978
rect 402874 100350 403494 117922
rect 402874 100294 402970 100350
rect 403026 100294 403094 100350
rect 403150 100294 403218 100350
rect 403274 100294 403342 100350
rect 403398 100294 403494 100350
rect 402874 100226 403494 100294
rect 402874 100170 402970 100226
rect 403026 100170 403094 100226
rect 403150 100170 403218 100226
rect 403274 100170 403342 100226
rect 403398 100170 403494 100226
rect 402874 100102 403494 100170
rect 402874 100046 402970 100102
rect 403026 100046 403094 100102
rect 403150 100046 403218 100102
rect 403274 100046 403342 100102
rect 403398 100046 403494 100102
rect 402874 99978 403494 100046
rect 402874 99922 402970 99978
rect 403026 99922 403094 99978
rect 403150 99922 403218 99978
rect 403274 99922 403342 99978
rect 403398 99922 403494 99978
rect 402874 82350 403494 99922
rect 402874 82294 402970 82350
rect 403026 82294 403094 82350
rect 403150 82294 403218 82350
rect 403274 82294 403342 82350
rect 403398 82294 403494 82350
rect 402874 82226 403494 82294
rect 402874 82170 402970 82226
rect 403026 82170 403094 82226
rect 403150 82170 403218 82226
rect 403274 82170 403342 82226
rect 403398 82170 403494 82226
rect 402874 82102 403494 82170
rect 402874 82046 402970 82102
rect 403026 82046 403094 82102
rect 403150 82046 403218 82102
rect 403274 82046 403342 82102
rect 403398 82046 403494 82102
rect 402874 81978 403494 82046
rect 402874 81922 402970 81978
rect 403026 81922 403094 81978
rect 403150 81922 403218 81978
rect 403274 81922 403342 81978
rect 403398 81922 403494 81978
rect 402874 64350 403494 81922
rect 402874 64294 402970 64350
rect 403026 64294 403094 64350
rect 403150 64294 403218 64350
rect 403274 64294 403342 64350
rect 403398 64294 403494 64350
rect 402874 64226 403494 64294
rect 402874 64170 402970 64226
rect 403026 64170 403094 64226
rect 403150 64170 403218 64226
rect 403274 64170 403342 64226
rect 403398 64170 403494 64226
rect 402874 64102 403494 64170
rect 402874 64046 402970 64102
rect 403026 64046 403094 64102
rect 403150 64046 403218 64102
rect 403274 64046 403342 64102
rect 403398 64046 403494 64102
rect 402874 63978 403494 64046
rect 402874 63922 402970 63978
rect 403026 63922 403094 63978
rect 403150 63922 403218 63978
rect 403274 63922 403342 63978
rect 403398 63922 403494 63978
rect 402874 46350 403494 63922
rect 402874 46294 402970 46350
rect 403026 46294 403094 46350
rect 403150 46294 403218 46350
rect 403274 46294 403342 46350
rect 403398 46294 403494 46350
rect 402874 46226 403494 46294
rect 402874 46170 402970 46226
rect 403026 46170 403094 46226
rect 403150 46170 403218 46226
rect 403274 46170 403342 46226
rect 403398 46170 403494 46226
rect 402874 46102 403494 46170
rect 402874 46046 402970 46102
rect 403026 46046 403094 46102
rect 403150 46046 403218 46102
rect 403274 46046 403342 46102
rect 403398 46046 403494 46102
rect 402874 45978 403494 46046
rect 402874 45922 402970 45978
rect 403026 45922 403094 45978
rect 403150 45922 403218 45978
rect 403274 45922 403342 45978
rect 403398 45922 403494 45978
rect 402874 28350 403494 45922
rect 402874 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 403494 28350
rect 402874 28226 403494 28294
rect 402874 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 403494 28226
rect 402874 28102 403494 28170
rect 402874 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 403494 28102
rect 402874 27978 403494 28046
rect 402874 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 403494 27978
rect 402874 10350 403494 27922
rect 402874 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 403494 10350
rect 402874 10226 403494 10294
rect 402874 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 403494 10226
rect 402874 10102 403494 10170
rect 402874 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 403494 10102
rect 402874 9978 403494 10046
rect 402874 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 403494 9978
rect 402874 -1120 403494 9922
rect 402874 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 403494 -1120
rect 402874 -1244 403494 -1176
rect 402874 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 403494 -1244
rect 402874 -1368 403494 -1300
rect 402874 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 403494 -1368
rect 402874 -1492 403494 -1424
rect 402874 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 403494 -1492
rect 402874 -1644 403494 -1548
rect 417154 202350 417774 210842
rect 417154 202294 417250 202350
rect 417306 202294 417374 202350
rect 417430 202294 417498 202350
rect 417554 202294 417622 202350
rect 417678 202294 417774 202350
rect 417154 202226 417774 202294
rect 417154 202170 417250 202226
rect 417306 202170 417374 202226
rect 417430 202170 417498 202226
rect 417554 202170 417622 202226
rect 417678 202170 417774 202226
rect 417154 202102 417774 202170
rect 417154 202046 417250 202102
rect 417306 202046 417374 202102
rect 417430 202046 417498 202102
rect 417554 202046 417622 202102
rect 417678 202046 417774 202102
rect 417154 201978 417774 202046
rect 417154 201922 417250 201978
rect 417306 201922 417374 201978
rect 417430 201922 417498 201978
rect 417554 201922 417622 201978
rect 417678 201922 417774 201978
rect 417154 184350 417774 201922
rect 417154 184294 417250 184350
rect 417306 184294 417374 184350
rect 417430 184294 417498 184350
rect 417554 184294 417622 184350
rect 417678 184294 417774 184350
rect 417154 184226 417774 184294
rect 417154 184170 417250 184226
rect 417306 184170 417374 184226
rect 417430 184170 417498 184226
rect 417554 184170 417622 184226
rect 417678 184170 417774 184226
rect 417154 184102 417774 184170
rect 417154 184046 417250 184102
rect 417306 184046 417374 184102
rect 417430 184046 417498 184102
rect 417554 184046 417622 184102
rect 417678 184046 417774 184102
rect 417154 183978 417774 184046
rect 417154 183922 417250 183978
rect 417306 183922 417374 183978
rect 417430 183922 417498 183978
rect 417554 183922 417622 183978
rect 417678 183922 417774 183978
rect 417154 166350 417774 183922
rect 417154 166294 417250 166350
rect 417306 166294 417374 166350
rect 417430 166294 417498 166350
rect 417554 166294 417622 166350
rect 417678 166294 417774 166350
rect 417154 166226 417774 166294
rect 417154 166170 417250 166226
rect 417306 166170 417374 166226
rect 417430 166170 417498 166226
rect 417554 166170 417622 166226
rect 417678 166170 417774 166226
rect 417154 166102 417774 166170
rect 417154 166046 417250 166102
rect 417306 166046 417374 166102
rect 417430 166046 417498 166102
rect 417554 166046 417622 166102
rect 417678 166046 417774 166102
rect 417154 165978 417774 166046
rect 417154 165922 417250 165978
rect 417306 165922 417374 165978
rect 417430 165922 417498 165978
rect 417554 165922 417622 165978
rect 417678 165922 417774 165978
rect 417154 148350 417774 165922
rect 417154 148294 417250 148350
rect 417306 148294 417374 148350
rect 417430 148294 417498 148350
rect 417554 148294 417622 148350
rect 417678 148294 417774 148350
rect 417154 148226 417774 148294
rect 417154 148170 417250 148226
rect 417306 148170 417374 148226
rect 417430 148170 417498 148226
rect 417554 148170 417622 148226
rect 417678 148170 417774 148226
rect 417154 148102 417774 148170
rect 417154 148046 417250 148102
rect 417306 148046 417374 148102
rect 417430 148046 417498 148102
rect 417554 148046 417622 148102
rect 417678 148046 417774 148102
rect 417154 147978 417774 148046
rect 417154 147922 417250 147978
rect 417306 147922 417374 147978
rect 417430 147922 417498 147978
rect 417554 147922 417622 147978
rect 417678 147922 417774 147978
rect 417154 130350 417774 147922
rect 417154 130294 417250 130350
rect 417306 130294 417374 130350
rect 417430 130294 417498 130350
rect 417554 130294 417622 130350
rect 417678 130294 417774 130350
rect 417154 130226 417774 130294
rect 417154 130170 417250 130226
rect 417306 130170 417374 130226
rect 417430 130170 417498 130226
rect 417554 130170 417622 130226
rect 417678 130170 417774 130226
rect 417154 130102 417774 130170
rect 417154 130046 417250 130102
rect 417306 130046 417374 130102
rect 417430 130046 417498 130102
rect 417554 130046 417622 130102
rect 417678 130046 417774 130102
rect 417154 129978 417774 130046
rect 417154 129922 417250 129978
rect 417306 129922 417374 129978
rect 417430 129922 417498 129978
rect 417554 129922 417622 129978
rect 417678 129922 417774 129978
rect 417154 112350 417774 129922
rect 417154 112294 417250 112350
rect 417306 112294 417374 112350
rect 417430 112294 417498 112350
rect 417554 112294 417622 112350
rect 417678 112294 417774 112350
rect 417154 112226 417774 112294
rect 417154 112170 417250 112226
rect 417306 112170 417374 112226
rect 417430 112170 417498 112226
rect 417554 112170 417622 112226
rect 417678 112170 417774 112226
rect 417154 112102 417774 112170
rect 417154 112046 417250 112102
rect 417306 112046 417374 112102
rect 417430 112046 417498 112102
rect 417554 112046 417622 112102
rect 417678 112046 417774 112102
rect 417154 111978 417774 112046
rect 417154 111922 417250 111978
rect 417306 111922 417374 111978
rect 417430 111922 417498 111978
rect 417554 111922 417622 111978
rect 417678 111922 417774 111978
rect 417154 94350 417774 111922
rect 417154 94294 417250 94350
rect 417306 94294 417374 94350
rect 417430 94294 417498 94350
rect 417554 94294 417622 94350
rect 417678 94294 417774 94350
rect 417154 94226 417774 94294
rect 417154 94170 417250 94226
rect 417306 94170 417374 94226
rect 417430 94170 417498 94226
rect 417554 94170 417622 94226
rect 417678 94170 417774 94226
rect 417154 94102 417774 94170
rect 417154 94046 417250 94102
rect 417306 94046 417374 94102
rect 417430 94046 417498 94102
rect 417554 94046 417622 94102
rect 417678 94046 417774 94102
rect 417154 93978 417774 94046
rect 417154 93922 417250 93978
rect 417306 93922 417374 93978
rect 417430 93922 417498 93978
rect 417554 93922 417622 93978
rect 417678 93922 417774 93978
rect 417154 76350 417774 93922
rect 417154 76294 417250 76350
rect 417306 76294 417374 76350
rect 417430 76294 417498 76350
rect 417554 76294 417622 76350
rect 417678 76294 417774 76350
rect 417154 76226 417774 76294
rect 417154 76170 417250 76226
rect 417306 76170 417374 76226
rect 417430 76170 417498 76226
rect 417554 76170 417622 76226
rect 417678 76170 417774 76226
rect 417154 76102 417774 76170
rect 417154 76046 417250 76102
rect 417306 76046 417374 76102
rect 417430 76046 417498 76102
rect 417554 76046 417622 76102
rect 417678 76046 417774 76102
rect 417154 75978 417774 76046
rect 417154 75922 417250 75978
rect 417306 75922 417374 75978
rect 417430 75922 417498 75978
rect 417554 75922 417622 75978
rect 417678 75922 417774 75978
rect 417154 58350 417774 75922
rect 417154 58294 417250 58350
rect 417306 58294 417374 58350
rect 417430 58294 417498 58350
rect 417554 58294 417622 58350
rect 417678 58294 417774 58350
rect 417154 58226 417774 58294
rect 417154 58170 417250 58226
rect 417306 58170 417374 58226
rect 417430 58170 417498 58226
rect 417554 58170 417622 58226
rect 417678 58170 417774 58226
rect 417154 58102 417774 58170
rect 417154 58046 417250 58102
rect 417306 58046 417374 58102
rect 417430 58046 417498 58102
rect 417554 58046 417622 58102
rect 417678 58046 417774 58102
rect 417154 57978 417774 58046
rect 417154 57922 417250 57978
rect 417306 57922 417374 57978
rect 417430 57922 417498 57978
rect 417554 57922 417622 57978
rect 417678 57922 417774 57978
rect 417154 40350 417774 57922
rect 417154 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 417774 40350
rect 417154 40226 417774 40294
rect 417154 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 417774 40226
rect 417154 40102 417774 40170
rect 417154 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 417774 40102
rect 417154 39978 417774 40046
rect 417154 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 417774 39978
rect 417154 22350 417774 39922
rect 417154 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 417774 22350
rect 417154 22226 417774 22294
rect 417154 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 417774 22226
rect 417154 22102 417774 22170
rect 417154 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 417774 22102
rect 417154 21978 417774 22046
rect 417154 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 417774 21978
rect 417154 4350 417774 21922
rect 417154 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 417774 4350
rect 417154 4226 417774 4294
rect 417154 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 417774 4226
rect 417154 4102 417774 4170
rect 417154 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 417774 4102
rect 417154 3978 417774 4046
rect 417154 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 417774 3978
rect 417154 -160 417774 3922
rect 417154 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 417774 -160
rect 417154 -284 417774 -216
rect 417154 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 417774 -284
rect 417154 -408 417774 -340
rect 417154 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 417774 -408
rect 417154 -532 417774 -464
rect 417154 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 417774 -532
rect 417154 -1644 417774 -588
rect 420874 208350 421494 210842
rect 420874 208294 420970 208350
rect 421026 208294 421094 208350
rect 421150 208294 421218 208350
rect 421274 208294 421342 208350
rect 421398 208294 421494 208350
rect 420874 208226 421494 208294
rect 420874 208170 420970 208226
rect 421026 208170 421094 208226
rect 421150 208170 421218 208226
rect 421274 208170 421342 208226
rect 421398 208170 421494 208226
rect 420874 208102 421494 208170
rect 420874 208046 420970 208102
rect 421026 208046 421094 208102
rect 421150 208046 421218 208102
rect 421274 208046 421342 208102
rect 421398 208046 421494 208102
rect 420874 207978 421494 208046
rect 420874 207922 420970 207978
rect 421026 207922 421094 207978
rect 421150 207922 421218 207978
rect 421274 207922 421342 207978
rect 421398 207922 421494 207978
rect 420874 190350 421494 207922
rect 434848 208350 435168 208384
rect 434848 208294 434918 208350
rect 434974 208294 435042 208350
rect 435098 208294 435168 208350
rect 434848 208226 435168 208294
rect 434848 208170 434918 208226
rect 434974 208170 435042 208226
rect 435098 208170 435168 208226
rect 434848 208102 435168 208170
rect 434848 208046 434918 208102
rect 434974 208046 435042 208102
rect 435098 208046 435168 208102
rect 434848 207978 435168 208046
rect 434848 207922 434918 207978
rect 434974 207922 435042 207978
rect 435098 207922 435168 207978
rect 434848 207888 435168 207922
rect 438874 208350 439494 210842
rect 438874 208294 438970 208350
rect 439026 208294 439094 208350
rect 439150 208294 439218 208350
rect 439274 208294 439342 208350
rect 439398 208294 439494 208350
rect 438874 208226 439494 208294
rect 438874 208170 438970 208226
rect 439026 208170 439094 208226
rect 439150 208170 439218 208226
rect 439274 208170 439342 208226
rect 439398 208170 439494 208226
rect 438874 208102 439494 208170
rect 438874 208046 438970 208102
rect 439026 208046 439094 208102
rect 439150 208046 439218 208102
rect 439274 208046 439342 208102
rect 439398 208046 439494 208102
rect 438874 207978 439494 208046
rect 438874 207922 438970 207978
rect 439026 207922 439094 207978
rect 439150 207922 439218 207978
rect 439274 207922 439342 207978
rect 439398 207922 439494 207978
rect 420874 190294 420970 190350
rect 421026 190294 421094 190350
rect 421150 190294 421218 190350
rect 421274 190294 421342 190350
rect 421398 190294 421494 190350
rect 420874 190226 421494 190294
rect 420874 190170 420970 190226
rect 421026 190170 421094 190226
rect 421150 190170 421218 190226
rect 421274 190170 421342 190226
rect 421398 190170 421494 190226
rect 420874 190102 421494 190170
rect 420874 190046 420970 190102
rect 421026 190046 421094 190102
rect 421150 190046 421218 190102
rect 421274 190046 421342 190102
rect 421398 190046 421494 190102
rect 420874 189978 421494 190046
rect 420874 189922 420970 189978
rect 421026 189922 421094 189978
rect 421150 189922 421218 189978
rect 421274 189922 421342 189978
rect 421398 189922 421494 189978
rect 420874 172350 421494 189922
rect 420874 172294 420970 172350
rect 421026 172294 421094 172350
rect 421150 172294 421218 172350
rect 421274 172294 421342 172350
rect 421398 172294 421494 172350
rect 420874 172226 421494 172294
rect 420874 172170 420970 172226
rect 421026 172170 421094 172226
rect 421150 172170 421218 172226
rect 421274 172170 421342 172226
rect 421398 172170 421494 172226
rect 420874 172102 421494 172170
rect 420874 172046 420970 172102
rect 421026 172046 421094 172102
rect 421150 172046 421218 172102
rect 421274 172046 421342 172102
rect 421398 172046 421494 172102
rect 420874 171978 421494 172046
rect 420874 171922 420970 171978
rect 421026 171922 421094 171978
rect 421150 171922 421218 171978
rect 421274 171922 421342 171978
rect 421398 171922 421494 171978
rect 420874 154350 421494 171922
rect 420874 154294 420970 154350
rect 421026 154294 421094 154350
rect 421150 154294 421218 154350
rect 421274 154294 421342 154350
rect 421398 154294 421494 154350
rect 420874 154226 421494 154294
rect 420874 154170 420970 154226
rect 421026 154170 421094 154226
rect 421150 154170 421218 154226
rect 421274 154170 421342 154226
rect 421398 154170 421494 154226
rect 420874 154102 421494 154170
rect 420874 154046 420970 154102
rect 421026 154046 421094 154102
rect 421150 154046 421218 154102
rect 421274 154046 421342 154102
rect 421398 154046 421494 154102
rect 420874 153978 421494 154046
rect 420874 153922 420970 153978
rect 421026 153922 421094 153978
rect 421150 153922 421218 153978
rect 421274 153922 421342 153978
rect 421398 153922 421494 153978
rect 420874 136350 421494 153922
rect 420874 136294 420970 136350
rect 421026 136294 421094 136350
rect 421150 136294 421218 136350
rect 421274 136294 421342 136350
rect 421398 136294 421494 136350
rect 420874 136226 421494 136294
rect 420874 136170 420970 136226
rect 421026 136170 421094 136226
rect 421150 136170 421218 136226
rect 421274 136170 421342 136226
rect 421398 136170 421494 136226
rect 420874 136102 421494 136170
rect 420874 136046 420970 136102
rect 421026 136046 421094 136102
rect 421150 136046 421218 136102
rect 421274 136046 421342 136102
rect 421398 136046 421494 136102
rect 420874 135978 421494 136046
rect 420874 135922 420970 135978
rect 421026 135922 421094 135978
rect 421150 135922 421218 135978
rect 421274 135922 421342 135978
rect 421398 135922 421494 135978
rect 420874 118350 421494 135922
rect 420874 118294 420970 118350
rect 421026 118294 421094 118350
rect 421150 118294 421218 118350
rect 421274 118294 421342 118350
rect 421398 118294 421494 118350
rect 420874 118226 421494 118294
rect 420874 118170 420970 118226
rect 421026 118170 421094 118226
rect 421150 118170 421218 118226
rect 421274 118170 421342 118226
rect 421398 118170 421494 118226
rect 420874 118102 421494 118170
rect 420874 118046 420970 118102
rect 421026 118046 421094 118102
rect 421150 118046 421218 118102
rect 421274 118046 421342 118102
rect 421398 118046 421494 118102
rect 420874 117978 421494 118046
rect 420874 117922 420970 117978
rect 421026 117922 421094 117978
rect 421150 117922 421218 117978
rect 421274 117922 421342 117978
rect 421398 117922 421494 117978
rect 420874 100350 421494 117922
rect 420874 100294 420970 100350
rect 421026 100294 421094 100350
rect 421150 100294 421218 100350
rect 421274 100294 421342 100350
rect 421398 100294 421494 100350
rect 420874 100226 421494 100294
rect 420874 100170 420970 100226
rect 421026 100170 421094 100226
rect 421150 100170 421218 100226
rect 421274 100170 421342 100226
rect 421398 100170 421494 100226
rect 420874 100102 421494 100170
rect 420874 100046 420970 100102
rect 421026 100046 421094 100102
rect 421150 100046 421218 100102
rect 421274 100046 421342 100102
rect 421398 100046 421494 100102
rect 420874 99978 421494 100046
rect 420874 99922 420970 99978
rect 421026 99922 421094 99978
rect 421150 99922 421218 99978
rect 421274 99922 421342 99978
rect 421398 99922 421494 99978
rect 420874 82350 421494 99922
rect 420874 82294 420970 82350
rect 421026 82294 421094 82350
rect 421150 82294 421218 82350
rect 421274 82294 421342 82350
rect 421398 82294 421494 82350
rect 420874 82226 421494 82294
rect 420874 82170 420970 82226
rect 421026 82170 421094 82226
rect 421150 82170 421218 82226
rect 421274 82170 421342 82226
rect 421398 82170 421494 82226
rect 420874 82102 421494 82170
rect 420874 82046 420970 82102
rect 421026 82046 421094 82102
rect 421150 82046 421218 82102
rect 421274 82046 421342 82102
rect 421398 82046 421494 82102
rect 420874 81978 421494 82046
rect 420874 81922 420970 81978
rect 421026 81922 421094 81978
rect 421150 81922 421218 81978
rect 421274 81922 421342 81978
rect 421398 81922 421494 81978
rect 420874 64350 421494 81922
rect 420874 64294 420970 64350
rect 421026 64294 421094 64350
rect 421150 64294 421218 64350
rect 421274 64294 421342 64350
rect 421398 64294 421494 64350
rect 420874 64226 421494 64294
rect 420874 64170 420970 64226
rect 421026 64170 421094 64226
rect 421150 64170 421218 64226
rect 421274 64170 421342 64226
rect 421398 64170 421494 64226
rect 420874 64102 421494 64170
rect 420874 64046 420970 64102
rect 421026 64046 421094 64102
rect 421150 64046 421218 64102
rect 421274 64046 421342 64102
rect 421398 64046 421494 64102
rect 420874 63978 421494 64046
rect 420874 63922 420970 63978
rect 421026 63922 421094 63978
rect 421150 63922 421218 63978
rect 421274 63922 421342 63978
rect 421398 63922 421494 63978
rect 420874 46350 421494 63922
rect 420874 46294 420970 46350
rect 421026 46294 421094 46350
rect 421150 46294 421218 46350
rect 421274 46294 421342 46350
rect 421398 46294 421494 46350
rect 420874 46226 421494 46294
rect 420874 46170 420970 46226
rect 421026 46170 421094 46226
rect 421150 46170 421218 46226
rect 421274 46170 421342 46226
rect 421398 46170 421494 46226
rect 420874 46102 421494 46170
rect 420874 46046 420970 46102
rect 421026 46046 421094 46102
rect 421150 46046 421218 46102
rect 421274 46046 421342 46102
rect 421398 46046 421494 46102
rect 420874 45978 421494 46046
rect 420874 45922 420970 45978
rect 421026 45922 421094 45978
rect 421150 45922 421218 45978
rect 421274 45922 421342 45978
rect 421398 45922 421494 45978
rect 420874 28350 421494 45922
rect 420874 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 421494 28350
rect 420874 28226 421494 28294
rect 420874 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 421494 28226
rect 420874 28102 421494 28170
rect 420874 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 421494 28102
rect 420874 27978 421494 28046
rect 420874 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 421494 27978
rect 420874 10350 421494 27922
rect 420874 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 421494 10350
rect 420874 10226 421494 10294
rect 420874 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 421494 10226
rect 420874 10102 421494 10170
rect 420874 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 421494 10102
rect 420874 9978 421494 10046
rect 420874 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 421494 9978
rect 420874 -1120 421494 9922
rect 420874 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 421494 -1120
rect 420874 -1244 421494 -1176
rect 420874 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 421494 -1244
rect 420874 -1368 421494 -1300
rect 420874 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 421494 -1368
rect 420874 -1492 421494 -1424
rect 420874 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 421494 -1492
rect 420874 -1644 421494 -1548
rect 435154 184350 435774 201020
rect 435154 184294 435250 184350
rect 435306 184294 435374 184350
rect 435430 184294 435498 184350
rect 435554 184294 435622 184350
rect 435678 184294 435774 184350
rect 435154 184226 435774 184294
rect 435154 184170 435250 184226
rect 435306 184170 435374 184226
rect 435430 184170 435498 184226
rect 435554 184170 435622 184226
rect 435678 184170 435774 184226
rect 435154 184102 435774 184170
rect 435154 184046 435250 184102
rect 435306 184046 435374 184102
rect 435430 184046 435498 184102
rect 435554 184046 435622 184102
rect 435678 184046 435774 184102
rect 435154 183978 435774 184046
rect 435154 183922 435250 183978
rect 435306 183922 435374 183978
rect 435430 183922 435498 183978
rect 435554 183922 435622 183978
rect 435678 183922 435774 183978
rect 435154 166350 435774 183922
rect 435154 166294 435250 166350
rect 435306 166294 435374 166350
rect 435430 166294 435498 166350
rect 435554 166294 435622 166350
rect 435678 166294 435774 166350
rect 435154 166226 435774 166294
rect 435154 166170 435250 166226
rect 435306 166170 435374 166226
rect 435430 166170 435498 166226
rect 435554 166170 435622 166226
rect 435678 166170 435774 166226
rect 435154 166102 435774 166170
rect 435154 166046 435250 166102
rect 435306 166046 435374 166102
rect 435430 166046 435498 166102
rect 435554 166046 435622 166102
rect 435678 166046 435774 166102
rect 435154 165978 435774 166046
rect 435154 165922 435250 165978
rect 435306 165922 435374 165978
rect 435430 165922 435498 165978
rect 435554 165922 435622 165978
rect 435678 165922 435774 165978
rect 435154 148350 435774 165922
rect 435154 148294 435250 148350
rect 435306 148294 435374 148350
rect 435430 148294 435498 148350
rect 435554 148294 435622 148350
rect 435678 148294 435774 148350
rect 435154 148226 435774 148294
rect 435154 148170 435250 148226
rect 435306 148170 435374 148226
rect 435430 148170 435498 148226
rect 435554 148170 435622 148226
rect 435678 148170 435774 148226
rect 435154 148102 435774 148170
rect 435154 148046 435250 148102
rect 435306 148046 435374 148102
rect 435430 148046 435498 148102
rect 435554 148046 435622 148102
rect 435678 148046 435774 148102
rect 435154 147978 435774 148046
rect 435154 147922 435250 147978
rect 435306 147922 435374 147978
rect 435430 147922 435498 147978
rect 435554 147922 435622 147978
rect 435678 147922 435774 147978
rect 435154 130350 435774 147922
rect 435154 130294 435250 130350
rect 435306 130294 435374 130350
rect 435430 130294 435498 130350
rect 435554 130294 435622 130350
rect 435678 130294 435774 130350
rect 435154 130226 435774 130294
rect 435154 130170 435250 130226
rect 435306 130170 435374 130226
rect 435430 130170 435498 130226
rect 435554 130170 435622 130226
rect 435678 130170 435774 130226
rect 435154 130102 435774 130170
rect 435154 130046 435250 130102
rect 435306 130046 435374 130102
rect 435430 130046 435498 130102
rect 435554 130046 435622 130102
rect 435678 130046 435774 130102
rect 435154 129978 435774 130046
rect 435154 129922 435250 129978
rect 435306 129922 435374 129978
rect 435430 129922 435498 129978
rect 435554 129922 435622 129978
rect 435678 129922 435774 129978
rect 435154 112350 435774 129922
rect 435154 112294 435250 112350
rect 435306 112294 435374 112350
rect 435430 112294 435498 112350
rect 435554 112294 435622 112350
rect 435678 112294 435774 112350
rect 435154 112226 435774 112294
rect 435154 112170 435250 112226
rect 435306 112170 435374 112226
rect 435430 112170 435498 112226
rect 435554 112170 435622 112226
rect 435678 112170 435774 112226
rect 435154 112102 435774 112170
rect 435154 112046 435250 112102
rect 435306 112046 435374 112102
rect 435430 112046 435498 112102
rect 435554 112046 435622 112102
rect 435678 112046 435774 112102
rect 435154 111978 435774 112046
rect 435154 111922 435250 111978
rect 435306 111922 435374 111978
rect 435430 111922 435498 111978
rect 435554 111922 435622 111978
rect 435678 111922 435774 111978
rect 435154 94350 435774 111922
rect 435154 94294 435250 94350
rect 435306 94294 435374 94350
rect 435430 94294 435498 94350
rect 435554 94294 435622 94350
rect 435678 94294 435774 94350
rect 435154 94226 435774 94294
rect 435154 94170 435250 94226
rect 435306 94170 435374 94226
rect 435430 94170 435498 94226
rect 435554 94170 435622 94226
rect 435678 94170 435774 94226
rect 435154 94102 435774 94170
rect 435154 94046 435250 94102
rect 435306 94046 435374 94102
rect 435430 94046 435498 94102
rect 435554 94046 435622 94102
rect 435678 94046 435774 94102
rect 435154 93978 435774 94046
rect 435154 93922 435250 93978
rect 435306 93922 435374 93978
rect 435430 93922 435498 93978
rect 435554 93922 435622 93978
rect 435678 93922 435774 93978
rect 435154 76350 435774 93922
rect 435154 76294 435250 76350
rect 435306 76294 435374 76350
rect 435430 76294 435498 76350
rect 435554 76294 435622 76350
rect 435678 76294 435774 76350
rect 435154 76226 435774 76294
rect 435154 76170 435250 76226
rect 435306 76170 435374 76226
rect 435430 76170 435498 76226
rect 435554 76170 435622 76226
rect 435678 76170 435774 76226
rect 435154 76102 435774 76170
rect 435154 76046 435250 76102
rect 435306 76046 435374 76102
rect 435430 76046 435498 76102
rect 435554 76046 435622 76102
rect 435678 76046 435774 76102
rect 435154 75978 435774 76046
rect 435154 75922 435250 75978
rect 435306 75922 435374 75978
rect 435430 75922 435498 75978
rect 435554 75922 435622 75978
rect 435678 75922 435774 75978
rect 435154 58350 435774 75922
rect 435154 58294 435250 58350
rect 435306 58294 435374 58350
rect 435430 58294 435498 58350
rect 435554 58294 435622 58350
rect 435678 58294 435774 58350
rect 435154 58226 435774 58294
rect 435154 58170 435250 58226
rect 435306 58170 435374 58226
rect 435430 58170 435498 58226
rect 435554 58170 435622 58226
rect 435678 58170 435774 58226
rect 435154 58102 435774 58170
rect 435154 58046 435250 58102
rect 435306 58046 435374 58102
rect 435430 58046 435498 58102
rect 435554 58046 435622 58102
rect 435678 58046 435774 58102
rect 435154 57978 435774 58046
rect 435154 57922 435250 57978
rect 435306 57922 435374 57978
rect 435430 57922 435498 57978
rect 435554 57922 435622 57978
rect 435678 57922 435774 57978
rect 435154 40350 435774 57922
rect 435154 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 435774 40350
rect 435154 40226 435774 40294
rect 435154 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 435774 40226
rect 435154 40102 435774 40170
rect 435154 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 435774 40102
rect 435154 39978 435774 40046
rect 435154 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 435774 39978
rect 435154 22350 435774 39922
rect 435154 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 435774 22350
rect 435154 22226 435774 22294
rect 435154 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 435774 22226
rect 435154 22102 435774 22170
rect 435154 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 435774 22102
rect 435154 21978 435774 22046
rect 435154 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 435774 21978
rect 435154 4350 435774 21922
rect 435154 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 435774 4350
rect 435154 4226 435774 4294
rect 435154 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 435774 4226
rect 435154 4102 435774 4170
rect 435154 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 435774 4102
rect 435154 3978 435774 4046
rect 435154 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 435774 3978
rect 435154 -160 435774 3922
rect 435154 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 435774 -160
rect 435154 -284 435774 -216
rect 435154 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 435774 -284
rect 435154 -408 435774 -340
rect 435154 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 435774 -408
rect 435154 -532 435774 -464
rect 435154 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 435774 -532
rect 435154 -1644 435774 -588
rect 438874 190350 439494 207922
rect 438874 190294 438970 190350
rect 439026 190294 439094 190350
rect 439150 190294 439218 190350
rect 439274 190294 439342 190350
rect 439398 190294 439494 190350
rect 438874 190226 439494 190294
rect 438874 190170 438970 190226
rect 439026 190170 439094 190226
rect 439150 190170 439218 190226
rect 439274 190170 439342 190226
rect 439398 190170 439494 190226
rect 438874 190102 439494 190170
rect 438874 190046 438970 190102
rect 439026 190046 439094 190102
rect 439150 190046 439218 190102
rect 439274 190046 439342 190102
rect 439398 190046 439494 190102
rect 438874 189978 439494 190046
rect 438874 189922 438970 189978
rect 439026 189922 439094 189978
rect 439150 189922 439218 189978
rect 439274 189922 439342 189978
rect 439398 189922 439494 189978
rect 438874 172350 439494 189922
rect 438874 172294 438970 172350
rect 439026 172294 439094 172350
rect 439150 172294 439218 172350
rect 439274 172294 439342 172350
rect 439398 172294 439494 172350
rect 438874 172226 439494 172294
rect 438874 172170 438970 172226
rect 439026 172170 439094 172226
rect 439150 172170 439218 172226
rect 439274 172170 439342 172226
rect 439398 172170 439494 172226
rect 438874 172102 439494 172170
rect 438874 172046 438970 172102
rect 439026 172046 439094 172102
rect 439150 172046 439218 172102
rect 439274 172046 439342 172102
rect 439398 172046 439494 172102
rect 438874 171978 439494 172046
rect 438874 171922 438970 171978
rect 439026 171922 439094 171978
rect 439150 171922 439218 171978
rect 439274 171922 439342 171978
rect 439398 171922 439494 171978
rect 438874 154350 439494 171922
rect 438874 154294 438970 154350
rect 439026 154294 439094 154350
rect 439150 154294 439218 154350
rect 439274 154294 439342 154350
rect 439398 154294 439494 154350
rect 438874 154226 439494 154294
rect 438874 154170 438970 154226
rect 439026 154170 439094 154226
rect 439150 154170 439218 154226
rect 439274 154170 439342 154226
rect 439398 154170 439494 154226
rect 438874 154102 439494 154170
rect 438874 154046 438970 154102
rect 439026 154046 439094 154102
rect 439150 154046 439218 154102
rect 439274 154046 439342 154102
rect 439398 154046 439494 154102
rect 438874 153978 439494 154046
rect 438874 153922 438970 153978
rect 439026 153922 439094 153978
rect 439150 153922 439218 153978
rect 439274 153922 439342 153978
rect 439398 153922 439494 153978
rect 438874 136350 439494 153922
rect 438874 136294 438970 136350
rect 439026 136294 439094 136350
rect 439150 136294 439218 136350
rect 439274 136294 439342 136350
rect 439398 136294 439494 136350
rect 438874 136226 439494 136294
rect 438874 136170 438970 136226
rect 439026 136170 439094 136226
rect 439150 136170 439218 136226
rect 439274 136170 439342 136226
rect 439398 136170 439494 136226
rect 438874 136102 439494 136170
rect 438874 136046 438970 136102
rect 439026 136046 439094 136102
rect 439150 136046 439218 136102
rect 439274 136046 439342 136102
rect 439398 136046 439494 136102
rect 438874 135978 439494 136046
rect 438874 135922 438970 135978
rect 439026 135922 439094 135978
rect 439150 135922 439218 135978
rect 439274 135922 439342 135978
rect 439398 135922 439494 135978
rect 438874 118350 439494 135922
rect 438874 118294 438970 118350
rect 439026 118294 439094 118350
rect 439150 118294 439218 118350
rect 439274 118294 439342 118350
rect 439398 118294 439494 118350
rect 438874 118226 439494 118294
rect 438874 118170 438970 118226
rect 439026 118170 439094 118226
rect 439150 118170 439218 118226
rect 439274 118170 439342 118226
rect 439398 118170 439494 118226
rect 438874 118102 439494 118170
rect 438874 118046 438970 118102
rect 439026 118046 439094 118102
rect 439150 118046 439218 118102
rect 439274 118046 439342 118102
rect 439398 118046 439494 118102
rect 438874 117978 439494 118046
rect 438874 117922 438970 117978
rect 439026 117922 439094 117978
rect 439150 117922 439218 117978
rect 439274 117922 439342 117978
rect 439398 117922 439494 117978
rect 438874 100350 439494 117922
rect 438874 100294 438970 100350
rect 439026 100294 439094 100350
rect 439150 100294 439218 100350
rect 439274 100294 439342 100350
rect 439398 100294 439494 100350
rect 438874 100226 439494 100294
rect 438874 100170 438970 100226
rect 439026 100170 439094 100226
rect 439150 100170 439218 100226
rect 439274 100170 439342 100226
rect 439398 100170 439494 100226
rect 438874 100102 439494 100170
rect 438874 100046 438970 100102
rect 439026 100046 439094 100102
rect 439150 100046 439218 100102
rect 439274 100046 439342 100102
rect 439398 100046 439494 100102
rect 438874 99978 439494 100046
rect 438874 99922 438970 99978
rect 439026 99922 439094 99978
rect 439150 99922 439218 99978
rect 439274 99922 439342 99978
rect 439398 99922 439494 99978
rect 438874 82350 439494 99922
rect 438874 82294 438970 82350
rect 439026 82294 439094 82350
rect 439150 82294 439218 82350
rect 439274 82294 439342 82350
rect 439398 82294 439494 82350
rect 438874 82226 439494 82294
rect 438874 82170 438970 82226
rect 439026 82170 439094 82226
rect 439150 82170 439218 82226
rect 439274 82170 439342 82226
rect 439398 82170 439494 82226
rect 438874 82102 439494 82170
rect 438874 82046 438970 82102
rect 439026 82046 439094 82102
rect 439150 82046 439218 82102
rect 439274 82046 439342 82102
rect 439398 82046 439494 82102
rect 438874 81978 439494 82046
rect 438874 81922 438970 81978
rect 439026 81922 439094 81978
rect 439150 81922 439218 81978
rect 439274 81922 439342 81978
rect 439398 81922 439494 81978
rect 438874 64350 439494 81922
rect 438874 64294 438970 64350
rect 439026 64294 439094 64350
rect 439150 64294 439218 64350
rect 439274 64294 439342 64350
rect 439398 64294 439494 64350
rect 438874 64226 439494 64294
rect 438874 64170 438970 64226
rect 439026 64170 439094 64226
rect 439150 64170 439218 64226
rect 439274 64170 439342 64226
rect 439398 64170 439494 64226
rect 438874 64102 439494 64170
rect 438874 64046 438970 64102
rect 439026 64046 439094 64102
rect 439150 64046 439218 64102
rect 439274 64046 439342 64102
rect 439398 64046 439494 64102
rect 438874 63978 439494 64046
rect 438874 63922 438970 63978
rect 439026 63922 439094 63978
rect 439150 63922 439218 63978
rect 439274 63922 439342 63978
rect 439398 63922 439494 63978
rect 438874 46350 439494 63922
rect 438874 46294 438970 46350
rect 439026 46294 439094 46350
rect 439150 46294 439218 46350
rect 439274 46294 439342 46350
rect 439398 46294 439494 46350
rect 438874 46226 439494 46294
rect 438874 46170 438970 46226
rect 439026 46170 439094 46226
rect 439150 46170 439218 46226
rect 439274 46170 439342 46226
rect 439398 46170 439494 46226
rect 438874 46102 439494 46170
rect 438874 46046 438970 46102
rect 439026 46046 439094 46102
rect 439150 46046 439218 46102
rect 439274 46046 439342 46102
rect 439398 46046 439494 46102
rect 438874 45978 439494 46046
rect 438874 45922 438970 45978
rect 439026 45922 439094 45978
rect 439150 45922 439218 45978
rect 439274 45922 439342 45978
rect 439398 45922 439494 45978
rect 438874 28350 439494 45922
rect 438874 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 439494 28350
rect 438874 28226 439494 28294
rect 438874 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 439494 28226
rect 438874 28102 439494 28170
rect 438874 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 439494 28102
rect 438874 27978 439494 28046
rect 438874 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 439494 27978
rect 438874 10350 439494 27922
rect 438874 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 439494 10350
rect 438874 10226 439494 10294
rect 438874 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 439494 10226
rect 438874 10102 439494 10170
rect 438874 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 439494 10102
rect 438874 9978 439494 10046
rect 438874 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 439494 9978
rect 438874 -1120 439494 9922
rect 438874 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 439494 -1120
rect 438874 -1244 439494 -1176
rect 438874 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 439494 -1244
rect 438874 -1368 439494 -1300
rect 438874 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 439494 -1368
rect 438874 -1492 439494 -1424
rect 438874 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 439494 -1492
rect 438874 -1644 439494 -1548
rect 453154 202350 453774 210842
rect 453154 202294 453250 202350
rect 453306 202294 453374 202350
rect 453430 202294 453498 202350
rect 453554 202294 453622 202350
rect 453678 202294 453774 202350
rect 453154 202226 453774 202294
rect 453154 202170 453250 202226
rect 453306 202170 453374 202226
rect 453430 202170 453498 202226
rect 453554 202170 453622 202226
rect 453678 202170 453774 202226
rect 453154 202102 453774 202170
rect 453154 202046 453250 202102
rect 453306 202046 453374 202102
rect 453430 202046 453498 202102
rect 453554 202046 453622 202102
rect 453678 202046 453774 202102
rect 453154 201978 453774 202046
rect 453154 201922 453250 201978
rect 453306 201922 453374 201978
rect 453430 201922 453498 201978
rect 453554 201922 453622 201978
rect 453678 201922 453774 201978
rect 453154 184350 453774 201922
rect 453154 184294 453250 184350
rect 453306 184294 453374 184350
rect 453430 184294 453498 184350
rect 453554 184294 453622 184350
rect 453678 184294 453774 184350
rect 453154 184226 453774 184294
rect 453154 184170 453250 184226
rect 453306 184170 453374 184226
rect 453430 184170 453498 184226
rect 453554 184170 453622 184226
rect 453678 184170 453774 184226
rect 453154 184102 453774 184170
rect 453154 184046 453250 184102
rect 453306 184046 453374 184102
rect 453430 184046 453498 184102
rect 453554 184046 453622 184102
rect 453678 184046 453774 184102
rect 453154 183978 453774 184046
rect 453154 183922 453250 183978
rect 453306 183922 453374 183978
rect 453430 183922 453498 183978
rect 453554 183922 453622 183978
rect 453678 183922 453774 183978
rect 453154 166350 453774 183922
rect 453154 166294 453250 166350
rect 453306 166294 453374 166350
rect 453430 166294 453498 166350
rect 453554 166294 453622 166350
rect 453678 166294 453774 166350
rect 453154 166226 453774 166294
rect 453154 166170 453250 166226
rect 453306 166170 453374 166226
rect 453430 166170 453498 166226
rect 453554 166170 453622 166226
rect 453678 166170 453774 166226
rect 453154 166102 453774 166170
rect 453154 166046 453250 166102
rect 453306 166046 453374 166102
rect 453430 166046 453498 166102
rect 453554 166046 453622 166102
rect 453678 166046 453774 166102
rect 453154 165978 453774 166046
rect 453154 165922 453250 165978
rect 453306 165922 453374 165978
rect 453430 165922 453498 165978
rect 453554 165922 453622 165978
rect 453678 165922 453774 165978
rect 453154 148350 453774 165922
rect 453154 148294 453250 148350
rect 453306 148294 453374 148350
rect 453430 148294 453498 148350
rect 453554 148294 453622 148350
rect 453678 148294 453774 148350
rect 453154 148226 453774 148294
rect 453154 148170 453250 148226
rect 453306 148170 453374 148226
rect 453430 148170 453498 148226
rect 453554 148170 453622 148226
rect 453678 148170 453774 148226
rect 453154 148102 453774 148170
rect 453154 148046 453250 148102
rect 453306 148046 453374 148102
rect 453430 148046 453498 148102
rect 453554 148046 453622 148102
rect 453678 148046 453774 148102
rect 453154 147978 453774 148046
rect 453154 147922 453250 147978
rect 453306 147922 453374 147978
rect 453430 147922 453498 147978
rect 453554 147922 453622 147978
rect 453678 147922 453774 147978
rect 453154 130350 453774 147922
rect 453154 130294 453250 130350
rect 453306 130294 453374 130350
rect 453430 130294 453498 130350
rect 453554 130294 453622 130350
rect 453678 130294 453774 130350
rect 453154 130226 453774 130294
rect 453154 130170 453250 130226
rect 453306 130170 453374 130226
rect 453430 130170 453498 130226
rect 453554 130170 453622 130226
rect 453678 130170 453774 130226
rect 453154 130102 453774 130170
rect 453154 130046 453250 130102
rect 453306 130046 453374 130102
rect 453430 130046 453498 130102
rect 453554 130046 453622 130102
rect 453678 130046 453774 130102
rect 453154 129978 453774 130046
rect 453154 129922 453250 129978
rect 453306 129922 453374 129978
rect 453430 129922 453498 129978
rect 453554 129922 453622 129978
rect 453678 129922 453774 129978
rect 453154 112350 453774 129922
rect 453154 112294 453250 112350
rect 453306 112294 453374 112350
rect 453430 112294 453498 112350
rect 453554 112294 453622 112350
rect 453678 112294 453774 112350
rect 453154 112226 453774 112294
rect 453154 112170 453250 112226
rect 453306 112170 453374 112226
rect 453430 112170 453498 112226
rect 453554 112170 453622 112226
rect 453678 112170 453774 112226
rect 453154 112102 453774 112170
rect 453154 112046 453250 112102
rect 453306 112046 453374 112102
rect 453430 112046 453498 112102
rect 453554 112046 453622 112102
rect 453678 112046 453774 112102
rect 453154 111978 453774 112046
rect 453154 111922 453250 111978
rect 453306 111922 453374 111978
rect 453430 111922 453498 111978
rect 453554 111922 453622 111978
rect 453678 111922 453774 111978
rect 453154 94350 453774 111922
rect 453154 94294 453250 94350
rect 453306 94294 453374 94350
rect 453430 94294 453498 94350
rect 453554 94294 453622 94350
rect 453678 94294 453774 94350
rect 453154 94226 453774 94294
rect 453154 94170 453250 94226
rect 453306 94170 453374 94226
rect 453430 94170 453498 94226
rect 453554 94170 453622 94226
rect 453678 94170 453774 94226
rect 453154 94102 453774 94170
rect 453154 94046 453250 94102
rect 453306 94046 453374 94102
rect 453430 94046 453498 94102
rect 453554 94046 453622 94102
rect 453678 94046 453774 94102
rect 453154 93978 453774 94046
rect 453154 93922 453250 93978
rect 453306 93922 453374 93978
rect 453430 93922 453498 93978
rect 453554 93922 453622 93978
rect 453678 93922 453774 93978
rect 453154 76350 453774 93922
rect 453154 76294 453250 76350
rect 453306 76294 453374 76350
rect 453430 76294 453498 76350
rect 453554 76294 453622 76350
rect 453678 76294 453774 76350
rect 453154 76226 453774 76294
rect 453154 76170 453250 76226
rect 453306 76170 453374 76226
rect 453430 76170 453498 76226
rect 453554 76170 453622 76226
rect 453678 76170 453774 76226
rect 453154 76102 453774 76170
rect 453154 76046 453250 76102
rect 453306 76046 453374 76102
rect 453430 76046 453498 76102
rect 453554 76046 453622 76102
rect 453678 76046 453774 76102
rect 453154 75978 453774 76046
rect 453154 75922 453250 75978
rect 453306 75922 453374 75978
rect 453430 75922 453498 75978
rect 453554 75922 453622 75978
rect 453678 75922 453774 75978
rect 453154 58350 453774 75922
rect 453154 58294 453250 58350
rect 453306 58294 453374 58350
rect 453430 58294 453498 58350
rect 453554 58294 453622 58350
rect 453678 58294 453774 58350
rect 453154 58226 453774 58294
rect 453154 58170 453250 58226
rect 453306 58170 453374 58226
rect 453430 58170 453498 58226
rect 453554 58170 453622 58226
rect 453678 58170 453774 58226
rect 453154 58102 453774 58170
rect 453154 58046 453250 58102
rect 453306 58046 453374 58102
rect 453430 58046 453498 58102
rect 453554 58046 453622 58102
rect 453678 58046 453774 58102
rect 453154 57978 453774 58046
rect 453154 57922 453250 57978
rect 453306 57922 453374 57978
rect 453430 57922 453498 57978
rect 453554 57922 453622 57978
rect 453678 57922 453774 57978
rect 453154 40350 453774 57922
rect 453154 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 453774 40350
rect 453154 40226 453774 40294
rect 453154 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 453774 40226
rect 453154 40102 453774 40170
rect 453154 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 453774 40102
rect 453154 39978 453774 40046
rect 453154 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 453774 39978
rect 453154 22350 453774 39922
rect 453154 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 453774 22350
rect 453154 22226 453774 22294
rect 453154 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 453774 22226
rect 453154 22102 453774 22170
rect 453154 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 453774 22102
rect 453154 21978 453774 22046
rect 453154 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 453774 21978
rect 453154 4350 453774 21922
rect 453154 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 453774 4350
rect 453154 4226 453774 4294
rect 453154 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 453774 4226
rect 453154 4102 453774 4170
rect 453154 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 453774 4102
rect 453154 3978 453774 4046
rect 453154 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 453774 3978
rect 453154 -160 453774 3922
rect 453154 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 453774 -160
rect 453154 -284 453774 -216
rect 453154 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 453774 -284
rect 453154 -408 453774 -340
rect 453154 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 453774 -408
rect 453154 -532 453774 -464
rect 453154 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 453774 -532
rect 453154 -1644 453774 -588
rect 456874 208350 457494 210842
rect 456874 208294 456970 208350
rect 457026 208294 457094 208350
rect 457150 208294 457218 208350
rect 457274 208294 457342 208350
rect 457398 208294 457494 208350
rect 456874 208226 457494 208294
rect 456874 208170 456970 208226
rect 457026 208170 457094 208226
rect 457150 208170 457218 208226
rect 457274 208170 457342 208226
rect 457398 208170 457494 208226
rect 456874 208102 457494 208170
rect 456874 208046 456970 208102
rect 457026 208046 457094 208102
rect 457150 208046 457218 208102
rect 457274 208046 457342 208102
rect 457398 208046 457494 208102
rect 456874 207978 457494 208046
rect 456874 207922 456970 207978
rect 457026 207922 457094 207978
rect 457150 207922 457218 207978
rect 457274 207922 457342 207978
rect 457398 207922 457494 207978
rect 456874 190350 457494 207922
rect 465568 208350 465888 208384
rect 465568 208294 465638 208350
rect 465694 208294 465762 208350
rect 465818 208294 465888 208350
rect 465568 208226 465888 208294
rect 465568 208170 465638 208226
rect 465694 208170 465762 208226
rect 465818 208170 465888 208226
rect 465568 208102 465888 208170
rect 465568 208046 465638 208102
rect 465694 208046 465762 208102
rect 465818 208046 465888 208102
rect 465568 207978 465888 208046
rect 465568 207922 465638 207978
rect 465694 207922 465762 207978
rect 465818 207922 465888 207978
rect 465568 207888 465888 207922
rect 456874 190294 456970 190350
rect 457026 190294 457094 190350
rect 457150 190294 457218 190350
rect 457274 190294 457342 190350
rect 457398 190294 457494 190350
rect 456874 190226 457494 190294
rect 456874 190170 456970 190226
rect 457026 190170 457094 190226
rect 457150 190170 457218 190226
rect 457274 190170 457342 190226
rect 457398 190170 457494 190226
rect 456874 190102 457494 190170
rect 456874 190046 456970 190102
rect 457026 190046 457094 190102
rect 457150 190046 457218 190102
rect 457274 190046 457342 190102
rect 457398 190046 457494 190102
rect 456874 189978 457494 190046
rect 456874 189922 456970 189978
rect 457026 189922 457094 189978
rect 457150 189922 457218 189978
rect 457274 189922 457342 189978
rect 457398 189922 457494 189978
rect 456874 172350 457494 189922
rect 456874 172294 456970 172350
rect 457026 172294 457094 172350
rect 457150 172294 457218 172350
rect 457274 172294 457342 172350
rect 457398 172294 457494 172350
rect 456874 172226 457494 172294
rect 456874 172170 456970 172226
rect 457026 172170 457094 172226
rect 457150 172170 457218 172226
rect 457274 172170 457342 172226
rect 457398 172170 457494 172226
rect 456874 172102 457494 172170
rect 456874 172046 456970 172102
rect 457026 172046 457094 172102
rect 457150 172046 457218 172102
rect 457274 172046 457342 172102
rect 457398 172046 457494 172102
rect 456874 171978 457494 172046
rect 456874 171922 456970 171978
rect 457026 171922 457094 171978
rect 457150 171922 457218 171978
rect 457274 171922 457342 171978
rect 457398 171922 457494 171978
rect 456874 154350 457494 171922
rect 456874 154294 456970 154350
rect 457026 154294 457094 154350
rect 457150 154294 457218 154350
rect 457274 154294 457342 154350
rect 457398 154294 457494 154350
rect 456874 154226 457494 154294
rect 456874 154170 456970 154226
rect 457026 154170 457094 154226
rect 457150 154170 457218 154226
rect 457274 154170 457342 154226
rect 457398 154170 457494 154226
rect 456874 154102 457494 154170
rect 456874 154046 456970 154102
rect 457026 154046 457094 154102
rect 457150 154046 457218 154102
rect 457274 154046 457342 154102
rect 457398 154046 457494 154102
rect 456874 153978 457494 154046
rect 456874 153922 456970 153978
rect 457026 153922 457094 153978
rect 457150 153922 457218 153978
rect 457274 153922 457342 153978
rect 457398 153922 457494 153978
rect 456874 136350 457494 153922
rect 456874 136294 456970 136350
rect 457026 136294 457094 136350
rect 457150 136294 457218 136350
rect 457274 136294 457342 136350
rect 457398 136294 457494 136350
rect 456874 136226 457494 136294
rect 456874 136170 456970 136226
rect 457026 136170 457094 136226
rect 457150 136170 457218 136226
rect 457274 136170 457342 136226
rect 457398 136170 457494 136226
rect 456874 136102 457494 136170
rect 456874 136046 456970 136102
rect 457026 136046 457094 136102
rect 457150 136046 457218 136102
rect 457274 136046 457342 136102
rect 457398 136046 457494 136102
rect 456874 135978 457494 136046
rect 456874 135922 456970 135978
rect 457026 135922 457094 135978
rect 457150 135922 457218 135978
rect 457274 135922 457342 135978
rect 457398 135922 457494 135978
rect 456874 118350 457494 135922
rect 456874 118294 456970 118350
rect 457026 118294 457094 118350
rect 457150 118294 457218 118350
rect 457274 118294 457342 118350
rect 457398 118294 457494 118350
rect 456874 118226 457494 118294
rect 456874 118170 456970 118226
rect 457026 118170 457094 118226
rect 457150 118170 457218 118226
rect 457274 118170 457342 118226
rect 457398 118170 457494 118226
rect 456874 118102 457494 118170
rect 456874 118046 456970 118102
rect 457026 118046 457094 118102
rect 457150 118046 457218 118102
rect 457274 118046 457342 118102
rect 457398 118046 457494 118102
rect 456874 117978 457494 118046
rect 456874 117922 456970 117978
rect 457026 117922 457094 117978
rect 457150 117922 457218 117978
rect 457274 117922 457342 117978
rect 457398 117922 457494 117978
rect 456874 100350 457494 117922
rect 456874 100294 456970 100350
rect 457026 100294 457094 100350
rect 457150 100294 457218 100350
rect 457274 100294 457342 100350
rect 457398 100294 457494 100350
rect 456874 100226 457494 100294
rect 456874 100170 456970 100226
rect 457026 100170 457094 100226
rect 457150 100170 457218 100226
rect 457274 100170 457342 100226
rect 457398 100170 457494 100226
rect 456874 100102 457494 100170
rect 456874 100046 456970 100102
rect 457026 100046 457094 100102
rect 457150 100046 457218 100102
rect 457274 100046 457342 100102
rect 457398 100046 457494 100102
rect 456874 99978 457494 100046
rect 456874 99922 456970 99978
rect 457026 99922 457094 99978
rect 457150 99922 457218 99978
rect 457274 99922 457342 99978
rect 457398 99922 457494 99978
rect 456874 82350 457494 99922
rect 456874 82294 456970 82350
rect 457026 82294 457094 82350
rect 457150 82294 457218 82350
rect 457274 82294 457342 82350
rect 457398 82294 457494 82350
rect 456874 82226 457494 82294
rect 456874 82170 456970 82226
rect 457026 82170 457094 82226
rect 457150 82170 457218 82226
rect 457274 82170 457342 82226
rect 457398 82170 457494 82226
rect 456874 82102 457494 82170
rect 456874 82046 456970 82102
rect 457026 82046 457094 82102
rect 457150 82046 457218 82102
rect 457274 82046 457342 82102
rect 457398 82046 457494 82102
rect 456874 81978 457494 82046
rect 456874 81922 456970 81978
rect 457026 81922 457094 81978
rect 457150 81922 457218 81978
rect 457274 81922 457342 81978
rect 457398 81922 457494 81978
rect 456874 64350 457494 81922
rect 456874 64294 456970 64350
rect 457026 64294 457094 64350
rect 457150 64294 457218 64350
rect 457274 64294 457342 64350
rect 457398 64294 457494 64350
rect 456874 64226 457494 64294
rect 456874 64170 456970 64226
rect 457026 64170 457094 64226
rect 457150 64170 457218 64226
rect 457274 64170 457342 64226
rect 457398 64170 457494 64226
rect 456874 64102 457494 64170
rect 456874 64046 456970 64102
rect 457026 64046 457094 64102
rect 457150 64046 457218 64102
rect 457274 64046 457342 64102
rect 457398 64046 457494 64102
rect 456874 63978 457494 64046
rect 456874 63922 456970 63978
rect 457026 63922 457094 63978
rect 457150 63922 457218 63978
rect 457274 63922 457342 63978
rect 457398 63922 457494 63978
rect 456874 46350 457494 63922
rect 456874 46294 456970 46350
rect 457026 46294 457094 46350
rect 457150 46294 457218 46350
rect 457274 46294 457342 46350
rect 457398 46294 457494 46350
rect 456874 46226 457494 46294
rect 456874 46170 456970 46226
rect 457026 46170 457094 46226
rect 457150 46170 457218 46226
rect 457274 46170 457342 46226
rect 457398 46170 457494 46226
rect 456874 46102 457494 46170
rect 456874 46046 456970 46102
rect 457026 46046 457094 46102
rect 457150 46046 457218 46102
rect 457274 46046 457342 46102
rect 457398 46046 457494 46102
rect 456874 45978 457494 46046
rect 456874 45922 456970 45978
rect 457026 45922 457094 45978
rect 457150 45922 457218 45978
rect 457274 45922 457342 45978
rect 457398 45922 457494 45978
rect 456874 28350 457494 45922
rect 456874 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 457494 28350
rect 456874 28226 457494 28294
rect 456874 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 457494 28226
rect 456874 28102 457494 28170
rect 456874 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 457494 28102
rect 456874 27978 457494 28046
rect 456874 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 457494 27978
rect 456874 10350 457494 27922
rect 456874 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 457494 10350
rect 456874 10226 457494 10294
rect 456874 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 457494 10226
rect 456874 10102 457494 10170
rect 456874 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 457494 10102
rect 456874 9978 457494 10046
rect 456874 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 457494 9978
rect 456874 -1120 457494 9922
rect 456874 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 457494 -1120
rect 456874 -1244 457494 -1176
rect 456874 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 457494 -1244
rect 456874 -1368 457494 -1300
rect 456874 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 457494 -1368
rect 456874 -1492 457494 -1424
rect 456874 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 457494 -1492
rect 456874 -1644 457494 -1548
rect 471154 202350 471774 210842
rect 471154 202294 471250 202350
rect 471306 202294 471374 202350
rect 471430 202294 471498 202350
rect 471554 202294 471622 202350
rect 471678 202294 471774 202350
rect 471154 202226 471774 202294
rect 471154 202170 471250 202226
rect 471306 202170 471374 202226
rect 471430 202170 471498 202226
rect 471554 202170 471622 202226
rect 471678 202170 471774 202226
rect 471154 202102 471774 202170
rect 471154 202046 471250 202102
rect 471306 202046 471374 202102
rect 471430 202046 471498 202102
rect 471554 202046 471622 202102
rect 471678 202046 471774 202102
rect 471154 201978 471774 202046
rect 471154 201922 471250 201978
rect 471306 201922 471374 201978
rect 471430 201922 471498 201978
rect 471554 201922 471622 201978
rect 471678 201922 471774 201978
rect 471154 184350 471774 201922
rect 471154 184294 471250 184350
rect 471306 184294 471374 184350
rect 471430 184294 471498 184350
rect 471554 184294 471622 184350
rect 471678 184294 471774 184350
rect 471154 184226 471774 184294
rect 471154 184170 471250 184226
rect 471306 184170 471374 184226
rect 471430 184170 471498 184226
rect 471554 184170 471622 184226
rect 471678 184170 471774 184226
rect 471154 184102 471774 184170
rect 471154 184046 471250 184102
rect 471306 184046 471374 184102
rect 471430 184046 471498 184102
rect 471554 184046 471622 184102
rect 471678 184046 471774 184102
rect 471154 183978 471774 184046
rect 471154 183922 471250 183978
rect 471306 183922 471374 183978
rect 471430 183922 471498 183978
rect 471554 183922 471622 183978
rect 471678 183922 471774 183978
rect 471154 166350 471774 183922
rect 471154 166294 471250 166350
rect 471306 166294 471374 166350
rect 471430 166294 471498 166350
rect 471554 166294 471622 166350
rect 471678 166294 471774 166350
rect 471154 166226 471774 166294
rect 471154 166170 471250 166226
rect 471306 166170 471374 166226
rect 471430 166170 471498 166226
rect 471554 166170 471622 166226
rect 471678 166170 471774 166226
rect 471154 166102 471774 166170
rect 471154 166046 471250 166102
rect 471306 166046 471374 166102
rect 471430 166046 471498 166102
rect 471554 166046 471622 166102
rect 471678 166046 471774 166102
rect 471154 165978 471774 166046
rect 471154 165922 471250 165978
rect 471306 165922 471374 165978
rect 471430 165922 471498 165978
rect 471554 165922 471622 165978
rect 471678 165922 471774 165978
rect 471154 148350 471774 165922
rect 471154 148294 471250 148350
rect 471306 148294 471374 148350
rect 471430 148294 471498 148350
rect 471554 148294 471622 148350
rect 471678 148294 471774 148350
rect 471154 148226 471774 148294
rect 471154 148170 471250 148226
rect 471306 148170 471374 148226
rect 471430 148170 471498 148226
rect 471554 148170 471622 148226
rect 471678 148170 471774 148226
rect 471154 148102 471774 148170
rect 471154 148046 471250 148102
rect 471306 148046 471374 148102
rect 471430 148046 471498 148102
rect 471554 148046 471622 148102
rect 471678 148046 471774 148102
rect 471154 147978 471774 148046
rect 471154 147922 471250 147978
rect 471306 147922 471374 147978
rect 471430 147922 471498 147978
rect 471554 147922 471622 147978
rect 471678 147922 471774 147978
rect 471154 130350 471774 147922
rect 471154 130294 471250 130350
rect 471306 130294 471374 130350
rect 471430 130294 471498 130350
rect 471554 130294 471622 130350
rect 471678 130294 471774 130350
rect 471154 130226 471774 130294
rect 471154 130170 471250 130226
rect 471306 130170 471374 130226
rect 471430 130170 471498 130226
rect 471554 130170 471622 130226
rect 471678 130170 471774 130226
rect 471154 130102 471774 130170
rect 471154 130046 471250 130102
rect 471306 130046 471374 130102
rect 471430 130046 471498 130102
rect 471554 130046 471622 130102
rect 471678 130046 471774 130102
rect 471154 129978 471774 130046
rect 471154 129922 471250 129978
rect 471306 129922 471374 129978
rect 471430 129922 471498 129978
rect 471554 129922 471622 129978
rect 471678 129922 471774 129978
rect 471154 112350 471774 129922
rect 471154 112294 471250 112350
rect 471306 112294 471374 112350
rect 471430 112294 471498 112350
rect 471554 112294 471622 112350
rect 471678 112294 471774 112350
rect 471154 112226 471774 112294
rect 471154 112170 471250 112226
rect 471306 112170 471374 112226
rect 471430 112170 471498 112226
rect 471554 112170 471622 112226
rect 471678 112170 471774 112226
rect 471154 112102 471774 112170
rect 471154 112046 471250 112102
rect 471306 112046 471374 112102
rect 471430 112046 471498 112102
rect 471554 112046 471622 112102
rect 471678 112046 471774 112102
rect 471154 111978 471774 112046
rect 471154 111922 471250 111978
rect 471306 111922 471374 111978
rect 471430 111922 471498 111978
rect 471554 111922 471622 111978
rect 471678 111922 471774 111978
rect 471154 94350 471774 111922
rect 471154 94294 471250 94350
rect 471306 94294 471374 94350
rect 471430 94294 471498 94350
rect 471554 94294 471622 94350
rect 471678 94294 471774 94350
rect 471154 94226 471774 94294
rect 471154 94170 471250 94226
rect 471306 94170 471374 94226
rect 471430 94170 471498 94226
rect 471554 94170 471622 94226
rect 471678 94170 471774 94226
rect 471154 94102 471774 94170
rect 471154 94046 471250 94102
rect 471306 94046 471374 94102
rect 471430 94046 471498 94102
rect 471554 94046 471622 94102
rect 471678 94046 471774 94102
rect 471154 93978 471774 94046
rect 471154 93922 471250 93978
rect 471306 93922 471374 93978
rect 471430 93922 471498 93978
rect 471554 93922 471622 93978
rect 471678 93922 471774 93978
rect 471154 76350 471774 93922
rect 471154 76294 471250 76350
rect 471306 76294 471374 76350
rect 471430 76294 471498 76350
rect 471554 76294 471622 76350
rect 471678 76294 471774 76350
rect 471154 76226 471774 76294
rect 471154 76170 471250 76226
rect 471306 76170 471374 76226
rect 471430 76170 471498 76226
rect 471554 76170 471622 76226
rect 471678 76170 471774 76226
rect 471154 76102 471774 76170
rect 471154 76046 471250 76102
rect 471306 76046 471374 76102
rect 471430 76046 471498 76102
rect 471554 76046 471622 76102
rect 471678 76046 471774 76102
rect 471154 75978 471774 76046
rect 471154 75922 471250 75978
rect 471306 75922 471374 75978
rect 471430 75922 471498 75978
rect 471554 75922 471622 75978
rect 471678 75922 471774 75978
rect 471154 58350 471774 75922
rect 471154 58294 471250 58350
rect 471306 58294 471374 58350
rect 471430 58294 471498 58350
rect 471554 58294 471622 58350
rect 471678 58294 471774 58350
rect 471154 58226 471774 58294
rect 471154 58170 471250 58226
rect 471306 58170 471374 58226
rect 471430 58170 471498 58226
rect 471554 58170 471622 58226
rect 471678 58170 471774 58226
rect 471154 58102 471774 58170
rect 471154 58046 471250 58102
rect 471306 58046 471374 58102
rect 471430 58046 471498 58102
rect 471554 58046 471622 58102
rect 471678 58046 471774 58102
rect 471154 57978 471774 58046
rect 471154 57922 471250 57978
rect 471306 57922 471374 57978
rect 471430 57922 471498 57978
rect 471554 57922 471622 57978
rect 471678 57922 471774 57978
rect 471154 40350 471774 57922
rect 471154 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 471774 40350
rect 471154 40226 471774 40294
rect 471154 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 471774 40226
rect 471154 40102 471774 40170
rect 471154 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 471774 40102
rect 471154 39978 471774 40046
rect 471154 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 471774 39978
rect 471154 22350 471774 39922
rect 471154 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 471774 22350
rect 471154 22226 471774 22294
rect 471154 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 471774 22226
rect 471154 22102 471774 22170
rect 471154 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 471774 22102
rect 471154 21978 471774 22046
rect 471154 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 471774 21978
rect 471154 4350 471774 21922
rect 471154 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 471774 4350
rect 471154 4226 471774 4294
rect 471154 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 471774 4226
rect 471154 4102 471774 4170
rect 471154 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 471774 4102
rect 471154 3978 471774 4046
rect 471154 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 471774 3978
rect 471154 -160 471774 3922
rect 471154 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 471774 -160
rect 471154 -284 471774 -216
rect 471154 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 471774 -284
rect 471154 -408 471774 -340
rect 471154 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 471774 -408
rect 471154 -532 471774 -464
rect 471154 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 471774 -532
rect 471154 -1644 471774 -588
rect 474874 208350 475494 210842
rect 474874 208294 474970 208350
rect 475026 208294 475094 208350
rect 475150 208294 475218 208350
rect 475274 208294 475342 208350
rect 475398 208294 475494 208350
rect 474874 208226 475494 208294
rect 474874 208170 474970 208226
rect 475026 208170 475094 208226
rect 475150 208170 475218 208226
rect 475274 208170 475342 208226
rect 475398 208170 475494 208226
rect 474874 208102 475494 208170
rect 474874 208046 474970 208102
rect 475026 208046 475094 208102
rect 475150 208046 475218 208102
rect 475274 208046 475342 208102
rect 475398 208046 475494 208102
rect 474874 207978 475494 208046
rect 474874 207922 474970 207978
rect 475026 207922 475094 207978
rect 475150 207922 475218 207978
rect 475274 207922 475342 207978
rect 475398 207922 475494 207978
rect 474874 190350 475494 207922
rect 474874 190294 474970 190350
rect 475026 190294 475094 190350
rect 475150 190294 475218 190350
rect 475274 190294 475342 190350
rect 475398 190294 475494 190350
rect 474874 190226 475494 190294
rect 474874 190170 474970 190226
rect 475026 190170 475094 190226
rect 475150 190170 475218 190226
rect 475274 190170 475342 190226
rect 475398 190170 475494 190226
rect 474874 190102 475494 190170
rect 474874 190046 474970 190102
rect 475026 190046 475094 190102
rect 475150 190046 475218 190102
rect 475274 190046 475342 190102
rect 475398 190046 475494 190102
rect 474874 189978 475494 190046
rect 474874 189922 474970 189978
rect 475026 189922 475094 189978
rect 475150 189922 475218 189978
rect 475274 189922 475342 189978
rect 475398 189922 475494 189978
rect 474874 172350 475494 189922
rect 474874 172294 474970 172350
rect 475026 172294 475094 172350
rect 475150 172294 475218 172350
rect 475274 172294 475342 172350
rect 475398 172294 475494 172350
rect 474874 172226 475494 172294
rect 474874 172170 474970 172226
rect 475026 172170 475094 172226
rect 475150 172170 475218 172226
rect 475274 172170 475342 172226
rect 475398 172170 475494 172226
rect 474874 172102 475494 172170
rect 474874 172046 474970 172102
rect 475026 172046 475094 172102
rect 475150 172046 475218 172102
rect 475274 172046 475342 172102
rect 475398 172046 475494 172102
rect 474874 171978 475494 172046
rect 474874 171922 474970 171978
rect 475026 171922 475094 171978
rect 475150 171922 475218 171978
rect 475274 171922 475342 171978
rect 475398 171922 475494 171978
rect 474874 154350 475494 171922
rect 474874 154294 474970 154350
rect 475026 154294 475094 154350
rect 475150 154294 475218 154350
rect 475274 154294 475342 154350
rect 475398 154294 475494 154350
rect 474874 154226 475494 154294
rect 474874 154170 474970 154226
rect 475026 154170 475094 154226
rect 475150 154170 475218 154226
rect 475274 154170 475342 154226
rect 475398 154170 475494 154226
rect 474874 154102 475494 154170
rect 474874 154046 474970 154102
rect 475026 154046 475094 154102
rect 475150 154046 475218 154102
rect 475274 154046 475342 154102
rect 475398 154046 475494 154102
rect 474874 153978 475494 154046
rect 474874 153922 474970 153978
rect 475026 153922 475094 153978
rect 475150 153922 475218 153978
rect 475274 153922 475342 153978
rect 475398 153922 475494 153978
rect 474874 136350 475494 153922
rect 474874 136294 474970 136350
rect 475026 136294 475094 136350
rect 475150 136294 475218 136350
rect 475274 136294 475342 136350
rect 475398 136294 475494 136350
rect 474874 136226 475494 136294
rect 474874 136170 474970 136226
rect 475026 136170 475094 136226
rect 475150 136170 475218 136226
rect 475274 136170 475342 136226
rect 475398 136170 475494 136226
rect 474874 136102 475494 136170
rect 474874 136046 474970 136102
rect 475026 136046 475094 136102
rect 475150 136046 475218 136102
rect 475274 136046 475342 136102
rect 475398 136046 475494 136102
rect 474874 135978 475494 136046
rect 474874 135922 474970 135978
rect 475026 135922 475094 135978
rect 475150 135922 475218 135978
rect 475274 135922 475342 135978
rect 475398 135922 475494 135978
rect 474874 118350 475494 135922
rect 474874 118294 474970 118350
rect 475026 118294 475094 118350
rect 475150 118294 475218 118350
rect 475274 118294 475342 118350
rect 475398 118294 475494 118350
rect 474874 118226 475494 118294
rect 474874 118170 474970 118226
rect 475026 118170 475094 118226
rect 475150 118170 475218 118226
rect 475274 118170 475342 118226
rect 475398 118170 475494 118226
rect 474874 118102 475494 118170
rect 474874 118046 474970 118102
rect 475026 118046 475094 118102
rect 475150 118046 475218 118102
rect 475274 118046 475342 118102
rect 475398 118046 475494 118102
rect 474874 117978 475494 118046
rect 474874 117922 474970 117978
rect 475026 117922 475094 117978
rect 475150 117922 475218 117978
rect 475274 117922 475342 117978
rect 475398 117922 475494 117978
rect 474874 100350 475494 117922
rect 474874 100294 474970 100350
rect 475026 100294 475094 100350
rect 475150 100294 475218 100350
rect 475274 100294 475342 100350
rect 475398 100294 475494 100350
rect 474874 100226 475494 100294
rect 474874 100170 474970 100226
rect 475026 100170 475094 100226
rect 475150 100170 475218 100226
rect 475274 100170 475342 100226
rect 475398 100170 475494 100226
rect 474874 100102 475494 100170
rect 474874 100046 474970 100102
rect 475026 100046 475094 100102
rect 475150 100046 475218 100102
rect 475274 100046 475342 100102
rect 475398 100046 475494 100102
rect 474874 99978 475494 100046
rect 474874 99922 474970 99978
rect 475026 99922 475094 99978
rect 475150 99922 475218 99978
rect 475274 99922 475342 99978
rect 475398 99922 475494 99978
rect 474874 82350 475494 99922
rect 474874 82294 474970 82350
rect 475026 82294 475094 82350
rect 475150 82294 475218 82350
rect 475274 82294 475342 82350
rect 475398 82294 475494 82350
rect 474874 82226 475494 82294
rect 474874 82170 474970 82226
rect 475026 82170 475094 82226
rect 475150 82170 475218 82226
rect 475274 82170 475342 82226
rect 475398 82170 475494 82226
rect 474874 82102 475494 82170
rect 474874 82046 474970 82102
rect 475026 82046 475094 82102
rect 475150 82046 475218 82102
rect 475274 82046 475342 82102
rect 475398 82046 475494 82102
rect 474874 81978 475494 82046
rect 474874 81922 474970 81978
rect 475026 81922 475094 81978
rect 475150 81922 475218 81978
rect 475274 81922 475342 81978
rect 475398 81922 475494 81978
rect 474874 64350 475494 81922
rect 474874 64294 474970 64350
rect 475026 64294 475094 64350
rect 475150 64294 475218 64350
rect 475274 64294 475342 64350
rect 475398 64294 475494 64350
rect 474874 64226 475494 64294
rect 474874 64170 474970 64226
rect 475026 64170 475094 64226
rect 475150 64170 475218 64226
rect 475274 64170 475342 64226
rect 475398 64170 475494 64226
rect 474874 64102 475494 64170
rect 474874 64046 474970 64102
rect 475026 64046 475094 64102
rect 475150 64046 475218 64102
rect 475274 64046 475342 64102
rect 475398 64046 475494 64102
rect 474874 63978 475494 64046
rect 474874 63922 474970 63978
rect 475026 63922 475094 63978
rect 475150 63922 475218 63978
rect 475274 63922 475342 63978
rect 475398 63922 475494 63978
rect 474874 46350 475494 63922
rect 474874 46294 474970 46350
rect 475026 46294 475094 46350
rect 475150 46294 475218 46350
rect 475274 46294 475342 46350
rect 475398 46294 475494 46350
rect 474874 46226 475494 46294
rect 474874 46170 474970 46226
rect 475026 46170 475094 46226
rect 475150 46170 475218 46226
rect 475274 46170 475342 46226
rect 475398 46170 475494 46226
rect 474874 46102 475494 46170
rect 474874 46046 474970 46102
rect 475026 46046 475094 46102
rect 475150 46046 475218 46102
rect 475274 46046 475342 46102
rect 475398 46046 475494 46102
rect 474874 45978 475494 46046
rect 474874 45922 474970 45978
rect 475026 45922 475094 45978
rect 475150 45922 475218 45978
rect 475274 45922 475342 45978
rect 475398 45922 475494 45978
rect 474874 28350 475494 45922
rect 474874 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 475494 28350
rect 474874 28226 475494 28294
rect 474874 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 475494 28226
rect 474874 28102 475494 28170
rect 474874 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 475494 28102
rect 474874 27978 475494 28046
rect 474874 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 475494 27978
rect 474874 10350 475494 27922
rect 474874 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 475494 10350
rect 474874 10226 475494 10294
rect 474874 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 475494 10226
rect 474874 10102 475494 10170
rect 474874 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 475494 10102
rect 474874 9978 475494 10046
rect 474874 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 475494 9978
rect 474874 -1120 475494 9922
rect 474874 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 475494 -1120
rect 474874 -1244 475494 -1176
rect 474874 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 475494 -1244
rect 474874 -1368 475494 -1300
rect 474874 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 475494 -1368
rect 474874 -1492 475494 -1424
rect 474874 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 475494 -1492
rect 474874 -1644 475494 -1548
rect 489154 202350 489774 210842
rect 489154 202294 489250 202350
rect 489306 202294 489374 202350
rect 489430 202294 489498 202350
rect 489554 202294 489622 202350
rect 489678 202294 489774 202350
rect 489154 202226 489774 202294
rect 489154 202170 489250 202226
rect 489306 202170 489374 202226
rect 489430 202170 489498 202226
rect 489554 202170 489622 202226
rect 489678 202170 489774 202226
rect 489154 202102 489774 202170
rect 489154 202046 489250 202102
rect 489306 202046 489374 202102
rect 489430 202046 489498 202102
rect 489554 202046 489622 202102
rect 489678 202046 489774 202102
rect 489154 201978 489774 202046
rect 489154 201922 489250 201978
rect 489306 201922 489374 201978
rect 489430 201922 489498 201978
rect 489554 201922 489622 201978
rect 489678 201922 489774 201978
rect 489154 184350 489774 201922
rect 489154 184294 489250 184350
rect 489306 184294 489374 184350
rect 489430 184294 489498 184350
rect 489554 184294 489622 184350
rect 489678 184294 489774 184350
rect 489154 184226 489774 184294
rect 489154 184170 489250 184226
rect 489306 184170 489374 184226
rect 489430 184170 489498 184226
rect 489554 184170 489622 184226
rect 489678 184170 489774 184226
rect 489154 184102 489774 184170
rect 489154 184046 489250 184102
rect 489306 184046 489374 184102
rect 489430 184046 489498 184102
rect 489554 184046 489622 184102
rect 489678 184046 489774 184102
rect 489154 183978 489774 184046
rect 489154 183922 489250 183978
rect 489306 183922 489374 183978
rect 489430 183922 489498 183978
rect 489554 183922 489622 183978
rect 489678 183922 489774 183978
rect 489154 166350 489774 183922
rect 489154 166294 489250 166350
rect 489306 166294 489374 166350
rect 489430 166294 489498 166350
rect 489554 166294 489622 166350
rect 489678 166294 489774 166350
rect 489154 166226 489774 166294
rect 489154 166170 489250 166226
rect 489306 166170 489374 166226
rect 489430 166170 489498 166226
rect 489554 166170 489622 166226
rect 489678 166170 489774 166226
rect 489154 166102 489774 166170
rect 489154 166046 489250 166102
rect 489306 166046 489374 166102
rect 489430 166046 489498 166102
rect 489554 166046 489622 166102
rect 489678 166046 489774 166102
rect 489154 165978 489774 166046
rect 489154 165922 489250 165978
rect 489306 165922 489374 165978
rect 489430 165922 489498 165978
rect 489554 165922 489622 165978
rect 489678 165922 489774 165978
rect 489154 148350 489774 165922
rect 489154 148294 489250 148350
rect 489306 148294 489374 148350
rect 489430 148294 489498 148350
rect 489554 148294 489622 148350
rect 489678 148294 489774 148350
rect 489154 148226 489774 148294
rect 489154 148170 489250 148226
rect 489306 148170 489374 148226
rect 489430 148170 489498 148226
rect 489554 148170 489622 148226
rect 489678 148170 489774 148226
rect 489154 148102 489774 148170
rect 489154 148046 489250 148102
rect 489306 148046 489374 148102
rect 489430 148046 489498 148102
rect 489554 148046 489622 148102
rect 489678 148046 489774 148102
rect 489154 147978 489774 148046
rect 489154 147922 489250 147978
rect 489306 147922 489374 147978
rect 489430 147922 489498 147978
rect 489554 147922 489622 147978
rect 489678 147922 489774 147978
rect 489154 130350 489774 147922
rect 489154 130294 489250 130350
rect 489306 130294 489374 130350
rect 489430 130294 489498 130350
rect 489554 130294 489622 130350
rect 489678 130294 489774 130350
rect 489154 130226 489774 130294
rect 489154 130170 489250 130226
rect 489306 130170 489374 130226
rect 489430 130170 489498 130226
rect 489554 130170 489622 130226
rect 489678 130170 489774 130226
rect 489154 130102 489774 130170
rect 489154 130046 489250 130102
rect 489306 130046 489374 130102
rect 489430 130046 489498 130102
rect 489554 130046 489622 130102
rect 489678 130046 489774 130102
rect 489154 129978 489774 130046
rect 489154 129922 489250 129978
rect 489306 129922 489374 129978
rect 489430 129922 489498 129978
rect 489554 129922 489622 129978
rect 489678 129922 489774 129978
rect 489154 112350 489774 129922
rect 489154 112294 489250 112350
rect 489306 112294 489374 112350
rect 489430 112294 489498 112350
rect 489554 112294 489622 112350
rect 489678 112294 489774 112350
rect 489154 112226 489774 112294
rect 489154 112170 489250 112226
rect 489306 112170 489374 112226
rect 489430 112170 489498 112226
rect 489554 112170 489622 112226
rect 489678 112170 489774 112226
rect 489154 112102 489774 112170
rect 489154 112046 489250 112102
rect 489306 112046 489374 112102
rect 489430 112046 489498 112102
rect 489554 112046 489622 112102
rect 489678 112046 489774 112102
rect 489154 111978 489774 112046
rect 489154 111922 489250 111978
rect 489306 111922 489374 111978
rect 489430 111922 489498 111978
rect 489554 111922 489622 111978
rect 489678 111922 489774 111978
rect 489154 94350 489774 111922
rect 489154 94294 489250 94350
rect 489306 94294 489374 94350
rect 489430 94294 489498 94350
rect 489554 94294 489622 94350
rect 489678 94294 489774 94350
rect 489154 94226 489774 94294
rect 489154 94170 489250 94226
rect 489306 94170 489374 94226
rect 489430 94170 489498 94226
rect 489554 94170 489622 94226
rect 489678 94170 489774 94226
rect 489154 94102 489774 94170
rect 489154 94046 489250 94102
rect 489306 94046 489374 94102
rect 489430 94046 489498 94102
rect 489554 94046 489622 94102
rect 489678 94046 489774 94102
rect 489154 93978 489774 94046
rect 489154 93922 489250 93978
rect 489306 93922 489374 93978
rect 489430 93922 489498 93978
rect 489554 93922 489622 93978
rect 489678 93922 489774 93978
rect 489154 76350 489774 93922
rect 489154 76294 489250 76350
rect 489306 76294 489374 76350
rect 489430 76294 489498 76350
rect 489554 76294 489622 76350
rect 489678 76294 489774 76350
rect 489154 76226 489774 76294
rect 489154 76170 489250 76226
rect 489306 76170 489374 76226
rect 489430 76170 489498 76226
rect 489554 76170 489622 76226
rect 489678 76170 489774 76226
rect 489154 76102 489774 76170
rect 489154 76046 489250 76102
rect 489306 76046 489374 76102
rect 489430 76046 489498 76102
rect 489554 76046 489622 76102
rect 489678 76046 489774 76102
rect 489154 75978 489774 76046
rect 489154 75922 489250 75978
rect 489306 75922 489374 75978
rect 489430 75922 489498 75978
rect 489554 75922 489622 75978
rect 489678 75922 489774 75978
rect 489154 58350 489774 75922
rect 489154 58294 489250 58350
rect 489306 58294 489374 58350
rect 489430 58294 489498 58350
rect 489554 58294 489622 58350
rect 489678 58294 489774 58350
rect 489154 58226 489774 58294
rect 489154 58170 489250 58226
rect 489306 58170 489374 58226
rect 489430 58170 489498 58226
rect 489554 58170 489622 58226
rect 489678 58170 489774 58226
rect 489154 58102 489774 58170
rect 489154 58046 489250 58102
rect 489306 58046 489374 58102
rect 489430 58046 489498 58102
rect 489554 58046 489622 58102
rect 489678 58046 489774 58102
rect 489154 57978 489774 58046
rect 489154 57922 489250 57978
rect 489306 57922 489374 57978
rect 489430 57922 489498 57978
rect 489554 57922 489622 57978
rect 489678 57922 489774 57978
rect 489154 40350 489774 57922
rect 489154 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 489774 40350
rect 489154 40226 489774 40294
rect 489154 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 489774 40226
rect 489154 40102 489774 40170
rect 489154 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 489774 40102
rect 489154 39978 489774 40046
rect 489154 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 489774 39978
rect 489154 22350 489774 39922
rect 489154 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 489774 22350
rect 489154 22226 489774 22294
rect 489154 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 489774 22226
rect 489154 22102 489774 22170
rect 489154 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 489774 22102
rect 489154 21978 489774 22046
rect 489154 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 489774 21978
rect 489154 4350 489774 21922
rect 489154 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 489774 4350
rect 489154 4226 489774 4294
rect 489154 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 489774 4226
rect 489154 4102 489774 4170
rect 489154 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 489774 4102
rect 489154 3978 489774 4046
rect 489154 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 489774 3978
rect 489154 -160 489774 3922
rect 489154 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 489774 -160
rect 489154 -284 489774 -216
rect 489154 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 489774 -284
rect 489154 -408 489774 -340
rect 489154 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 489774 -408
rect 489154 -532 489774 -464
rect 489154 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 489774 -532
rect 489154 -1644 489774 -588
rect 492874 208350 493494 210842
rect 492874 208294 492970 208350
rect 493026 208294 493094 208350
rect 493150 208294 493218 208350
rect 493274 208294 493342 208350
rect 493398 208294 493494 208350
rect 492874 208226 493494 208294
rect 492874 208170 492970 208226
rect 493026 208170 493094 208226
rect 493150 208170 493218 208226
rect 493274 208170 493342 208226
rect 493398 208170 493494 208226
rect 492874 208102 493494 208170
rect 492874 208046 492970 208102
rect 493026 208046 493094 208102
rect 493150 208046 493218 208102
rect 493274 208046 493342 208102
rect 493398 208046 493494 208102
rect 492874 207978 493494 208046
rect 492874 207922 492970 207978
rect 493026 207922 493094 207978
rect 493150 207922 493218 207978
rect 493274 207922 493342 207978
rect 493398 207922 493494 207978
rect 492874 190350 493494 207922
rect 496288 208350 496608 208384
rect 496288 208294 496358 208350
rect 496414 208294 496482 208350
rect 496538 208294 496608 208350
rect 496288 208226 496608 208294
rect 496288 208170 496358 208226
rect 496414 208170 496482 208226
rect 496538 208170 496608 208226
rect 496288 208102 496608 208170
rect 496288 208046 496358 208102
rect 496414 208046 496482 208102
rect 496538 208046 496608 208102
rect 496288 207978 496608 208046
rect 496288 207922 496358 207978
rect 496414 207922 496482 207978
rect 496538 207922 496608 207978
rect 496288 207888 496608 207922
rect 492874 190294 492970 190350
rect 493026 190294 493094 190350
rect 493150 190294 493218 190350
rect 493274 190294 493342 190350
rect 493398 190294 493494 190350
rect 492874 190226 493494 190294
rect 492874 190170 492970 190226
rect 493026 190170 493094 190226
rect 493150 190170 493218 190226
rect 493274 190170 493342 190226
rect 493398 190170 493494 190226
rect 492874 190102 493494 190170
rect 492874 190046 492970 190102
rect 493026 190046 493094 190102
rect 493150 190046 493218 190102
rect 493274 190046 493342 190102
rect 493398 190046 493494 190102
rect 492874 189978 493494 190046
rect 492874 189922 492970 189978
rect 493026 189922 493094 189978
rect 493150 189922 493218 189978
rect 493274 189922 493342 189978
rect 493398 189922 493494 189978
rect 492874 172350 493494 189922
rect 492874 172294 492970 172350
rect 493026 172294 493094 172350
rect 493150 172294 493218 172350
rect 493274 172294 493342 172350
rect 493398 172294 493494 172350
rect 492874 172226 493494 172294
rect 492874 172170 492970 172226
rect 493026 172170 493094 172226
rect 493150 172170 493218 172226
rect 493274 172170 493342 172226
rect 493398 172170 493494 172226
rect 492874 172102 493494 172170
rect 492874 172046 492970 172102
rect 493026 172046 493094 172102
rect 493150 172046 493218 172102
rect 493274 172046 493342 172102
rect 493398 172046 493494 172102
rect 492874 171978 493494 172046
rect 492874 171922 492970 171978
rect 493026 171922 493094 171978
rect 493150 171922 493218 171978
rect 493274 171922 493342 171978
rect 493398 171922 493494 171978
rect 492874 154350 493494 171922
rect 492874 154294 492970 154350
rect 493026 154294 493094 154350
rect 493150 154294 493218 154350
rect 493274 154294 493342 154350
rect 493398 154294 493494 154350
rect 492874 154226 493494 154294
rect 492874 154170 492970 154226
rect 493026 154170 493094 154226
rect 493150 154170 493218 154226
rect 493274 154170 493342 154226
rect 493398 154170 493494 154226
rect 492874 154102 493494 154170
rect 492874 154046 492970 154102
rect 493026 154046 493094 154102
rect 493150 154046 493218 154102
rect 493274 154046 493342 154102
rect 493398 154046 493494 154102
rect 492874 153978 493494 154046
rect 492874 153922 492970 153978
rect 493026 153922 493094 153978
rect 493150 153922 493218 153978
rect 493274 153922 493342 153978
rect 493398 153922 493494 153978
rect 492874 136350 493494 153922
rect 492874 136294 492970 136350
rect 493026 136294 493094 136350
rect 493150 136294 493218 136350
rect 493274 136294 493342 136350
rect 493398 136294 493494 136350
rect 492874 136226 493494 136294
rect 492874 136170 492970 136226
rect 493026 136170 493094 136226
rect 493150 136170 493218 136226
rect 493274 136170 493342 136226
rect 493398 136170 493494 136226
rect 492874 136102 493494 136170
rect 492874 136046 492970 136102
rect 493026 136046 493094 136102
rect 493150 136046 493218 136102
rect 493274 136046 493342 136102
rect 493398 136046 493494 136102
rect 492874 135978 493494 136046
rect 492874 135922 492970 135978
rect 493026 135922 493094 135978
rect 493150 135922 493218 135978
rect 493274 135922 493342 135978
rect 493398 135922 493494 135978
rect 492874 118350 493494 135922
rect 492874 118294 492970 118350
rect 493026 118294 493094 118350
rect 493150 118294 493218 118350
rect 493274 118294 493342 118350
rect 493398 118294 493494 118350
rect 492874 118226 493494 118294
rect 492874 118170 492970 118226
rect 493026 118170 493094 118226
rect 493150 118170 493218 118226
rect 493274 118170 493342 118226
rect 493398 118170 493494 118226
rect 492874 118102 493494 118170
rect 492874 118046 492970 118102
rect 493026 118046 493094 118102
rect 493150 118046 493218 118102
rect 493274 118046 493342 118102
rect 493398 118046 493494 118102
rect 492874 117978 493494 118046
rect 492874 117922 492970 117978
rect 493026 117922 493094 117978
rect 493150 117922 493218 117978
rect 493274 117922 493342 117978
rect 493398 117922 493494 117978
rect 492874 100350 493494 117922
rect 492874 100294 492970 100350
rect 493026 100294 493094 100350
rect 493150 100294 493218 100350
rect 493274 100294 493342 100350
rect 493398 100294 493494 100350
rect 492874 100226 493494 100294
rect 492874 100170 492970 100226
rect 493026 100170 493094 100226
rect 493150 100170 493218 100226
rect 493274 100170 493342 100226
rect 493398 100170 493494 100226
rect 492874 100102 493494 100170
rect 492874 100046 492970 100102
rect 493026 100046 493094 100102
rect 493150 100046 493218 100102
rect 493274 100046 493342 100102
rect 493398 100046 493494 100102
rect 492874 99978 493494 100046
rect 492874 99922 492970 99978
rect 493026 99922 493094 99978
rect 493150 99922 493218 99978
rect 493274 99922 493342 99978
rect 493398 99922 493494 99978
rect 492874 82350 493494 99922
rect 492874 82294 492970 82350
rect 493026 82294 493094 82350
rect 493150 82294 493218 82350
rect 493274 82294 493342 82350
rect 493398 82294 493494 82350
rect 492874 82226 493494 82294
rect 492874 82170 492970 82226
rect 493026 82170 493094 82226
rect 493150 82170 493218 82226
rect 493274 82170 493342 82226
rect 493398 82170 493494 82226
rect 492874 82102 493494 82170
rect 492874 82046 492970 82102
rect 493026 82046 493094 82102
rect 493150 82046 493218 82102
rect 493274 82046 493342 82102
rect 493398 82046 493494 82102
rect 492874 81978 493494 82046
rect 492874 81922 492970 81978
rect 493026 81922 493094 81978
rect 493150 81922 493218 81978
rect 493274 81922 493342 81978
rect 493398 81922 493494 81978
rect 492874 64350 493494 81922
rect 492874 64294 492970 64350
rect 493026 64294 493094 64350
rect 493150 64294 493218 64350
rect 493274 64294 493342 64350
rect 493398 64294 493494 64350
rect 492874 64226 493494 64294
rect 492874 64170 492970 64226
rect 493026 64170 493094 64226
rect 493150 64170 493218 64226
rect 493274 64170 493342 64226
rect 493398 64170 493494 64226
rect 492874 64102 493494 64170
rect 492874 64046 492970 64102
rect 493026 64046 493094 64102
rect 493150 64046 493218 64102
rect 493274 64046 493342 64102
rect 493398 64046 493494 64102
rect 492874 63978 493494 64046
rect 492874 63922 492970 63978
rect 493026 63922 493094 63978
rect 493150 63922 493218 63978
rect 493274 63922 493342 63978
rect 493398 63922 493494 63978
rect 492874 46350 493494 63922
rect 492874 46294 492970 46350
rect 493026 46294 493094 46350
rect 493150 46294 493218 46350
rect 493274 46294 493342 46350
rect 493398 46294 493494 46350
rect 492874 46226 493494 46294
rect 492874 46170 492970 46226
rect 493026 46170 493094 46226
rect 493150 46170 493218 46226
rect 493274 46170 493342 46226
rect 493398 46170 493494 46226
rect 492874 46102 493494 46170
rect 492874 46046 492970 46102
rect 493026 46046 493094 46102
rect 493150 46046 493218 46102
rect 493274 46046 493342 46102
rect 493398 46046 493494 46102
rect 492874 45978 493494 46046
rect 492874 45922 492970 45978
rect 493026 45922 493094 45978
rect 493150 45922 493218 45978
rect 493274 45922 493342 45978
rect 493398 45922 493494 45978
rect 492874 28350 493494 45922
rect 492874 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 493494 28350
rect 492874 28226 493494 28294
rect 492874 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 493494 28226
rect 492874 28102 493494 28170
rect 492874 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 493494 28102
rect 492874 27978 493494 28046
rect 492874 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 493494 27978
rect 492874 10350 493494 27922
rect 492874 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 493494 10350
rect 492874 10226 493494 10294
rect 492874 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 493494 10226
rect 492874 10102 493494 10170
rect 492874 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 493494 10102
rect 492874 9978 493494 10046
rect 492874 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 493494 9978
rect 492874 -1120 493494 9922
rect 492874 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 493494 -1120
rect 492874 -1244 493494 -1176
rect 492874 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 493494 -1244
rect 492874 -1368 493494 -1300
rect 492874 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 493494 -1368
rect 492874 -1492 493494 -1424
rect 492874 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 493494 -1492
rect 492874 -1644 493494 -1548
rect 507154 202350 507774 219922
rect 507154 202294 507250 202350
rect 507306 202294 507374 202350
rect 507430 202294 507498 202350
rect 507554 202294 507622 202350
rect 507678 202294 507774 202350
rect 507154 202226 507774 202294
rect 507154 202170 507250 202226
rect 507306 202170 507374 202226
rect 507430 202170 507498 202226
rect 507554 202170 507622 202226
rect 507678 202170 507774 202226
rect 507154 202102 507774 202170
rect 507154 202046 507250 202102
rect 507306 202046 507374 202102
rect 507430 202046 507498 202102
rect 507554 202046 507622 202102
rect 507678 202046 507774 202102
rect 507154 201978 507774 202046
rect 507154 201922 507250 201978
rect 507306 201922 507374 201978
rect 507430 201922 507498 201978
rect 507554 201922 507622 201978
rect 507678 201922 507774 201978
rect 507154 184350 507774 201922
rect 507154 184294 507250 184350
rect 507306 184294 507374 184350
rect 507430 184294 507498 184350
rect 507554 184294 507622 184350
rect 507678 184294 507774 184350
rect 507154 184226 507774 184294
rect 507154 184170 507250 184226
rect 507306 184170 507374 184226
rect 507430 184170 507498 184226
rect 507554 184170 507622 184226
rect 507678 184170 507774 184226
rect 507154 184102 507774 184170
rect 507154 184046 507250 184102
rect 507306 184046 507374 184102
rect 507430 184046 507498 184102
rect 507554 184046 507622 184102
rect 507678 184046 507774 184102
rect 507154 183978 507774 184046
rect 507154 183922 507250 183978
rect 507306 183922 507374 183978
rect 507430 183922 507498 183978
rect 507554 183922 507622 183978
rect 507678 183922 507774 183978
rect 507154 166350 507774 183922
rect 507154 166294 507250 166350
rect 507306 166294 507374 166350
rect 507430 166294 507498 166350
rect 507554 166294 507622 166350
rect 507678 166294 507774 166350
rect 507154 166226 507774 166294
rect 507154 166170 507250 166226
rect 507306 166170 507374 166226
rect 507430 166170 507498 166226
rect 507554 166170 507622 166226
rect 507678 166170 507774 166226
rect 507154 166102 507774 166170
rect 507154 166046 507250 166102
rect 507306 166046 507374 166102
rect 507430 166046 507498 166102
rect 507554 166046 507622 166102
rect 507678 166046 507774 166102
rect 507154 165978 507774 166046
rect 507154 165922 507250 165978
rect 507306 165922 507374 165978
rect 507430 165922 507498 165978
rect 507554 165922 507622 165978
rect 507678 165922 507774 165978
rect 507154 148350 507774 165922
rect 507154 148294 507250 148350
rect 507306 148294 507374 148350
rect 507430 148294 507498 148350
rect 507554 148294 507622 148350
rect 507678 148294 507774 148350
rect 507154 148226 507774 148294
rect 507154 148170 507250 148226
rect 507306 148170 507374 148226
rect 507430 148170 507498 148226
rect 507554 148170 507622 148226
rect 507678 148170 507774 148226
rect 507154 148102 507774 148170
rect 507154 148046 507250 148102
rect 507306 148046 507374 148102
rect 507430 148046 507498 148102
rect 507554 148046 507622 148102
rect 507678 148046 507774 148102
rect 507154 147978 507774 148046
rect 507154 147922 507250 147978
rect 507306 147922 507374 147978
rect 507430 147922 507498 147978
rect 507554 147922 507622 147978
rect 507678 147922 507774 147978
rect 507154 130350 507774 147922
rect 507154 130294 507250 130350
rect 507306 130294 507374 130350
rect 507430 130294 507498 130350
rect 507554 130294 507622 130350
rect 507678 130294 507774 130350
rect 507154 130226 507774 130294
rect 507154 130170 507250 130226
rect 507306 130170 507374 130226
rect 507430 130170 507498 130226
rect 507554 130170 507622 130226
rect 507678 130170 507774 130226
rect 507154 130102 507774 130170
rect 507154 130046 507250 130102
rect 507306 130046 507374 130102
rect 507430 130046 507498 130102
rect 507554 130046 507622 130102
rect 507678 130046 507774 130102
rect 507154 129978 507774 130046
rect 507154 129922 507250 129978
rect 507306 129922 507374 129978
rect 507430 129922 507498 129978
rect 507554 129922 507622 129978
rect 507678 129922 507774 129978
rect 507154 112350 507774 129922
rect 507154 112294 507250 112350
rect 507306 112294 507374 112350
rect 507430 112294 507498 112350
rect 507554 112294 507622 112350
rect 507678 112294 507774 112350
rect 507154 112226 507774 112294
rect 507154 112170 507250 112226
rect 507306 112170 507374 112226
rect 507430 112170 507498 112226
rect 507554 112170 507622 112226
rect 507678 112170 507774 112226
rect 507154 112102 507774 112170
rect 507154 112046 507250 112102
rect 507306 112046 507374 112102
rect 507430 112046 507498 112102
rect 507554 112046 507622 112102
rect 507678 112046 507774 112102
rect 507154 111978 507774 112046
rect 507154 111922 507250 111978
rect 507306 111922 507374 111978
rect 507430 111922 507498 111978
rect 507554 111922 507622 111978
rect 507678 111922 507774 111978
rect 507154 94350 507774 111922
rect 507154 94294 507250 94350
rect 507306 94294 507374 94350
rect 507430 94294 507498 94350
rect 507554 94294 507622 94350
rect 507678 94294 507774 94350
rect 507154 94226 507774 94294
rect 507154 94170 507250 94226
rect 507306 94170 507374 94226
rect 507430 94170 507498 94226
rect 507554 94170 507622 94226
rect 507678 94170 507774 94226
rect 507154 94102 507774 94170
rect 507154 94046 507250 94102
rect 507306 94046 507374 94102
rect 507430 94046 507498 94102
rect 507554 94046 507622 94102
rect 507678 94046 507774 94102
rect 507154 93978 507774 94046
rect 507154 93922 507250 93978
rect 507306 93922 507374 93978
rect 507430 93922 507498 93978
rect 507554 93922 507622 93978
rect 507678 93922 507774 93978
rect 507154 76350 507774 93922
rect 507154 76294 507250 76350
rect 507306 76294 507374 76350
rect 507430 76294 507498 76350
rect 507554 76294 507622 76350
rect 507678 76294 507774 76350
rect 507154 76226 507774 76294
rect 507154 76170 507250 76226
rect 507306 76170 507374 76226
rect 507430 76170 507498 76226
rect 507554 76170 507622 76226
rect 507678 76170 507774 76226
rect 507154 76102 507774 76170
rect 507154 76046 507250 76102
rect 507306 76046 507374 76102
rect 507430 76046 507498 76102
rect 507554 76046 507622 76102
rect 507678 76046 507774 76102
rect 507154 75978 507774 76046
rect 507154 75922 507250 75978
rect 507306 75922 507374 75978
rect 507430 75922 507498 75978
rect 507554 75922 507622 75978
rect 507678 75922 507774 75978
rect 507154 58350 507774 75922
rect 507154 58294 507250 58350
rect 507306 58294 507374 58350
rect 507430 58294 507498 58350
rect 507554 58294 507622 58350
rect 507678 58294 507774 58350
rect 507154 58226 507774 58294
rect 507154 58170 507250 58226
rect 507306 58170 507374 58226
rect 507430 58170 507498 58226
rect 507554 58170 507622 58226
rect 507678 58170 507774 58226
rect 507154 58102 507774 58170
rect 507154 58046 507250 58102
rect 507306 58046 507374 58102
rect 507430 58046 507498 58102
rect 507554 58046 507622 58102
rect 507678 58046 507774 58102
rect 507154 57978 507774 58046
rect 507154 57922 507250 57978
rect 507306 57922 507374 57978
rect 507430 57922 507498 57978
rect 507554 57922 507622 57978
rect 507678 57922 507774 57978
rect 507154 40350 507774 57922
rect 507154 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 507774 40350
rect 507154 40226 507774 40294
rect 507154 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 507774 40226
rect 507154 40102 507774 40170
rect 507154 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 507774 40102
rect 507154 39978 507774 40046
rect 507154 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 507774 39978
rect 507154 22350 507774 39922
rect 507154 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 507774 22350
rect 507154 22226 507774 22294
rect 507154 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 507774 22226
rect 507154 22102 507774 22170
rect 507154 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 507774 22102
rect 507154 21978 507774 22046
rect 507154 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 507774 21978
rect 507154 4350 507774 21922
rect 507154 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 507774 4350
rect 507154 4226 507774 4294
rect 507154 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 507774 4226
rect 507154 4102 507774 4170
rect 507154 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 507774 4102
rect 507154 3978 507774 4046
rect 507154 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 507774 3978
rect 507154 -160 507774 3922
rect 507154 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 507774 -160
rect 507154 -284 507774 -216
rect 507154 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 507774 -284
rect 507154 -408 507774 -340
rect 507154 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 507774 -408
rect 507154 -532 507774 -464
rect 507154 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 507774 -532
rect 507154 -1644 507774 -588
rect 510874 598172 511494 598268
rect 510874 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 511494 598172
rect 510874 598048 511494 598116
rect 510874 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 511494 598048
rect 510874 597924 511494 597992
rect 510874 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 511494 597924
rect 510874 597800 511494 597868
rect 510874 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 511494 597800
rect 510874 586350 511494 597744
rect 510874 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 511494 586350
rect 510874 586226 511494 586294
rect 510874 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 511494 586226
rect 510874 586102 511494 586170
rect 510874 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 511494 586102
rect 510874 585978 511494 586046
rect 510874 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 511494 585978
rect 510874 568350 511494 585922
rect 510874 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 511494 568350
rect 510874 568226 511494 568294
rect 510874 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 511494 568226
rect 510874 568102 511494 568170
rect 510874 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 511494 568102
rect 510874 567978 511494 568046
rect 510874 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 511494 567978
rect 510874 550350 511494 567922
rect 510874 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 511494 550350
rect 510874 550226 511494 550294
rect 510874 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 511494 550226
rect 510874 550102 511494 550170
rect 510874 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 511494 550102
rect 510874 549978 511494 550046
rect 510874 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 511494 549978
rect 510874 532350 511494 549922
rect 510874 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 511494 532350
rect 510874 532226 511494 532294
rect 510874 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 511494 532226
rect 510874 532102 511494 532170
rect 510874 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 511494 532102
rect 510874 531978 511494 532046
rect 510874 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 511494 531978
rect 510874 514350 511494 531922
rect 510874 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 511494 514350
rect 510874 514226 511494 514294
rect 510874 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 511494 514226
rect 510874 514102 511494 514170
rect 510874 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 511494 514102
rect 510874 513978 511494 514046
rect 510874 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 511494 513978
rect 510874 496350 511494 513922
rect 510874 496294 510970 496350
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 511494 496350
rect 510874 496226 511494 496294
rect 510874 496170 510970 496226
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 511494 496226
rect 510874 496102 511494 496170
rect 510874 496046 510970 496102
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 511494 496102
rect 510874 495978 511494 496046
rect 510874 495922 510970 495978
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 511494 495978
rect 510874 478350 511494 495922
rect 510874 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 511494 478350
rect 510874 478226 511494 478294
rect 510874 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 511494 478226
rect 510874 478102 511494 478170
rect 510874 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 511494 478102
rect 510874 477978 511494 478046
rect 510874 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 511494 477978
rect 510874 460350 511494 477922
rect 510874 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 511494 460350
rect 510874 460226 511494 460294
rect 510874 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 511494 460226
rect 510874 460102 511494 460170
rect 510874 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 511494 460102
rect 510874 459978 511494 460046
rect 510874 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 511494 459978
rect 510874 442350 511494 459922
rect 510874 442294 510970 442350
rect 511026 442294 511094 442350
rect 511150 442294 511218 442350
rect 511274 442294 511342 442350
rect 511398 442294 511494 442350
rect 510874 442226 511494 442294
rect 510874 442170 510970 442226
rect 511026 442170 511094 442226
rect 511150 442170 511218 442226
rect 511274 442170 511342 442226
rect 511398 442170 511494 442226
rect 510874 442102 511494 442170
rect 510874 442046 510970 442102
rect 511026 442046 511094 442102
rect 511150 442046 511218 442102
rect 511274 442046 511342 442102
rect 511398 442046 511494 442102
rect 510874 441978 511494 442046
rect 510874 441922 510970 441978
rect 511026 441922 511094 441978
rect 511150 441922 511218 441978
rect 511274 441922 511342 441978
rect 511398 441922 511494 441978
rect 510874 424350 511494 441922
rect 510874 424294 510970 424350
rect 511026 424294 511094 424350
rect 511150 424294 511218 424350
rect 511274 424294 511342 424350
rect 511398 424294 511494 424350
rect 510874 424226 511494 424294
rect 510874 424170 510970 424226
rect 511026 424170 511094 424226
rect 511150 424170 511218 424226
rect 511274 424170 511342 424226
rect 511398 424170 511494 424226
rect 510874 424102 511494 424170
rect 510874 424046 510970 424102
rect 511026 424046 511094 424102
rect 511150 424046 511218 424102
rect 511274 424046 511342 424102
rect 511398 424046 511494 424102
rect 510874 423978 511494 424046
rect 510874 423922 510970 423978
rect 511026 423922 511094 423978
rect 511150 423922 511218 423978
rect 511274 423922 511342 423978
rect 511398 423922 511494 423978
rect 510874 406350 511494 423922
rect 510874 406294 510970 406350
rect 511026 406294 511094 406350
rect 511150 406294 511218 406350
rect 511274 406294 511342 406350
rect 511398 406294 511494 406350
rect 510874 406226 511494 406294
rect 510874 406170 510970 406226
rect 511026 406170 511094 406226
rect 511150 406170 511218 406226
rect 511274 406170 511342 406226
rect 511398 406170 511494 406226
rect 510874 406102 511494 406170
rect 510874 406046 510970 406102
rect 511026 406046 511094 406102
rect 511150 406046 511218 406102
rect 511274 406046 511342 406102
rect 511398 406046 511494 406102
rect 510874 405978 511494 406046
rect 510874 405922 510970 405978
rect 511026 405922 511094 405978
rect 511150 405922 511218 405978
rect 511274 405922 511342 405978
rect 511398 405922 511494 405978
rect 510874 388350 511494 405922
rect 510874 388294 510970 388350
rect 511026 388294 511094 388350
rect 511150 388294 511218 388350
rect 511274 388294 511342 388350
rect 511398 388294 511494 388350
rect 510874 388226 511494 388294
rect 510874 388170 510970 388226
rect 511026 388170 511094 388226
rect 511150 388170 511218 388226
rect 511274 388170 511342 388226
rect 511398 388170 511494 388226
rect 510874 388102 511494 388170
rect 510874 388046 510970 388102
rect 511026 388046 511094 388102
rect 511150 388046 511218 388102
rect 511274 388046 511342 388102
rect 511398 388046 511494 388102
rect 510874 387978 511494 388046
rect 510874 387922 510970 387978
rect 511026 387922 511094 387978
rect 511150 387922 511218 387978
rect 511274 387922 511342 387978
rect 511398 387922 511494 387978
rect 510874 370350 511494 387922
rect 510874 370294 510970 370350
rect 511026 370294 511094 370350
rect 511150 370294 511218 370350
rect 511274 370294 511342 370350
rect 511398 370294 511494 370350
rect 510874 370226 511494 370294
rect 510874 370170 510970 370226
rect 511026 370170 511094 370226
rect 511150 370170 511218 370226
rect 511274 370170 511342 370226
rect 511398 370170 511494 370226
rect 510874 370102 511494 370170
rect 510874 370046 510970 370102
rect 511026 370046 511094 370102
rect 511150 370046 511218 370102
rect 511274 370046 511342 370102
rect 511398 370046 511494 370102
rect 510874 369978 511494 370046
rect 510874 369922 510970 369978
rect 511026 369922 511094 369978
rect 511150 369922 511218 369978
rect 511274 369922 511342 369978
rect 511398 369922 511494 369978
rect 510874 352350 511494 369922
rect 510874 352294 510970 352350
rect 511026 352294 511094 352350
rect 511150 352294 511218 352350
rect 511274 352294 511342 352350
rect 511398 352294 511494 352350
rect 510874 352226 511494 352294
rect 510874 352170 510970 352226
rect 511026 352170 511094 352226
rect 511150 352170 511218 352226
rect 511274 352170 511342 352226
rect 511398 352170 511494 352226
rect 510874 352102 511494 352170
rect 510874 352046 510970 352102
rect 511026 352046 511094 352102
rect 511150 352046 511218 352102
rect 511274 352046 511342 352102
rect 511398 352046 511494 352102
rect 510874 351978 511494 352046
rect 510874 351922 510970 351978
rect 511026 351922 511094 351978
rect 511150 351922 511218 351978
rect 511274 351922 511342 351978
rect 511398 351922 511494 351978
rect 510874 334350 511494 351922
rect 510874 334294 510970 334350
rect 511026 334294 511094 334350
rect 511150 334294 511218 334350
rect 511274 334294 511342 334350
rect 511398 334294 511494 334350
rect 510874 334226 511494 334294
rect 510874 334170 510970 334226
rect 511026 334170 511094 334226
rect 511150 334170 511218 334226
rect 511274 334170 511342 334226
rect 511398 334170 511494 334226
rect 510874 334102 511494 334170
rect 510874 334046 510970 334102
rect 511026 334046 511094 334102
rect 511150 334046 511218 334102
rect 511274 334046 511342 334102
rect 511398 334046 511494 334102
rect 510874 333978 511494 334046
rect 510874 333922 510970 333978
rect 511026 333922 511094 333978
rect 511150 333922 511218 333978
rect 511274 333922 511342 333978
rect 511398 333922 511494 333978
rect 510874 316350 511494 333922
rect 510874 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 511494 316350
rect 510874 316226 511494 316294
rect 510874 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 511494 316226
rect 510874 316102 511494 316170
rect 510874 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 511494 316102
rect 510874 315978 511494 316046
rect 510874 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 511494 315978
rect 510874 298350 511494 315922
rect 510874 298294 510970 298350
rect 511026 298294 511094 298350
rect 511150 298294 511218 298350
rect 511274 298294 511342 298350
rect 511398 298294 511494 298350
rect 510874 298226 511494 298294
rect 510874 298170 510970 298226
rect 511026 298170 511094 298226
rect 511150 298170 511218 298226
rect 511274 298170 511342 298226
rect 511398 298170 511494 298226
rect 510874 298102 511494 298170
rect 510874 298046 510970 298102
rect 511026 298046 511094 298102
rect 511150 298046 511218 298102
rect 511274 298046 511342 298102
rect 511398 298046 511494 298102
rect 510874 297978 511494 298046
rect 510874 297922 510970 297978
rect 511026 297922 511094 297978
rect 511150 297922 511218 297978
rect 511274 297922 511342 297978
rect 511398 297922 511494 297978
rect 510874 280350 511494 297922
rect 510874 280294 510970 280350
rect 511026 280294 511094 280350
rect 511150 280294 511218 280350
rect 511274 280294 511342 280350
rect 511398 280294 511494 280350
rect 510874 280226 511494 280294
rect 510874 280170 510970 280226
rect 511026 280170 511094 280226
rect 511150 280170 511218 280226
rect 511274 280170 511342 280226
rect 511398 280170 511494 280226
rect 510874 280102 511494 280170
rect 510874 280046 510970 280102
rect 511026 280046 511094 280102
rect 511150 280046 511218 280102
rect 511274 280046 511342 280102
rect 511398 280046 511494 280102
rect 510874 279978 511494 280046
rect 510874 279922 510970 279978
rect 511026 279922 511094 279978
rect 511150 279922 511218 279978
rect 511274 279922 511342 279978
rect 511398 279922 511494 279978
rect 510874 262350 511494 279922
rect 510874 262294 510970 262350
rect 511026 262294 511094 262350
rect 511150 262294 511218 262350
rect 511274 262294 511342 262350
rect 511398 262294 511494 262350
rect 510874 262226 511494 262294
rect 510874 262170 510970 262226
rect 511026 262170 511094 262226
rect 511150 262170 511218 262226
rect 511274 262170 511342 262226
rect 511398 262170 511494 262226
rect 510874 262102 511494 262170
rect 510874 262046 510970 262102
rect 511026 262046 511094 262102
rect 511150 262046 511218 262102
rect 511274 262046 511342 262102
rect 511398 262046 511494 262102
rect 510874 261978 511494 262046
rect 510874 261922 510970 261978
rect 511026 261922 511094 261978
rect 511150 261922 511218 261978
rect 511274 261922 511342 261978
rect 511398 261922 511494 261978
rect 510874 244350 511494 261922
rect 510874 244294 510970 244350
rect 511026 244294 511094 244350
rect 511150 244294 511218 244350
rect 511274 244294 511342 244350
rect 511398 244294 511494 244350
rect 510874 244226 511494 244294
rect 510874 244170 510970 244226
rect 511026 244170 511094 244226
rect 511150 244170 511218 244226
rect 511274 244170 511342 244226
rect 511398 244170 511494 244226
rect 510874 244102 511494 244170
rect 510874 244046 510970 244102
rect 511026 244046 511094 244102
rect 511150 244046 511218 244102
rect 511274 244046 511342 244102
rect 511398 244046 511494 244102
rect 510874 243978 511494 244046
rect 510874 243922 510970 243978
rect 511026 243922 511094 243978
rect 511150 243922 511218 243978
rect 511274 243922 511342 243978
rect 511398 243922 511494 243978
rect 510874 226350 511494 243922
rect 510874 226294 510970 226350
rect 511026 226294 511094 226350
rect 511150 226294 511218 226350
rect 511274 226294 511342 226350
rect 511398 226294 511494 226350
rect 510874 226226 511494 226294
rect 510874 226170 510970 226226
rect 511026 226170 511094 226226
rect 511150 226170 511218 226226
rect 511274 226170 511342 226226
rect 511398 226170 511494 226226
rect 510874 226102 511494 226170
rect 510874 226046 510970 226102
rect 511026 226046 511094 226102
rect 511150 226046 511218 226102
rect 511274 226046 511342 226102
rect 511398 226046 511494 226102
rect 510874 225978 511494 226046
rect 510874 225922 510970 225978
rect 511026 225922 511094 225978
rect 511150 225922 511218 225978
rect 511274 225922 511342 225978
rect 511398 225922 511494 225978
rect 510874 208350 511494 225922
rect 510874 208294 510970 208350
rect 511026 208294 511094 208350
rect 511150 208294 511218 208350
rect 511274 208294 511342 208350
rect 511398 208294 511494 208350
rect 510874 208226 511494 208294
rect 510874 208170 510970 208226
rect 511026 208170 511094 208226
rect 511150 208170 511218 208226
rect 511274 208170 511342 208226
rect 511398 208170 511494 208226
rect 510874 208102 511494 208170
rect 510874 208046 510970 208102
rect 511026 208046 511094 208102
rect 511150 208046 511218 208102
rect 511274 208046 511342 208102
rect 511398 208046 511494 208102
rect 510874 207978 511494 208046
rect 510874 207922 510970 207978
rect 511026 207922 511094 207978
rect 511150 207922 511218 207978
rect 511274 207922 511342 207978
rect 511398 207922 511494 207978
rect 510874 190350 511494 207922
rect 510874 190294 510970 190350
rect 511026 190294 511094 190350
rect 511150 190294 511218 190350
rect 511274 190294 511342 190350
rect 511398 190294 511494 190350
rect 510874 190226 511494 190294
rect 510874 190170 510970 190226
rect 511026 190170 511094 190226
rect 511150 190170 511218 190226
rect 511274 190170 511342 190226
rect 511398 190170 511494 190226
rect 510874 190102 511494 190170
rect 510874 190046 510970 190102
rect 511026 190046 511094 190102
rect 511150 190046 511218 190102
rect 511274 190046 511342 190102
rect 511398 190046 511494 190102
rect 510874 189978 511494 190046
rect 510874 189922 510970 189978
rect 511026 189922 511094 189978
rect 511150 189922 511218 189978
rect 511274 189922 511342 189978
rect 511398 189922 511494 189978
rect 510874 172350 511494 189922
rect 510874 172294 510970 172350
rect 511026 172294 511094 172350
rect 511150 172294 511218 172350
rect 511274 172294 511342 172350
rect 511398 172294 511494 172350
rect 510874 172226 511494 172294
rect 510874 172170 510970 172226
rect 511026 172170 511094 172226
rect 511150 172170 511218 172226
rect 511274 172170 511342 172226
rect 511398 172170 511494 172226
rect 510874 172102 511494 172170
rect 510874 172046 510970 172102
rect 511026 172046 511094 172102
rect 511150 172046 511218 172102
rect 511274 172046 511342 172102
rect 511398 172046 511494 172102
rect 510874 171978 511494 172046
rect 510874 171922 510970 171978
rect 511026 171922 511094 171978
rect 511150 171922 511218 171978
rect 511274 171922 511342 171978
rect 511398 171922 511494 171978
rect 510874 154350 511494 171922
rect 510874 154294 510970 154350
rect 511026 154294 511094 154350
rect 511150 154294 511218 154350
rect 511274 154294 511342 154350
rect 511398 154294 511494 154350
rect 510874 154226 511494 154294
rect 510874 154170 510970 154226
rect 511026 154170 511094 154226
rect 511150 154170 511218 154226
rect 511274 154170 511342 154226
rect 511398 154170 511494 154226
rect 510874 154102 511494 154170
rect 510874 154046 510970 154102
rect 511026 154046 511094 154102
rect 511150 154046 511218 154102
rect 511274 154046 511342 154102
rect 511398 154046 511494 154102
rect 510874 153978 511494 154046
rect 510874 153922 510970 153978
rect 511026 153922 511094 153978
rect 511150 153922 511218 153978
rect 511274 153922 511342 153978
rect 511398 153922 511494 153978
rect 510874 136350 511494 153922
rect 510874 136294 510970 136350
rect 511026 136294 511094 136350
rect 511150 136294 511218 136350
rect 511274 136294 511342 136350
rect 511398 136294 511494 136350
rect 510874 136226 511494 136294
rect 510874 136170 510970 136226
rect 511026 136170 511094 136226
rect 511150 136170 511218 136226
rect 511274 136170 511342 136226
rect 511398 136170 511494 136226
rect 510874 136102 511494 136170
rect 510874 136046 510970 136102
rect 511026 136046 511094 136102
rect 511150 136046 511218 136102
rect 511274 136046 511342 136102
rect 511398 136046 511494 136102
rect 510874 135978 511494 136046
rect 510874 135922 510970 135978
rect 511026 135922 511094 135978
rect 511150 135922 511218 135978
rect 511274 135922 511342 135978
rect 511398 135922 511494 135978
rect 510874 118350 511494 135922
rect 510874 118294 510970 118350
rect 511026 118294 511094 118350
rect 511150 118294 511218 118350
rect 511274 118294 511342 118350
rect 511398 118294 511494 118350
rect 510874 118226 511494 118294
rect 510874 118170 510970 118226
rect 511026 118170 511094 118226
rect 511150 118170 511218 118226
rect 511274 118170 511342 118226
rect 511398 118170 511494 118226
rect 510874 118102 511494 118170
rect 510874 118046 510970 118102
rect 511026 118046 511094 118102
rect 511150 118046 511218 118102
rect 511274 118046 511342 118102
rect 511398 118046 511494 118102
rect 510874 117978 511494 118046
rect 510874 117922 510970 117978
rect 511026 117922 511094 117978
rect 511150 117922 511218 117978
rect 511274 117922 511342 117978
rect 511398 117922 511494 117978
rect 510874 100350 511494 117922
rect 510874 100294 510970 100350
rect 511026 100294 511094 100350
rect 511150 100294 511218 100350
rect 511274 100294 511342 100350
rect 511398 100294 511494 100350
rect 510874 100226 511494 100294
rect 510874 100170 510970 100226
rect 511026 100170 511094 100226
rect 511150 100170 511218 100226
rect 511274 100170 511342 100226
rect 511398 100170 511494 100226
rect 510874 100102 511494 100170
rect 510874 100046 510970 100102
rect 511026 100046 511094 100102
rect 511150 100046 511218 100102
rect 511274 100046 511342 100102
rect 511398 100046 511494 100102
rect 510874 99978 511494 100046
rect 510874 99922 510970 99978
rect 511026 99922 511094 99978
rect 511150 99922 511218 99978
rect 511274 99922 511342 99978
rect 511398 99922 511494 99978
rect 510874 82350 511494 99922
rect 510874 82294 510970 82350
rect 511026 82294 511094 82350
rect 511150 82294 511218 82350
rect 511274 82294 511342 82350
rect 511398 82294 511494 82350
rect 510874 82226 511494 82294
rect 510874 82170 510970 82226
rect 511026 82170 511094 82226
rect 511150 82170 511218 82226
rect 511274 82170 511342 82226
rect 511398 82170 511494 82226
rect 510874 82102 511494 82170
rect 510874 82046 510970 82102
rect 511026 82046 511094 82102
rect 511150 82046 511218 82102
rect 511274 82046 511342 82102
rect 511398 82046 511494 82102
rect 510874 81978 511494 82046
rect 510874 81922 510970 81978
rect 511026 81922 511094 81978
rect 511150 81922 511218 81978
rect 511274 81922 511342 81978
rect 511398 81922 511494 81978
rect 510874 64350 511494 81922
rect 510874 64294 510970 64350
rect 511026 64294 511094 64350
rect 511150 64294 511218 64350
rect 511274 64294 511342 64350
rect 511398 64294 511494 64350
rect 510874 64226 511494 64294
rect 510874 64170 510970 64226
rect 511026 64170 511094 64226
rect 511150 64170 511218 64226
rect 511274 64170 511342 64226
rect 511398 64170 511494 64226
rect 510874 64102 511494 64170
rect 510874 64046 510970 64102
rect 511026 64046 511094 64102
rect 511150 64046 511218 64102
rect 511274 64046 511342 64102
rect 511398 64046 511494 64102
rect 510874 63978 511494 64046
rect 510874 63922 510970 63978
rect 511026 63922 511094 63978
rect 511150 63922 511218 63978
rect 511274 63922 511342 63978
rect 511398 63922 511494 63978
rect 510874 46350 511494 63922
rect 510874 46294 510970 46350
rect 511026 46294 511094 46350
rect 511150 46294 511218 46350
rect 511274 46294 511342 46350
rect 511398 46294 511494 46350
rect 510874 46226 511494 46294
rect 510874 46170 510970 46226
rect 511026 46170 511094 46226
rect 511150 46170 511218 46226
rect 511274 46170 511342 46226
rect 511398 46170 511494 46226
rect 510874 46102 511494 46170
rect 510874 46046 510970 46102
rect 511026 46046 511094 46102
rect 511150 46046 511218 46102
rect 511274 46046 511342 46102
rect 511398 46046 511494 46102
rect 510874 45978 511494 46046
rect 510874 45922 510970 45978
rect 511026 45922 511094 45978
rect 511150 45922 511218 45978
rect 511274 45922 511342 45978
rect 511398 45922 511494 45978
rect 510874 28350 511494 45922
rect 510874 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 511494 28350
rect 510874 28226 511494 28294
rect 510874 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 511494 28226
rect 510874 28102 511494 28170
rect 510874 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 511494 28102
rect 510874 27978 511494 28046
rect 510874 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 511494 27978
rect 510874 10350 511494 27922
rect 510874 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 511494 10350
rect 510874 10226 511494 10294
rect 510874 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 511494 10226
rect 510874 10102 511494 10170
rect 510874 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 511494 10102
rect 510874 9978 511494 10046
rect 510874 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 511494 9978
rect 510874 -1120 511494 9922
rect 510874 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 511494 -1120
rect 510874 -1244 511494 -1176
rect 510874 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 511494 -1244
rect 510874 -1368 511494 -1300
rect 510874 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 511494 -1368
rect 510874 -1492 511494 -1424
rect 510874 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 511494 -1492
rect 510874 -1644 511494 -1548
rect 525154 597212 525774 598268
rect 525154 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 525774 597212
rect 525154 597088 525774 597156
rect 525154 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 525774 597088
rect 525154 596964 525774 597032
rect 525154 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 525774 596964
rect 525154 596840 525774 596908
rect 525154 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 525774 596840
rect 525154 580350 525774 596784
rect 525154 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 525774 580350
rect 525154 580226 525774 580294
rect 525154 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 525774 580226
rect 525154 580102 525774 580170
rect 525154 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 525774 580102
rect 525154 579978 525774 580046
rect 525154 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 525774 579978
rect 525154 562350 525774 579922
rect 525154 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 525774 562350
rect 525154 562226 525774 562294
rect 525154 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 525774 562226
rect 525154 562102 525774 562170
rect 525154 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 525774 562102
rect 525154 561978 525774 562046
rect 525154 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 525774 561978
rect 525154 544350 525774 561922
rect 525154 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 525774 544350
rect 525154 544226 525774 544294
rect 525154 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 525774 544226
rect 525154 544102 525774 544170
rect 525154 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 525774 544102
rect 525154 543978 525774 544046
rect 525154 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 525774 543978
rect 525154 526350 525774 543922
rect 525154 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 525774 526350
rect 525154 526226 525774 526294
rect 525154 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 525774 526226
rect 525154 526102 525774 526170
rect 525154 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 525774 526102
rect 525154 525978 525774 526046
rect 525154 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 525774 525978
rect 525154 508350 525774 525922
rect 525154 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 525774 508350
rect 525154 508226 525774 508294
rect 525154 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 525774 508226
rect 525154 508102 525774 508170
rect 525154 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 525774 508102
rect 525154 507978 525774 508046
rect 525154 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 525774 507978
rect 525154 490350 525774 507922
rect 525154 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 525774 490350
rect 525154 490226 525774 490294
rect 525154 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 525774 490226
rect 525154 490102 525774 490170
rect 525154 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 525774 490102
rect 525154 489978 525774 490046
rect 525154 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 525774 489978
rect 525154 472350 525774 489922
rect 525154 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 525774 472350
rect 525154 472226 525774 472294
rect 525154 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 525774 472226
rect 525154 472102 525774 472170
rect 525154 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 525774 472102
rect 525154 471978 525774 472046
rect 525154 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 525774 471978
rect 525154 454350 525774 471922
rect 525154 454294 525250 454350
rect 525306 454294 525374 454350
rect 525430 454294 525498 454350
rect 525554 454294 525622 454350
rect 525678 454294 525774 454350
rect 525154 454226 525774 454294
rect 525154 454170 525250 454226
rect 525306 454170 525374 454226
rect 525430 454170 525498 454226
rect 525554 454170 525622 454226
rect 525678 454170 525774 454226
rect 525154 454102 525774 454170
rect 525154 454046 525250 454102
rect 525306 454046 525374 454102
rect 525430 454046 525498 454102
rect 525554 454046 525622 454102
rect 525678 454046 525774 454102
rect 525154 453978 525774 454046
rect 525154 453922 525250 453978
rect 525306 453922 525374 453978
rect 525430 453922 525498 453978
rect 525554 453922 525622 453978
rect 525678 453922 525774 453978
rect 525154 436350 525774 453922
rect 525154 436294 525250 436350
rect 525306 436294 525374 436350
rect 525430 436294 525498 436350
rect 525554 436294 525622 436350
rect 525678 436294 525774 436350
rect 525154 436226 525774 436294
rect 525154 436170 525250 436226
rect 525306 436170 525374 436226
rect 525430 436170 525498 436226
rect 525554 436170 525622 436226
rect 525678 436170 525774 436226
rect 525154 436102 525774 436170
rect 525154 436046 525250 436102
rect 525306 436046 525374 436102
rect 525430 436046 525498 436102
rect 525554 436046 525622 436102
rect 525678 436046 525774 436102
rect 525154 435978 525774 436046
rect 525154 435922 525250 435978
rect 525306 435922 525374 435978
rect 525430 435922 525498 435978
rect 525554 435922 525622 435978
rect 525678 435922 525774 435978
rect 525154 418350 525774 435922
rect 525154 418294 525250 418350
rect 525306 418294 525374 418350
rect 525430 418294 525498 418350
rect 525554 418294 525622 418350
rect 525678 418294 525774 418350
rect 525154 418226 525774 418294
rect 525154 418170 525250 418226
rect 525306 418170 525374 418226
rect 525430 418170 525498 418226
rect 525554 418170 525622 418226
rect 525678 418170 525774 418226
rect 525154 418102 525774 418170
rect 525154 418046 525250 418102
rect 525306 418046 525374 418102
rect 525430 418046 525498 418102
rect 525554 418046 525622 418102
rect 525678 418046 525774 418102
rect 525154 417978 525774 418046
rect 525154 417922 525250 417978
rect 525306 417922 525374 417978
rect 525430 417922 525498 417978
rect 525554 417922 525622 417978
rect 525678 417922 525774 417978
rect 525154 400350 525774 417922
rect 525154 400294 525250 400350
rect 525306 400294 525374 400350
rect 525430 400294 525498 400350
rect 525554 400294 525622 400350
rect 525678 400294 525774 400350
rect 525154 400226 525774 400294
rect 525154 400170 525250 400226
rect 525306 400170 525374 400226
rect 525430 400170 525498 400226
rect 525554 400170 525622 400226
rect 525678 400170 525774 400226
rect 525154 400102 525774 400170
rect 525154 400046 525250 400102
rect 525306 400046 525374 400102
rect 525430 400046 525498 400102
rect 525554 400046 525622 400102
rect 525678 400046 525774 400102
rect 525154 399978 525774 400046
rect 525154 399922 525250 399978
rect 525306 399922 525374 399978
rect 525430 399922 525498 399978
rect 525554 399922 525622 399978
rect 525678 399922 525774 399978
rect 525154 382350 525774 399922
rect 525154 382294 525250 382350
rect 525306 382294 525374 382350
rect 525430 382294 525498 382350
rect 525554 382294 525622 382350
rect 525678 382294 525774 382350
rect 525154 382226 525774 382294
rect 525154 382170 525250 382226
rect 525306 382170 525374 382226
rect 525430 382170 525498 382226
rect 525554 382170 525622 382226
rect 525678 382170 525774 382226
rect 525154 382102 525774 382170
rect 525154 382046 525250 382102
rect 525306 382046 525374 382102
rect 525430 382046 525498 382102
rect 525554 382046 525622 382102
rect 525678 382046 525774 382102
rect 525154 381978 525774 382046
rect 525154 381922 525250 381978
rect 525306 381922 525374 381978
rect 525430 381922 525498 381978
rect 525554 381922 525622 381978
rect 525678 381922 525774 381978
rect 525154 364350 525774 381922
rect 525154 364294 525250 364350
rect 525306 364294 525374 364350
rect 525430 364294 525498 364350
rect 525554 364294 525622 364350
rect 525678 364294 525774 364350
rect 525154 364226 525774 364294
rect 525154 364170 525250 364226
rect 525306 364170 525374 364226
rect 525430 364170 525498 364226
rect 525554 364170 525622 364226
rect 525678 364170 525774 364226
rect 525154 364102 525774 364170
rect 525154 364046 525250 364102
rect 525306 364046 525374 364102
rect 525430 364046 525498 364102
rect 525554 364046 525622 364102
rect 525678 364046 525774 364102
rect 525154 363978 525774 364046
rect 525154 363922 525250 363978
rect 525306 363922 525374 363978
rect 525430 363922 525498 363978
rect 525554 363922 525622 363978
rect 525678 363922 525774 363978
rect 525154 346350 525774 363922
rect 525154 346294 525250 346350
rect 525306 346294 525374 346350
rect 525430 346294 525498 346350
rect 525554 346294 525622 346350
rect 525678 346294 525774 346350
rect 525154 346226 525774 346294
rect 525154 346170 525250 346226
rect 525306 346170 525374 346226
rect 525430 346170 525498 346226
rect 525554 346170 525622 346226
rect 525678 346170 525774 346226
rect 525154 346102 525774 346170
rect 525154 346046 525250 346102
rect 525306 346046 525374 346102
rect 525430 346046 525498 346102
rect 525554 346046 525622 346102
rect 525678 346046 525774 346102
rect 525154 345978 525774 346046
rect 525154 345922 525250 345978
rect 525306 345922 525374 345978
rect 525430 345922 525498 345978
rect 525554 345922 525622 345978
rect 525678 345922 525774 345978
rect 525154 328350 525774 345922
rect 525154 328294 525250 328350
rect 525306 328294 525374 328350
rect 525430 328294 525498 328350
rect 525554 328294 525622 328350
rect 525678 328294 525774 328350
rect 525154 328226 525774 328294
rect 525154 328170 525250 328226
rect 525306 328170 525374 328226
rect 525430 328170 525498 328226
rect 525554 328170 525622 328226
rect 525678 328170 525774 328226
rect 525154 328102 525774 328170
rect 525154 328046 525250 328102
rect 525306 328046 525374 328102
rect 525430 328046 525498 328102
rect 525554 328046 525622 328102
rect 525678 328046 525774 328102
rect 525154 327978 525774 328046
rect 525154 327922 525250 327978
rect 525306 327922 525374 327978
rect 525430 327922 525498 327978
rect 525554 327922 525622 327978
rect 525678 327922 525774 327978
rect 525154 310350 525774 327922
rect 525154 310294 525250 310350
rect 525306 310294 525374 310350
rect 525430 310294 525498 310350
rect 525554 310294 525622 310350
rect 525678 310294 525774 310350
rect 525154 310226 525774 310294
rect 525154 310170 525250 310226
rect 525306 310170 525374 310226
rect 525430 310170 525498 310226
rect 525554 310170 525622 310226
rect 525678 310170 525774 310226
rect 525154 310102 525774 310170
rect 525154 310046 525250 310102
rect 525306 310046 525374 310102
rect 525430 310046 525498 310102
rect 525554 310046 525622 310102
rect 525678 310046 525774 310102
rect 525154 309978 525774 310046
rect 525154 309922 525250 309978
rect 525306 309922 525374 309978
rect 525430 309922 525498 309978
rect 525554 309922 525622 309978
rect 525678 309922 525774 309978
rect 525154 292350 525774 309922
rect 525154 292294 525250 292350
rect 525306 292294 525374 292350
rect 525430 292294 525498 292350
rect 525554 292294 525622 292350
rect 525678 292294 525774 292350
rect 525154 292226 525774 292294
rect 525154 292170 525250 292226
rect 525306 292170 525374 292226
rect 525430 292170 525498 292226
rect 525554 292170 525622 292226
rect 525678 292170 525774 292226
rect 525154 292102 525774 292170
rect 525154 292046 525250 292102
rect 525306 292046 525374 292102
rect 525430 292046 525498 292102
rect 525554 292046 525622 292102
rect 525678 292046 525774 292102
rect 525154 291978 525774 292046
rect 525154 291922 525250 291978
rect 525306 291922 525374 291978
rect 525430 291922 525498 291978
rect 525554 291922 525622 291978
rect 525678 291922 525774 291978
rect 525154 274350 525774 291922
rect 525154 274294 525250 274350
rect 525306 274294 525374 274350
rect 525430 274294 525498 274350
rect 525554 274294 525622 274350
rect 525678 274294 525774 274350
rect 525154 274226 525774 274294
rect 525154 274170 525250 274226
rect 525306 274170 525374 274226
rect 525430 274170 525498 274226
rect 525554 274170 525622 274226
rect 525678 274170 525774 274226
rect 525154 274102 525774 274170
rect 525154 274046 525250 274102
rect 525306 274046 525374 274102
rect 525430 274046 525498 274102
rect 525554 274046 525622 274102
rect 525678 274046 525774 274102
rect 525154 273978 525774 274046
rect 525154 273922 525250 273978
rect 525306 273922 525374 273978
rect 525430 273922 525498 273978
rect 525554 273922 525622 273978
rect 525678 273922 525774 273978
rect 525154 256350 525774 273922
rect 525154 256294 525250 256350
rect 525306 256294 525374 256350
rect 525430 256294 525498 256350
rect 525554 256294 525622 256350
rect 525678 256294 525774 256350
rect 525154 256226 525774 256294
rect 525154 256170 525250 256226
rect 525306 256170 525374 256226
rect 525430 256170 525498 256226
rect 525554 256170 525622 256226
rect 525678 256170 525774 256226
rect 525154 256102 525774 256170
rect 525154 256046 525250 256102
rect 525306 256046 525374 256102
rect 525430 256046 525498 256102
rect 525554 256046 525622 256102
rect 525678 256046 525774 256102
rect 525154 255978 525774 256046
rect 525154 255922 525250 255978
rect 525306 255922 525374 255978
rect 525430 255922 525498 255978
rect 525554 255922 525622 255978
rect 525678 255922 525774 255978
rect 525154 238350 525774 255922
rect 525154 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 525774 238350
rect 525154 238226 525774 238294
rect 525154 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 525774 238226
rect 525154 238102 525774 238170
rect 525154 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 525774 238102
rect 525154 237978 525774 238046
rect 525154 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 525774 237978
rect 525154 220350 525774 237922
rect 525154 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 525774 220350
rect 525154 220226 525774 220294
rect 525154 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 525774 220226
rect 525154 220102 525774 220170
rect 525154 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 525774 220102
rect 525154 219978 525774 220046
rect 525154 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 525774 219978
rect 525154 202350 525774 219922
rect 525154 202294 525250 202350
rect 525306 202294 525374 202350
rect 525430 202294 525498 202350
rect 525554 202294 525622 202350
rect 525678 202294 525774 202350
rect 525154 202226 525774 202294
rect 525154 202170 525250 202226
rect 525306 202170 525374 202226
rect 525430 202170 525498 202226
rect 525554 202170 525622 202226
rect 525678 202170 525774 202226
rect 525154 202102 525774 202170
rect 525154 202046 525250 202102
rect 525306 202046 525374 202102
rect 525430 202046 525498 202102
rect 525554 202046 525622 202102
rect 525678 202046 525774 202102
rect 525154 201978 525774 202046
rect 525154 201922 525250 201978
rect 525306 201922 525374 201978
rect 525430 201922 525498 201978
rect 525554 201922 525622 201978
rect 525678 201922 525774 201978
rect 525154 184350 525774 201922
rect 525154 184294 525250 184350
rect 525306 184294 525374 184350
rect 525430 184294 525498 184350
rect 525554 184294 525622 184350
rect 525678 184294 525774 184350
rect 525154 184226 525774 184294
rect 525154 184170 525250 184226
rect 525306 184170 525374 184226
rect 525430 184170 525498 184226
rect 525554 184170 525622 184226
rect 525678 184170 525774 184226
rect 525154 184102 525774 184170
rect 525154 184046 525250 184102
rect 525306 184046 525374 184102
rect 525430 184046 525498 184102
rect 525554 184046 525622 184102
rect 525678 184046 525774 184102
rect 525154 183978 525774 184046
rect 525154 183922 525250 183978
rect 525306 183922 525374 183978
rect 525430 183922 525498 183978
rect 525554 183922 525622 183978
rect 525678 183922 525774 183978
rect 525154 166350 525774 183922
rect 525154 166294 525250 166350
rect 525306 166294 525374 166350
rect 525430 166294 525498 166350
rect 525554 166294 525622 166350
rect 525678 166294 525774 166350
rect 525154 166226 525774 166294
rect 525154 166170 525250 166226
rect 525306 166170 525374 166226
rect 525430 166170 525498 166226
rect 525554 166170 525622 166226
rect 525678 166170 525774 166226
rect 525154 166102 525774 166170
rect 525154 166046 525250 166102
rect 525306 166046 525374 166102
rect 525430 166046 525498 166102
rect 525554 166046 525622 166102
rect 525678 166046 525774 166102
rect 525154 165978 525774 166046
rect 525154 165922 525250 165978
rect 525306 165922 525374 165978
rect 525430 165922 525498 165978
rect 525554 165922 525622 165978
rect 525678 165922 525774 165978
rect 525154 148350 525774 165922
rect 525154 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 525774 148350
rect 525154 148226 525774 148294
rect 525154 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 525774 148226
rect 525154 148102 525774 148170
rect 525154 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 525774 148102
rect 525154 147978 525774 148046
rect 525154 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 525774 147978
rect 525154 130350 525774 147922
rect 525154 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 525774 130350
rect 525154 130226 525774 130294
rect 525154 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 525774 130226
rect 525154 130102 525774 130170
rect 525154 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 525774 130102
rect 525154 129978 525774 130046
rect 525154 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 525774 129978
rect 525154 112350 525774 129922
rect 525154 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 525774 112350
rect 525154 112226 525774 112294
rect 525154 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 525774 112226
rect 525154 112102 525774 112170
rect 525154 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 525774 112102
rect 525154 111978 525774 112046
rect 525154 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 525774 111978
rect 525154 94350 525774 111922
rect 525154 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 525774 94350
rect 525154 94226 525774 94294
rect 525154 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 525774 94226
rect 525154 94102 525774 94170
rect 525154 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 525774 94102
rect 525154 93978 525774 94046
rect 525154 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 525774 93978
rect 525154 76350 525774 93922
rect 525154 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 525774 76350
rect 525154 76226 525774 76294
rect 525154 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 525774 76226
rect 525154 76102 525774 76170
rect 525154 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 525774 76102
rect 525154 75978 525774 76046
rect 525154 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 525774 75978
rect 525154 58350 525774 75922
rect 525154 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 525774 58350
rect 525154 58226 525774 58294
rect 525154 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 525774 58226
rect 525154 58102 525774 58170
rect 525154 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 525774 58102
rect 525154 57978 525774 58046
rect 525154 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 525774 57978
rect 525154 40350 525774 57922
rect 525154 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 525774 40350
rect 525154 40226 525774 40294
rect 525154 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 525774 40226
rect 525154 40102 525774 40170
rect 525154 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 525774 40102
rect 525154 39978 525774 40046
rect 525154 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 525774 39978
rect 525154 22350 525774 39922
rect 525154 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 525774 22350
rect 525154 22226 525774 22294
rect 525154 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 525774 22226
rect 525154 22102 525774 22170
rect 525154 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 525774 22102
rect 525154 21978 525774 22046
rect 525154 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 525774 21978
rect 525154 4350 525774 21922
rect 525154 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 525774 4350
rect 525154 4226 525774 4294
rect 525154 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 525774 4226
rect 525154 4102 525774 4170
rect 525154 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 525774 4102
rect 525154 3978 525774 4046
rect 525154 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 525774 3978
rect 525154 -160 525774 3922
rect 525154 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 525774 -160
rect 525154 -284 525774 -216
rect 525154 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 525774 -284
rect 525154 -408 525774 -340
rect 525154 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 525774 -408
rect 525154 -532 525774 -464
rect 525154 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 525774 -532
rect 525154 -1644 525774 -588
rect 528874 598172 529494 598268
rect 528874 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 529494 598172
rect 528874 598048 529494 598116
rect 528874 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 529494 598048
rect 528874 597924 529494 597992
rect 528874 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 529494 597924
rect 528874 597800 529494 597868
rect 528874 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 529494 597800
rect 528874 586350 529494 597744
rect 528874 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 529494 586350
rect 528874 586226 529494 586294
rect 528874 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 529494 586226
rect 528874 586102 529494 586170
rect 528874 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 529494 586102
rect 528874 585978 529494 586046
rect 528874 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 529494 585978
rect 528874 568350 529494 585922
rect 528874 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 529494 568350
rect 528874 568226 529494 568294
rect 528874 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 529494 568226
rect 528874 568102 529494 568170
rect 528874 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 529494 568102
rect 528874 567978 529494 568046
rect 528874 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 529494 567978
rect 528874 550350 529494 567922
rect 528874 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 529494 550350
rect 528874 550226 529494 550294
rect 528874 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 529494 550226
rect 528874 550102 529494 550170
rect 528874 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 529494 550102
rect 528874 549978 529494 550046
rect 528874 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 529494 549978
rect 528874 532350 529494 549922
rect 528874 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 529494 532350
rect 528874 532226 529494 532294
rect 528874 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 529494 532226
rect 528874 532102 529494 532170
rect 528874 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 529494 532102
rect 528874 531978 529494 532046
rect 528874 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 529494 531978
rect 528874 514350 529494 531922
rect 528874 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 529494 514350
rect 528874 514226 529494 514294
rect 528874 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 529494 514226
rect 528874 514102 529494 514170
rect 528874 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 529494 514102
rect 528874 513978 529494 514046
rect 528874 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 529494 513978
rect 528874 496350 529494 513922
rect 528874 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 529494 496350
rect 528874 496226 529494 496294
rect 528874 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 529494 496226
rect 528874 496102 529494 496170
rect 528874 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 529494 496102
rect 528874 495978 529494 496046
rect 528874 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 529494 495978
rect 528874 478350 529494 495922
rect 528874 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 529494 478350
rect 528874 478226 529494 478294
rect 528874 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 529494 478226
rect 528874 478102 529494 478170
rect 528874 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 529494 478102
rect 528874 477978 529494 478046
rect 528874 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 529494 477978
rect 528874 460350 529494 477922
rect 528874 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 529494 460350
rect 528874 460226 529494 460294
rect 528874 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 529494 460226
rect 528874 460102 529494 460170
rect 528874 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 529494 460102
rect 528874 459978 529494 460046
rect 528874 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 529494 459978
rect 528874 442350 529494 459922
rect 528874 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 529494 442350
rect 528874 442226 529494 442294
rect 528874 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 529494 442226
rect 528874 442102 529494 442170
rect 528874 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 529494 442102
rect 528874 441978 529494 442046
rect 528874 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 529494 441978
rect 528874 424350 529494 441922
rect 528874 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 529494 424350
rect 528874 424226 529494 424294
rect 528874 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 529494 424226
rect 528874 424102 529494 424170
rect 528874 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 529494 424102
rect 528874 423978 529494 424046
rect 528874 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 529494 423978
rect 528874 406350 529494 423922
rect 528874 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 529494 406350
rect 528874 406226 529494 406294
rect 528874 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 529494 406226
rect 528874 406102 529494 406170
rect 528874 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 529494 406102
rect 528874 405978 529494 406046
rect 528874 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 529494 405978
rect 528874 388350 529494 405922
rect 528874 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 529494 388350
rect 528874 388226 529494 388294
rect 528874 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 529494 388226
rect 528874 388102 529494 388170
rect 528874 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 529494 388102
rect 528874 387978 529494 388046
rect 528874 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 529494 387978
rect 528874 370350 529494 387922
rect 528874 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 529494 370350
rect 528874 370226 529494 370294
rect 528874 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 529494 370226
rect 528874 370102 529494 370170
rect 528874 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 529494 370102
rect 528874 369978 529494 370046
rect 528874 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 529494 369978
rect 528874 352350 529494 369922
rect 528874 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 529494 352350
rect 528874 352226 529494 352294
rect 528874 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 529494 352226
rect 528874 352102 529494 352170
rect 528874 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 529494 352102
rect 528874 351978 529494 352046
rect 528874 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 529494 351978
rect 528874 334350 529494 351922
rect 528874 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 529494 334350
rect 528874 334226 529494 334294
rect 528874 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 529494 334226
rect 528874 334102 529494 334170
rect 528874 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 529494 334102
rect 528874 333978 529494 334046
rect 528874 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 529494 333978
rect 528874 316350 529494 333922
rect 528874 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 529494 316350
rect 528874 316226 529494 316294
rect 528874 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 529494 316226
rect 528874 316102 529494 316170
rect 528874 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 529494 316102
rect 528874 315978 529494 316046
rect 528874 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 529494 315978
rect 528874 298350 529494 315922
rect 528874 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 529494 298350
rect 528874 298226 529494 298294
rect 528874 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 529494 298226
rect 528874 298102 529494 298170
rect 528874 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 529494 298102
rect 528874 297978 529494 298046
rect 528874 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 529494 297978
rect 528874 280350 529494 297922
rect 528874 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 529494 280350
rect 528874 280226 529494 280294
rect 528874 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 529494 280226
rect 528874 280102 529494 280170
rect 528874 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 529494 280102
rect 528874 279978 529494 280046
rect 528874 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 529494 279978
rect 528874 262350 529494 279922
rect 528874 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 529494 262350
rect 528874 262226 529494 262294
rect 528874 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 529494 262226
rect 528874 262102 529494 262170
rect 528874 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 529494 262102
rect 528874 261978 529494 262046
rect 528874 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 529494 261978
rect 528874 244350 529494 261922
rect 528874 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 529494 244350
rect 528874 244226 529494 244294
rect 528874 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 529494 244226
rect 528874 244102 529494 244170
rect 528874 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 529494 244102
rect 528874 243978 529494 244046
rect 528874 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 529494 243978
rect 528874 226350 529494 243922
rect 528874 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 529494 226350
rect 528874 226226 529494 226294
rect 528874 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 529494 226226
rect 528874 226102 529494 226170
rect 528874 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 529494 226102
rect 528874 225978 529494 226046
rect 528874 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 529494 225978
rect 528874 208350 529494 225922
rect 528874 208294 528970 208350
rect 529026 208294 529094 208350
rect 529150 208294 529218 208350
rect 529274 208294 529342 208350
rect 529398 208294 529494 208350
rect 528874 208226 529494 208294
rect 528874 208170 528970 208226
rect 529026 208170 529094 208226
rect 529150 208170 529218 208226
rect 529274 208170 529342 208226
rect 529398 208170 529494 208226
rect 528874 208102 529494 208170
rect 528874 208046 528970 208102
rect 529026 208046 529094 208102
rect 529150 208046 529218 208102
rect 529274 208046 529342 208102
rect 529398 208046 529494 208102
rect 528874 207978 529494 208046
rect 528874 207922 528970 207978
rect 529026 207922 529094 207978
rect 529150 207922 529218 207978
rect 529274 207922 529342 207978
rect 529398 207922 529494 207978
rect 528874 190350 529494 207922
rect 528874 190294 528970 190350
rect 529026 190294 529094 190350
rect 529150 190294 529218 190350
rect 529274 190294 529342 190350
rect 529398 190294 529494 190350
rect 528874 190226 529494 190294
rect 528874 190170 528970 190226
rect 529026 190170 529094 190226
rect 529150 190170 529218 190226
rect 529274 190170 529342 190226
rect 529398 190170 529494 190226
rect 528874 190102 529494 190170
rect 528874 190046 528970 190102
rect 529026 190046 529094 190102
rect 529150 190046 529218 190102
rect 529274 190046 529342 190102
rect 529398 190046 529494 190102
rect 528874 189978 529494 190046
rect 528874 189922 528970 189978
rect 529026 189922 529094 189978
rect 529150 189922 529218 189978
rect 529274 189922 529342 189978
rect 529398 189922 529494 189978
rect 528874 172350 529494 189922
rect 528874 172294 528970 172350
rect 529026 172294 529094 172350
rect 529150 172294 529218 172350
rect 529274 172294 529342 172350
rect 529398 172294 529494 172350
rect 528874 172226 529494 172294
rect 528874 172170 528970 172226
rect 529026 172170 529094 172226
rect 529150 172170 529218 172226
rect 529274 172170 529342 172226
rect 529398 172170 529494 172226
rect 528874 172102 529494 172170
rect 528874 172046 528970 172102
rect 529026 172046 529094 172102
rect 529150 172046 529218 172102
rect 529274 172046 529342 172102
rect 529398 172046 529494 172102
rect 528874 171978 529494 172046
rect 528874 171922 528970 171978
rect 529026 171922 529094 171978
rect 529150 171922 529218 171978
rect 529274 171922 529342 171978
rect 529398 171922 529494 171978
rect 528874 154350 529494 171922
rect 528874 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 529494 154350
rect 528874 154226 529494 154294
rect 528874 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 529494 154226
rect 528874 154102 529494 154170
rect 528874 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 529494 154102
rect 528874 153978 529494 154046
rect 528874 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 529494 153978
rect 528874 136350 529494 153922
rect 528874 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 529494 136350
rect 528874 136226 529494 136294
rect 528874 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 529494 136226
rect 528874 136102 529494 136170
rect 528874 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 529494 136102
rect 528874 135978 529494 136046
rect 528874 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 529494 135978
rect 528874 118350 529494 135922
rect 528874 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 529494 118350
rect 528874 118226 529494 118294
rect 528874 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 529494 118226
rect 528874 118102 529494 118170
rect 528874 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 529494 118102
rect 528874 117978 529494 118046
rect 528874 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 529494 117978
rect 528874 100350 529494 117922
rect 528874 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 529494 100350
rect 528874 100226 529494 100294
rect 528874 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 529494 100226
rect 528874 100102 529494 100170
rect 528874 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 529494 100102
rect 528874 99978 529494 100046
rect 528874 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 529494 99978
rect 528874 82350 529494 99922
rect 528874 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 529494 82350
rect 528874 82226 529494 82294
rect 528874 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 529494 82226
rect 528874 82102 529494 82170
rect 528874 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 529494 82102
rect 528874 81978 529494 82046
rect 528874 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 529494 81978
rect 528874 64350 529494 81922
rect 528874 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 529494 64350
rect 528874 64226 529494 64294
rect 528874 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 529494 64226
rect 528874 64102 529494 64170
rect 528874 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 529494 64102
rect 528874 63978 529494 64046
rect 528874 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 529494 63978
rect 528874 46350 529494 63922
rect 528874 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 529494 46350
rect 528874 46226 529494 46294
rect 528874 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 529494 46226
rect 528874 46102 529494 46170
rect 528874 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 529494 46102
rect 528874 45978 529494 46046
rect 528874 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 529494 45978
rect 528874 28350 529494 45922
rect 528874 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 529494 28350
rect 528874 28226 529494 28294
rect 528874 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 529494 28226
rect 528874 28102 529494 28170
rect 528874 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 529494 28102
rect 528874 27978 529494 28046
rect 528874 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 529494 27978
rect 528874 10350 529494 27922
rect 528874 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 529494 10350
rect 528874 10226 529494 10294
rect 528874 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 529494 10226
rect 528874 10102 529494 10170
rect 528874 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 529494 10102
rect 528874 9978 529494 10046
rect 528874 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 529494 9978
rect 528874 -1120 529494 9922
rect 528874 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 529494 -1120
rect 528874 -1244 529494 -1176
rect 528874 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 529494 -1244
rect 528874 -1368 529494 -1300
rect 528874 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 529494 -1368
rect 528874 -1492 529494 -1424
rect 528874 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 529494 -1492
rect 528874 -1644 529494 -1548
rect 543154 597212 543774 598268
rect 543154 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 543774 597212
rect 543154 597088 543774 597156
rect 543154 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 543774 597088
rect 543154 596964 543774 597032
rect 543154 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 543774 596964
rect 543154 596840 543774 596908
rect 543154 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 543774 596840
rect 543154 580350 543774 596784
rect 543154 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 543774 580350
rect 543154 580226 543774 580294
rect 543154 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 543774 580226
rect 543154 580102 543774 580170
rect 543154 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 543774 580102
rect 543154 579978 543774 580046
rect 543154 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 543774 579978
rect 543154 562350 543774 579922
rect 543154 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 543774 562350
rect 543154 562226 543774 562294
rect 543154 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 543774 562226
rect 543154 562102 543774 562170
rect 543154 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 543774 562102
rect 543154 561978 543774 562046
rect 543154 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 543774 561978
rect 543154 544350 543774 561922
rect 543154 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 543774 544350
rect 543154 544226 543774 544294
rect 543154 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 543774 544226
rect 543154 544102 543774 544170
rect 543154 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 543774 544102
rect 543154 543978 543774 544046
rect 543154 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 543774 543978
rect 543154 526350 543774 543922
rect 543154 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 543774 526350
rect 543154 526226 543774 526294
rect 543154 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 543774 526226
rect 543154 526102 543774 526170
rect 543154 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 543774 526102
rect 543154 525978 543774 526046
rect 543154 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 543774 525978
rect 543154 508350 543774 525922
rect 543154 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 543774 508350
rect 543154 508226 543774 508294
rect 543154 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 543774 508226
rect 543154 508102 543774 508170
rect 543154 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 543774 508102
rect 543154 507978 543774 508046
rect 543154 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 543774 507978
rect 543154 490350 543774 507922
rect 543154 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 543774 490350
rect 543154 490226 543774 490294
rect 543154 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 543774 490226
rect 543154 490102 543774 490170
rect 543154 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 543774 490102
rect 543154 489978 543774 490046
rect 543154 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 543774 489978
rect 543154 472350 543774 489922
rect 543154 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 543774 472350
rect 543154 472226 543774 472294
rect 543154 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 543774 472226
rect 543154 472102 543774 472170
rect 543154 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 543774 472102
rect 543154 471978 543774 472046
rect 543154 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 543774 471978
rect 543154 454350 543774 471922
rect 543154 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 543774 454350
rect 543154 454226 543774 454294
rect 543154 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 543774 454226
rect 543154 454102 543774 454170
rect 543154 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 543774 454102
rect 543154 453978 543774 454046
rect 543154 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 543774 453978
rect 543154 436350 543774 453922
rect 543154 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 543774 436350
rect 543154 436226 543774 436294
rect 543154 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 543774 436226
rect 543154 436102 543774 436170
rect 543154 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 543774 436102
rect 543154 435978 543774 436046
rect 543154 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 543774 435978
rect 543154 418350 543774 435922
rect 543154 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 543774 418350
rect 543154 418226 543774 418294
rect 543154 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 543774 418226
rect 543154 418102 543774 418170
rect 543154 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 543774 418102
rect 543154 417978 543774 418046
rect 543154 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 543774 417978
rect 543154 400350 543774 417922
rect 543154 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 543774 400350
rect 543154 400226 543774 400294
rect 543154 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 543774 400226
rect 543154 400102 543774 400170
rect 543154 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 543774 400102
rect 543154 399978 543774 400046
rect 543154 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 543774 399978
rect 543154 382350 543774 399922
rect 543154 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 543774 382350
rect 543154 382226 543774 382294
rect 543154 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 543774 382226
rect 543154 382102 543774 382170
rect 543154 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 543774 382102
rect 543154 381978 543774 382046
rect 543154 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 543774 381978
rect 543154 364350 543774 381922
rect 543154 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 543774 364350
rect 543154 364226 543774 364294
rect 543154 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 543774 364226
rect 543154 364102 543774 364170
rect 543154 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 543774 364102
rect 543154 363978 543774 364046
rect 543154 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 543774 363978
rect 543154 346350 543774 363922
rect 543154 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 543774 346350
rect 543154 346226 543774 346294
rect 543154 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 543774 346226
rect 543154 346102 543774 346170
rect 543154 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 543774 346102
rect 543154 345978 543774 346046
rect 543154 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 543774 345978
rect 543154 328350 543774 345922
rect 543154 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 543774 328350
rect 543154 328226 543774 328294
rect 543154 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 543774 328226
rect 543154 328102 543774 328170
rect 543154 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 543774 328102
rect 543154 327978 543774 328046
rect 543154 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 543774 327978
rect 543154 310350 543774 327922
rect 543154 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 543774 310350
rect 543154 310226 543774 310294
rect 543154 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 543774 310226
rect 543154 310102 543774 310170
rect 543154 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 543774 310102
rect 543154 309978 543774 310046
rect 543154 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 543774 309978
rect 543154 292350 543774 309922
rect 543154 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 543774 292350
rect 543154 292226 543774 292294
rect 543154 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 543774 292226
rect 543154 292102 543774 292170
rect 543154 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 543774 292102
rect 543154 291978 543774 292046
rect 543154 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 543774 291978
rect 543154 274350 543774 291922
rect 543154 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 543774 274350
rect 543154 274226 543774 274294
rect 543154 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 543774 274226
rect 543154 274102 543774 274170
rect 543154 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 543774 274102
rect 543154 273978 543774 274046
rect 543154 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 543774 273978
rect 543154 256350 543774 273922
rect 543154 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 543774 256350
rect 543154 256226 543774 256294
rect 543154 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 543774 256226
rect 543154 256102 543774 256170
rect 543154 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 543774 256102
rect 543154 255978 543774 256046
rect 543154 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 543774 255978
rect 543154 238350 543774 255922
rect 543154 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 543774 238350
rect 543154 238226 543774 238294
rect 543154 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 543774 238226
rect 543154 238102 543774 238170
rect 543154 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 543774 238102
rect 543154 237978 543774 238046
rect 543154 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 543774 237978
rect 543154 220350 543774 237922
rect 543154 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 543774 220350
rect 543154 220226 543774 220294
rect 543154 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 543774 220226
rect 543154 220102 543774 220170
rect 543154 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 543774 220102
rect 543154 219978 543774 220046
rect 543154 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 543774 219978
rect 543154 202350 543774 219922
rect 543154 202294 543250 202350
rect 543306 202294 543374 202350
rect 543430 202294 543498 202350
rect 543554 202294 543622 202350
rect 543678 202294 543774 202350
rect 543154 202226 543774 202294
rect 543154 202170 543250 202226
rect 543306 202170 543374 202226
rect 543430 202170 543498 202226
rect 543554 202170 543622 202226
rect 543678 202170 543774 202226
rect 543154 202102 543774 202170
rect 543154 202046 543250 202102
rect 543306 202046 543374 202102
rect 543430 202046 543498 202102
rect 543554 202046 543622 202102
rect 543678 202046 543774 202102
rect 543154 201978 543774 202046
rect 543154 201922 543250 201978
rect 543306 201922 543374 201978
rect 543430 201922 543498 201978
rect 543554 201922 543622 201978
rect 543678 201922 543774 201978
rect 543154 184350 543774 201922
rect 543154 184294 543250 184350
rect 543306 184294 543374 184350
rect 543430 184294 543498 184350
rect 543554 184294 543622 184350
rect 543678 184294 543774 184350
rect 543154 184226 543774 184294
rect 543154 184170 543250 184226
rect 543306 184170 543374 184226
rect 543430 184170 543498 184226
rect 543554 184170 543622 184226
rect 543678 184170 543774 184226
rect 543154 184102 543774 184170
rect 543154 184046 543250 184102
rect 543306 184046 543374 184102
rect 543430 184046 543498 184102
rect 543554 184046 543622 184102
rect 543678 184046 543774 184102
rect 543154 183978 543774 184046
rect 543154 183922 543250 183978
rect 543306 183922 543374 183978
rect 543430 183922 543498 183978
rect 543554 183922 543622 183978
rect 543678 183922 543774 183978
rect 543154 166350 543774 183922
rect 543154 166294 543250 166350
rect 543306 166294 543374 166350
rect 543430 166294 543498 166350
rect 543554 166294 543622 166350
rect 543678 166294 543774 166350
rect 543154 166226 543774 166294
rect 543154 166170 543250 166226
rect 543306 166170 543374 166226
rect 543430 166170 543498 166226
rect 543554 166170 543622 166226
rect 543678 166170 543774 166226
rect 543154 166102 543774 166170
rect 543154 166046 543250 166102
rect 543306 166046 543374 166102
rect 543430 166046 543498 166102
rect 543554 166046 543622 166102
rect 543678 166046 543774 166102
rect 543154 165978 543774 166046
rect 543154 165922 543250 165978
rect 543306 165922 543374 165978
rect 543430 165922 543498 165978
rect 543554 165922 543622 165978
rect 543678 165922 543774 165978
rect 543154 148350 543774 165922
rect 543154 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 543774 148350
rect 543154 148226 543774 148294
rect 543154 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 543774 148226
rect 543154 148102 543774 148170
rect 543154 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 543774 148102
rect 543154 147978 543774 148046
rect 543154 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 543774 147978
rect 543154 130350 543774 147922
rect 543154 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 543774 130350
rect 543154 130226 543774 130294
rect 543154 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 543774 130226
rect 543154 130102 543774 130170
rect 543154 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 543774 130102
rect 543154 129978 543774 130046
rect 543154 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 543774 129978
rect 543154 112350 543774 129922
rect 543154 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 543774 112350
rect 543154 112226 543774 112294
rect 543154 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 543774 112226
rect 543154 112102 543774 112170
rect 543154 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 543774 112102
rect 543154 111978 543774 112046
rect 543154 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 543774 111978
rect 543154 94350 543774 111922
rect 543154 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 543774 94350
rect 543154 94226 543774 94294
rect 543154 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 543774 94226
rect 543154 94102 543774 94170
rect 543154 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 543774 94102
rect 543154 93978 543774 94046
rect 543154 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 543774 93978
rect 543154 76350 543774 93922
rect 543154 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 543774 76350
rect 543154 76226 543774 76294
rect 543154 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 543774 76226
rect 543154 76102 543774 76170
rect 543154 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 543774 76102
rect 543154 75978 543774 76046
rect 543154 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 543774 75978
rect 543154 58350 543774 75922
rect 543154 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 543774 58350
rect 543154 58226 543774 58294
rect 543154 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 543774 58226
rect 543154 58102 543774 58170
rect 543154 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 543774 58102
rect 543154 57978 543774 58046
rect 543154 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 543774 57978
rect 543154 40350 543774 57922
rect 543154 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 543774 40350
rect 543154 40226 543774 40294
rect 543154 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 543774 40226
rect 543154 40102 543774 40170
rect 543154 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 543774 40102
rect 543154 39978 543774 40046
rect 543154 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 543774 39978
rect 543154 22350 543774 39922
rect 543154 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 543774 22350
rect 543154 22226 543774 22294
rect 543154 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 543774 22226
rect 543154 22102 543774 22170
rect 543154 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 543774 22102
rect 543154 21978 543774 22046
rect 543154 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 543774 21978
rect 543154 4350 543774 21922
rect 543154 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 543774 4350
rect 543154 4226 543774 4294
rect 543154 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 543774 4226
rect 543154 4102 543774 4170
rect 543154 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 543774 4102
rect 543154 3978 543774 4046
rect 543154 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 543774 3978
rect 543154 -160 543774 3922
rect 543154 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 543774 -160
rect 543154 -284 543774 -216
rect 543154 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 543774 -284
rect 543154 -408 543774 -340
rect 543154 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 543774 -408
rect 543154 -532 543774 -464
rect 543154 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 543774 -532
rect 543154 -1644 543774 -588
rect 546874 598172 547494 598268
rect 546874 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 547494 598172
rect 546874 598048 547494 598116
rect 546874 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 547494 598048
rect 546874 597924 547494 597992
rect 546874 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 547494 597924
rect 546874 597800 547494 597868
rect 546874 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 547494 597800
rect 546874 586350 547494 597744
rect 546874 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 547494 586350
rect 546874 586226 547494 586294
rect 546874 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 547494 586226
rect 546874 586102 547494 586170
rect 546874 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 547494 586102
rect 546874 585978 547494 586046
rect 546874 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 547494 585978
rect 546874 568350 547494 585922
rect 546874 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 547494 568350
rect 546874 568226 547494 568294
rect 546874 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 547494 568226
rect 546874 568102 547494 568170
rect 546874 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 547494 568102
rect 546874 567978 547494 568046
rect 546874 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 547494 567978
rect 546874 550350 547494 567922
rect 546874 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 547494 550350
rect 546874 550226 547494 550294
rect 546874 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 547494 550226
rect 546874 550102 547494 550170
rect 546874 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 547494 550102
rect 546874 549978 547494 550046
rect 546874 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 547494 549978
rect 546874 532350 547494 549922
rect 546874 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 547494 532350
rect 546874 532226 547494 532294
rect 546874 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 547494 532226
rect 546874 532102 547494 532170
rect 546874 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 547494 532102
rect 546874 531978 547494 532046
rect 546874 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 547494 531978
rect 546874 514350 547494 531922
rect 546874 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 547494 514350
rect 546874 514226 547494 514294
rect 546874 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 547494 514226
rect 546874 514102 547494 514170
rect 546874 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 547494 514102
rect 546874 513978 547494 514046
rect 546874 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 547494 513978
rect 546874 496350 547494 513922
rect 546874 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 547494 496350
rect 546874 496226 547494 496294
rect 546874 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 547494 496226
rect 546874 496102 547494 496170
rect 546874 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 547494 496102
rect 546874 495978 547494 496046
rect 546874 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 547494 495978
rect 546874 478350 547494 495922
rect 546874 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 547494 478350
rect 546874 478226 547494 478294
rect 546874 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 547494 478226
rect 546874 478102 547494 478170
rect 546874 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 547494 478102
rect 546874 477978 547494 478046
rect 546874 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 547494 477978
rect 546874 460350 547494 477922
rect 546874 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 547494 460350
rect 546874 460226 547494 460294
rect 546874 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 547494 460226
rect 546874 460102 547494 460170
rect 546874 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 547494 460102
rect 546874 459978 547494 460046
rect 546874 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 547494 459978
rect 546874 442350 547494 459922
rect 546874 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 547494 442350
rect 546874 442226 547494 442294
rect 546874 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 547494 442226
rect 546874 442102 547494 442170
rect 546874 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 547494 442102
rect 546874 441978 547494 442046
rect 546874 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 547494 441978
rect 546874 424350 547494 441922
rect 546874 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 547494 424350
rect 546874 424226 547494 424294
rect 546874 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 547494 424226
rect 546874 424102 547494 424170
rect 546874 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 547494 424102
rect 546874 423978 547494 424046
rect 546874 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 547494 423978
rect 546874 406350 547494 423922
rect 546874 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 547494 406350
rect 546874 406226 547494 406294
rect 546874 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 547494 406226
rect 546874 406102 547494 406170
rect 546874 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 547494 406102
rect 546874 405978 547494 406046
rect 546874 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 547494 405978
rect 546874 388350 547494 405922
rect 546874 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 547494 388350
rect 546874 388226 547494 388294
rect 546874 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 547494 388226
rect 546874 388102 547494 388170
rect 546874 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 547494 388102
rect 546874 387978 547494 388046
rect 546874 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 547494 387978
rect 546874 370350 547494 387922
rect 546874 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 547494 370350
rect 546874 370226 547494 370294
rect 546874 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 547494 370226
rect 546874 370102 547494 370170
rect 546874 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 547494 370102
rect 546874 369978 547494 370046
rect 546874 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 547494 369978
rect 546874 352350 547494 369922
rect 546874 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 547494 352350
rect 546874 352226 547494 352294
rect 546874 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 547494 352226
rect 546874 352102 547494 352170
rect 546874 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 547494 352102
rect 546874 351978 547494 352046
rect 546874 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 547494 351978
rect 546874 334350 547494 351922
rect 546874 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 547494 334350
rect 546874 334226 547494 334294
rect 546874 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 547494 334226
rect 546874 334102 547494 334170
rect 546874 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 547494 334102
rect 546874 333978 547494 334046
rect 546874 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 547494 333978
rect 546874 316350 547494 333922
rect 546874 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 547494 316350
rect 546874 316226 547494 316294
rect 546874 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 547494 316226
rect 546874 316102 547494 316170
rect 546874 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 547494 316102
rect 546874 315978 547494 316046
rect 546874 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 547494 315978
rect 546874 298350 547494 315922
rect 546874 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 547494 298350
rect 546874 298226 547494 298294
rect 546874 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 547494 298226
rect 546874 298102 547494 298170
rect 546874 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 547494 298102
rect 546874 297978 547494 298046
rect 546874 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 547494 297978
rect 546874 280350 547494 297922
rect 546874 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 547494 280350
rect 546874 280226 547494 280294
rect 546874 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 547494 280226
rect 546874 280102 547494 280170
rect 546874 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 547494 280102
rect 546874 279978 547494 280046
rect 546874 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 547494 279978
rect 546874 262350 547494 279922
rect 546874 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 547494 262350
rect 546874 262226 547494 262294
rect 546874 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 547494 262226
rect 546874 262102 547494 262170
rect 546874 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 547494 262102
rect 546874 261978 547494 262046
rect 546874 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 547494 261978
rect 546874 244350 547494 261922
rect 546874 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 547494 244350
rect 546874 244226 547494 244294
rect 546874 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 547494 244226
rect 546874 244102 547494 244170
rect 546874 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 547494 244102
rect 546874 243978 547494 244046
rect 546874 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 547494 243978
rect 546874 226350 547494 243922
rect 546874 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 547494 226350
rect 546874 226226 547494 226294
rect 546874 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 547494 226226
rect 546874 226102 547494 226170
rect 546874 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 547494 226102
rect 546874 225978 547494 226046
rect 546874 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 547494 225978
rect 546874 208350 547494 225922
rect 546874 208294 546970 208350
rect 547026 208294 547094 208350
rect 547150 208294 547218 208350
rect 547274 208294 547342 208350
rect 547398 208294 547494 208350
rect 546874 208226 547494 208294
rect 546874 208170 546970 208226
rect 547026 208170 547094 208226
rect 547150 208170 547218 208226
rect 547274 208170 547342 208226
rect 547398 208170 547494 208226
rect 546874 208102 547494 208170
rect 546874 208046 546970 208102
rect 547026 208046 547094 208102
rect 547150 208046 547218 208102
rect 547274 208046 547342 208102
rect 547398 208046 547494 208102
rect 546874 207978 547494 208046
rect 546874 207922 546970 207978
rect 547026 207922 547094 207978
rect 547150 207922 547218 207978
rect 547274 207922 547342 207978
rect 547398 207922 547494 207978
rect 546874 190350 547494 207922
rect 546874 190294 546970 190350
rect 547026 190294 547094 190350
rect 547150 190294 547218 190350
rect 547274 190294 547342 190350
rect 547398 190294 547494 190350
rect 546874 190226 547494 190294
rect 546874 190170 546970 190226
rect 547026 190170 547094 190226
rect 547150 190170 547218 190226
rect 547274 190170 547342 190226
rect 547398 190170 547494 190226
rect 546874 190102 547494 190170
rect 546874 190046 546970 190102
rect 547026 190046 547094 190102
rect 547150 190046 547218 190102
rect 547274 190046 547342 190102
rect 547398 190046 547494 190102
rect 546874 189978 547494 190046
rect 546874 189922 546970 189978
rect 547026 189922 547094 189978
rect 547150 189922 547218 189978
rect 547274 189922 547342 189978
rect 547398 189922 547494 189978
rect 546874 172350 547494 189922
rect 546874 172294 546970 172350
rect 547026 172294 547094 172350
rect 547150 172294 547218 172350
rect 547274 172294 547342 172350
rect 547398 172294 547494 172350
rect 546874 172226 547494 172294
rect 546874 172170 546970 172226
rect 547026 172170 547094 172226
rect 547150 172170 547218 172226
rect 547274 172170 547342 172226
rect 547398 172170 547494 172226
rect 546874 172102 547494 172170
rect 546874 172046 546970 172102
rect 547026 172046 547094 172102
rect 547150 172046 547218 172102
rect 547274 172046 547342 172102
rect 547398 172046 547494 172102
rect 546874 171978 547494 172046
rect 546874 171922 546970 171978
rect 547026 171922 547094 171978
rect 547150 171922 547218 171978
rect 547274 171922 547342 171978
rect 547398 171922 547494 171978
rect 546874 154350 547494 171922
rect 546874 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 547494 154350
rect 546874 154226 547494 154294
rect 546874 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 547494 154226
rect 546874 154102 547494 154170
rect 546874 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 547494 154102
rect 546874 153978 547494 154046
rect 546874 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 547494 153978
rect 546874 136350 547494 153922
rect 546874 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 547494 136350
rect 546874 136226 547494 136294
rect 546874 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 547494 136226
rect 546874 136102 547494 136170
rect 546874 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 547494 136102
rect 546874 135978 547494 136046
rect 546874 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 547494 135978
rect 546874 118350 547494 135922
rect 546874 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 547494 118350
rect 546874 118226 547494 118294
rect 546874 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 547494 118226
rect 546874 118102 547494 118170
rect 546874 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 547494 118102
rect 546874 117978 547494 118046
rect 546874 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 547494 117978
rect 546874 100350 547494 117922
rect 546874 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 547494 100350
rect 546874 100226 547494 100294
rect 546874 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 547494 100226
rect 546874 100102 547494 100170
rect 546874 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 547494 100102
rect 546874 99978 547494 100046
rect 546874 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 547494 99978
rect 546874 82350 547494 99922
rect 546874 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 547494 82350
rect 546874 82226 547494 82294
rect 546874 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 547494 82226
rect 546874 82102 547494 82170
rect 546874 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 547494 82102
rect 546874 81978 547494 82046
rect 546874 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 547494 81978
rect 546874 64350 547494 81922
rect 546874 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 547494 64350
rect 546874 64226 547494 64294
rect 546874 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 547494 64226
rect 546874 64102 547494 64170
rect 546874 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 547494 64102
rect 546874 63978 547494 64046
rect 546874 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 547494 63978
rect 546874 46350 547494 63922
rect 546874 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 547494 46350
rect 546874 46226 547494 46294
rect 546874 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 547494 46226
rect 546874 46102 547494 46170
rect 546874 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 547494 46102
rect 546874 45978 547494 46046
rect 546874 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 547494 45978
rect 546874 28350 547494 45922
rect 546874 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 547494 28350
rect 546874 28226 547494 28294
rect 546874 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 547494 28226
rect 546874 28102 547494 28170
rect 546874 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 547494 28102
rect 546874 27978 547494 28046
rect 546874 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 547494 27978
rect 546874 10350 547494 27922
rect 546874 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 547494 10350
rect 546874 10226 547494 10294
rect 546874 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 547494 10226
rect 546874 10102 547494 10170
rect 546874 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 547494 10102
rect 546874 9978 547494 10046
rect 546874 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 547494 9978
rect 546874 -1120 547494 9922
rect 546874 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 547494 -1120
rect 546874 -1244 547494 -1176
rect 546874 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 547494 -1244
rect 546874 -1368 547494 -1300
rect 546874 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 547494 -1368
rect 546874 -1492 547494 -1424
rect 546874 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 547494 -1492
rect 546874 -1644 547494 -1548
rect 561154 597212 561774 598268
rect 561154 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 561774 597212
rect 561154 597088 561774 597156
rect 561154 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 561774 597088
rect 561154 596964 561774 597032
rect 561154 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 561774 596964
rect 561154 596840 561774 596908
rect 561154 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 561774 596840
rect 561154 580350 561774 596784
rect 561154 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 561774 580350
rect 561154 580226 561774 580294
rect 561154 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 561774 580226
rect 561154 580102 561774 580170
rect 561154 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 561774 580102
rect 561154 579978 561774 580046
rect 561154 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 561774 579978
rect 561154 562350 561774 579922
rect 561154 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 561774 562350
rect 561154 562226 561774 562294
rect 561154 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 561774 562226
rect 561154 562102 561774 562170
rect 561154 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 561774 562102
rect 561154 561978 561774 562046
rect 561154 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 561774 561978
rect 561154 544350 561774 561922
rect 561154 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 561774 544350
rect 561154 544226 561774 544294
rect 561154 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 561774 544226
rect 561154 544102 561774 544170
rect 561154 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 561774 544102
rect 561154 543978 561774 544046
rect 561154 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 561774 543978
rect 561154 526350 561774 543922
rect 561154 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 561774 526350
rect 561154 526226 561774 526294
rect 561154 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 561774 526226
rect 561154 526102 561774 526170
rect 561154 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 561774 526102
rect 561154 525978 561774 526046
rect 561154 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 561774 525978
rect 561154 508350 561774 525922
rect 561154 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 561774 508350
rect 561154 508226 561774 508294
rect 561154 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 561774 508226
rect 561154 508102 561774 508170
rect 561154 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 561774 508102
rect 561154 507978 561774 508046
rect 561154 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 561774 507978
rect 561154 490350 561774 507922
rect 561154 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 561774 490350
rect 561154 490226 561774 490294
rect 561154 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 561774 490226
rect 561154 490102 561774 490170
rect 561154 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 561774 490102
rect 561154 489978 561774 490046
rect 561154 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 561774 489978
rect 561154 472350 561774 489922
rect 561154 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 561774 472350
rect 561154 472226 561774 472294
rect 561154 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 561774 472226
rect 561154 472102 561774 472170
rect 561154 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 561774 472102
rect 561154 471978 561774 472046
rect 561154 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 561774 471978
rect 561154 454350 561774 471922
rect 561154 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 561774 454350
rect 561154 454226 561774 454294
rect 561154 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 561774 454226
rect 561154 454102 561774 454170
rect 561154 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 561774 454102
rect 561154 453978 561774 454046
rect 561154 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 561774 453978
rect 561154 436350 561774 453922
rect 561154 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 561774 436350
rect 561154 436226 561774 436294
rect 561154 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 561774 436226
rect 561154 436102 561774 436170
rect 561154 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 561774 436102
rect 561154 435978 561774 436046
rect 561154 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 561774 435978
rect 561154 418350 561774 435922
rect 561154 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 561774 418350
rect 561154 418226 561774 418294
rect 561154 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 561774 418226
rect 561154 418102 561774 418170
rect 561154 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 561774 418102
rect 561154 417978 561774 418046
rect 561154 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 561774 417978
rect 561154 400350 561774 417922
rect 561154 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 561774 400350
rect 561154 400226 561774 400294
rect 561154 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 561774 400226
rect 561154 400102 561774 400170
rect 561154 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 561774 400102
rect 561154 399978 561774 400046
rect 561154 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 561774 399978
rect 561154 382350 561774 399922
rect 561154 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 561774 382350
rect 561154 382226 561774 382294
rect 561154 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 561774 382226
rect 561154 382102 561774 382170
rect 561154 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 561774 382102
rect 561154 381978 561774 382046
rect 561154 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 561774 381978
rect 561154 364350 561774 381922
rect 561154 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 561774 364350
rect 561154 364226 561774 364294
rect 561154 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 561774 364226
rect 561154 364102 561774 364170
rect 561154 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 561774 364102
rect 561154 363978 561774 364046
rect 561154 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 561774 363978
rect 561154 346350 561774 363922
rect 561154 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 561774 346350
rect 561154 346226 561774 346294
rect 561154 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 561774 346226
rect 561154 346102 561774 346170
rect 561154 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 561774 346102
rect 561154 345978 561774 346046
rect 561154 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 561774 345978
rect 561154 328350 561774 345922
rect 561154 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 561774 328350
rect 561154 328226 561774 328294
rect 561154 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 561774 328226
rect 561154 328102 561774 328170
rect 561154 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 561774 328102
rect 561154 327978 561774 328046
rect 561154 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 561774 327978
rect 561154 310350 561774 327922
rect 561154 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 561774 310350
rect 561154 310226 561774 310294
rect 561154 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 561774 310226
rect 561154 310102 561774 310170
rect 561154 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 561774 310102
rect 561154 309978 561774 310046
rect 561154 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 561774 309978
rect 561154 292350 561774 309922
rect 561154 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 561774 292350
rect 561154 292226 561774 292294
rect 561154 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 561774 292226
rect 561154 292102 561774 292170
rect 561154 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 561774 292102
rect 561154 291978 561774 292046
rect 561154 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 561774 291978
rect 561154 274350 561774 291922
rect 561154 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 561774 274350
rect 561154 274226 561774 274294
rect 561154 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 561774 274226
rect 561154 274102 561774 274170
rect 561154 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 561774 274102
rect 561154 273978 561774 274046
rect 561154 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 561774 273978
rect 561154 256350 561774 273922
rect 561154 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 561774 256350
rect 561154 256226 561774 256294
rect 561154 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 561774 256226
rect 561154 256102 561774 256170
rect 561154 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 561774 256102
rect 561154 255978 561774 256046
rect 561154 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 561774 255978
rect 561154 238350 561774 255922
rect 561154 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 561774 238350
rect 561154 238226 561774 238294
rect 561154 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 561774 238226
rect 561154 238102 561774 238170
rect 561154 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 561774 238102
rect 561154 237978 561774 238046
rect 561154 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 561774 237978
rect 561154 220350 561774 237922
rect 561154 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 561774 220350
rect 561154 220226 561774 220294
rect 561154 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 561774 220226
rect 561154 220102 561774 220170
rect 561154 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 561774 220102
rect 561154 219978 561774 220046
rect 561154 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 561774 219978
rect 561154 202350 561774 219922
rect 561154 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 561774 202350
rect 561154 202226 561774 202294
rect 561154 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 561774 202226
rect 561154 202102 561774 202170
rect 561154 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 561774 202102
rect 561154 201978 561774 202046
rect 561154 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 561774 201978
rect 561154 184350 561774 201922
rect 561154 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 561774 184350
rect 561154 184226 561774 184294
rect 561154 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 561774 184226
rect 561154 184102 561774 184170
rect 561154 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 561774 184102
rect 561154 183978 561774 184046
rect 561154 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 561774 183978
rect 561154 166350 561774 183922
rect 561154 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 561774 166350
rect 561154 166226 561774 166294
rect 561154 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 561774 166226
rect 561154 166102 561774 166170
rect 561154 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 561774 166102
rect 561154 165978 561774 166046
rect 561154 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 561774 165978
rect 561154 148350 561774 165922
rect 561154 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 561774 148350
rect 561154 148226 561774 148294
rect 561154 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 561774 148226
rect 561154 148102 561774 148170
rect 561154 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 561774 148102
rect 561154 147978 561774 148046
rect 561154 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 561774 147978
rect 561154 130350 561774 147922
rect 561154 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 561774 130350
rect 561154 130226 561774 130294
rect 561154 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 561774 130226
rect 561154 130102 561774 130170
rect 561154 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 561774 130102
rect 561154 129978 561774 130046
rect 561154 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 561774 129978
rect 561154 112350 561774 129922
rect 561154 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 561774 112350
rect 561154 112226 561774 112294
rect 561154 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 561774 112226
rect 561154 112102 561774 112170
rect 561154 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 561774 112102
rect 561154 111978 561774 112046
rect 561154 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 561774 111978
rect 561154 94350 561774 111922
rect 561154 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 561774 94350
rect 561154 94226 561774 94294
rect 561154 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 561774 94226
rect 561154 94102 561774 94170
rect 561154 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 561774 94102
rect 561154 93978 561774 94046
rect 561154 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 561774 93978
rect 561154 76350 561774 93922
rect 561154 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 561774 76350
rect 561154 76226 561774 76294
rect 561154 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 561774 76226
rect 561154 76102 561774 76170
rect 561154 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 561774 76102
rect 561154 75978 561774 76046
rect 561154 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 561774 75978
rect 561154 58350 561774 75922
rect 561154 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 561774 58350
rect 561154 58226 561774 58294
rect 561154 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 561774 58226
rect 561154 58102 561774 58170
rect 561154 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 561774 58102
rect 561154 57978 561774 58046
rect 561154 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 561774 57978
rect 561154 40350 561774 57922
rect 561154 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 561774 40350
rect 561154 40226 561774 40294
rect 561154 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 561774 40226
rect 561154 40102 561774 40170
rect 561154 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 561774 40102
rect 561154 39978 561774 40046
rect 561154 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 561774 39978
rect 561154 22350 561774 39922
rect 561154 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 561774 22350
rect 561154 22226 561774 22294
rect 561154 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 561774 22226
rect 561154 22102 561774 22170
rect 561154 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 561774 22102
rect 561154 21978 561774 22046
rect 561154 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 561774 21978
rect 561154 4350 561774 21922
rect 561154 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 561774 4350
rect 561154 4226 561774 4294
rect 561154 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 561774 4226
rect 561154 4102 561774 4170
rect 561154 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 561774 4102
rect 561154 3978 561774 4046
rect 561154 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 561774 3978
rect 561154 -160 561774 3922
rect 561154 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 561774 -160
rect 561154 -284 561774 -216
rect 561154 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 561774 -284
rect 561154 -408 561774 -340
rect 561154 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 561774 -408
rect 561154 -532 561774 -464
rect 561154 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 561774 -532
rect 561154 -1644 561774 -588
rect 564874 598172 565494 598268
rect 564874 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 565494 598172
rect 564874 598048 565494 598116
rect 564874 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 565494 598048
rect 564874 597924 565494 597992
rect 564874 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 565494 597924
rect 564874 597800 565494 597868
rect 564874 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 565494 597800
rect 564874 586350 565494 597744
rect 564874 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 565494 586350
rect 564874 586226 565494 586294
rect 564874 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 565494 586226
rect 564874 586102 565494 586170
rect 564874 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 565494 586102
rect 564874 585978 565494 586046
rect 564874 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 565494 585978
rect 564874 568350 565494 585922
rect 564874 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 565494 568350
rect 564874 568226 565494 568294
rect 564874 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 565494 568226
rect 564874 568102 565494 568170
rect 564874 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 565494 568102
rect 564874 567978 565494 568046
rect 564874 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 565494 567978
rect 564874 550350 565494 567922
rect 564874 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 565494 550350
rect 564874 550226 565494 550294
rect 564874 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 565494 550226
rect 564874 550102 565494 550170
rect 564874 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 565494 550102
rect 564874 549978 565494 550046
rect 564874 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 565494 549978
rect 564874 532350 565494 549922
rect 564874 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 565494 532350
rect 564874 532226 565494 532294
rect 564874 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 565494 532226
rect 564874 532102 565494 532170
rect 564874 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 565494 532102
rect 564874 531978 565494 532046
rect 564874 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 565494 531978
rect 564874 514350 565494 531922
rect 564874 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 565494 514350
rect 564874 514226 565494 514294
rect 564874 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 565494 514226
rect 564874 514102 565494 514170
rect 564874 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 565494 514102
rect 564874 513978 565494 514046
rect 564874 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 565494 513978
rect 564874 496350 565494 513922
rect 564874 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 565494 496350
rect 564874 496226 565494 496294
rect 564874 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 565494 496226
rect 564874 496102 565494 496170
rect 564874 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 565494 496102
rect 564874 495978 565494 496046
rect 564874 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 565494 495978
rect 564874 478350 565494 495922
rect 564874 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 565494 478350
rect 564874 478226 565494 478294
rect 564874 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 565494 478226
rect 564874 478102 565494 478170
rect 564874 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 565494 478102
rect 564874 477978 565494 478046
rect 564874 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 565494 477978
rect 564874 460350 565494 477922
rect 564874 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 565494 460350
rect 564874 460226 565494 460294
rect 564874 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 565494 460226
rect 564874 460102 565494 460170
rect 564874 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 565494 460102
rect 564874 459978 565494 460046
rect 564874 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 565494 459978
rect 564874 442350 565494 459922
rect 564874 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 565494 442350
rect 564874 442226 565494 442294
rect 564874 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 565494 442226
rect 564874 442102 565494 442170
rect 564874 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 565494 442102
rect 564874 441978 565494 442046
rect 564874 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 565494 441978
rect 564874 424350 565494 441922
rect 564874 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 565494 424350
rect 564874 424226 565494 424294
rect 564874 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 565494 424226
rect 564874 424102 565494 424170
rect 564874 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 565494 424102
rect 564874 423978 565494 424046
rect 564874 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 565494 423978
rect 564874 406350 565494 423922
rect 564874 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 565494 406350
rect 564874 406226 565494 406294
rect 564874 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 565494 406226
rect 564874 406102 565494 406170
rect 564874 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 565494 406102
rect 564874 405978 565494 406046
rect 564874 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 565494 405978
rect 564874 388350 565494 405922
rect 564874 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 565494 388350
rect 564874 388226 565494 388294
rect 564874 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 565494 388226
rect 564874 388102 565494 388170
rect 564874 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 565494 388102
rect 564874 387978 565494 388046
rect 564874 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 565494 387978
rect 564874 370350 565494 387922
rect 564874 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 565494 370350
rect 564874 370226 565494 370294
rect 564874 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 565494 370226
rect 564874 370102 565494 370170
rect 564874 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 565494 370102
rect 564874 369978 565494 370046
rect 564874 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 565494 369978
rect 564874 352350 565494 369922
rect 564874 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 565494 352350
rect 564874 352226 565494 352294
rect 564874 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 565494 352226
rect 564874 352102 565494 352170
rect 564874 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 565494 352102
rect 564874 351978 565494 352046
rect 564874 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 565494 351978
rect 564874 334350 565494 351922
rect 564874 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 565494 334350
rect 564874 334226 565494 334294
rect 564874 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 565494 334226
rect 564874 334102 565494 334170
rect 564874 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 565494 334102
rect 564874 333978 565494 334046
rect 564874 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 565494 333978
rect 564874 316350 565494 333922
rect 564874 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 565494 316350
rect 564874 316226 565494 316294
rect 564874 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 565494 316226
rect 564874 316102 565494 316170
rect 564874 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 565494 316102
rect 564874 315978 565494 316046
rect 564874 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 565494 315978
rect 564874 298350 565494 315922
rect 564874 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 565494 298350
rect 564874 298226 565494 298294
rect 564874 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 565494 298226
rect 564874 298102 565494 298170
rect 564874 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 565494 298102
rect 564874 297978 565494 298046
rect 564874 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 565494 297978
rect 564874 280350 565494 297922
rect 564874 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 565494 280350
rect 564874 280226 565494 280294
rect 564874 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 565494 280226
rect 564874 280102 565494 280170
rect 564874 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 565494 280102
rect 564874 279978 565494 280046
rect 564874 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 565494 279978
rect 564874 262350 565494 279922
rect 564874 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 565494 262350
rect 564874 262226 565494 262294
rect 564874 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 565494 262226
rect 564874 262102 565494 262170
rect 564874 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 565494 262102
rect 564874 261978 565494 262046
rect 564874 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 565494 261978
rect 564874 244350 565494 261922
rect 564874 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 565494 244350
rect 564874 244226 565494 244294
rect 564874 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 565494 244226
rect 564874 244102 565494 244170
rect 564874 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 565494 244102
rect 564874 243978 565494 244046
rect 564874 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 565494 243978
rect 564874 226350 565494 243922
rect 564874 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 565494 226350
rect 564874 226226 565494 226294
rect 564874 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 565494 226226
rect 564874 226102 565494 226170
rect 564874 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 565494 226102
rect 564874 225978 565494 226046
rect 564874 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 565494 225978
rect 564874 208350 565494 225922
rect 564874 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 565494 208350
rect 564874 208226 565494 208294
rect 564874 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 565494 208226
rect 564874 208102 565494 208170
rect 564874 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 565494 208102
rect 564874 207978 565494 208046
rect 564874 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 565494 207978
rect 564874 190350 565494 207922
rect 564874 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 565494 190350
rect 564874 190226 565494 190294
rect 564874 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 565494 190226
rect 564874 190102 565494 190170
rect 564874 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 565494 190102
rect 564874 189978 565494 190046
rect 564874 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 565494 189978
rect 564874 172350 565494 189922
rect 564874 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 565494 172350
rect 564874 172226 565494 172294
rect 564874 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 565494 172226
rect 564874 172102 565494 172170
rect 564874 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 565494 172102
rect 564874 171978 565494 172046
rect 564874 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 565494 171978
rect 564874 154350 565494 171922
rect 564874 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 565494 154350
rect 564874 154226 565494 154294
rect 564874 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 565494 154226
rect 564874 154102 565494 154170
rect 564874 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 565494 154102
rect 564874 153978 565494 154046
rect 564874 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 565494 153978
rect 564874 136350 565494 153922
rect 564874 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 565494 136350
rect 564874 136226 565494 136294
rect 564874 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 565494 136226
rect 564874 136102 565494 136170
rect 564874 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 565494 136102
rect 564874 135978 565494 136046
rect 564874 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 565494 135978
rect 564874 118350 565494 135922
rect 564874 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 565494 118350
rect 564874 118226 565494 118294
rect 564874 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 565494 118226
rect 564874 118102 565494 118170
rect 564874 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 565494 118102
rect 564874 117978 565494 118046
rect 564874 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 565494 117978
rect 564874 100350 565494 117922
rect 564874 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 565494 100350
rect 564874 100226 565494 100294
rect 564874 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 565494 100226
rect 564874 100102 565494 100170
rect 564874 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 565494 100102
rect 564874 99978 565494 100046
rect 564874 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 565494 99978
rect 564874 82350 565494 99922
rect 564874 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 565494 82350
rect 564874 82226 565494 82294
rect 564874 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 565494 82226
rect 564874 82102 565494 82170
rect 564874 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 565494 82102
rect 564874 81978 565494 82046
rect 564874 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 565494 81978
rect 564874 64350 565494 81922
rect 564874 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 565494 64350
rect 564874 64226 565494 64294
rect 564874 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 565494 64226
rect 564874 64102 565494 64170
rect 564874 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 565494 64102
rect 564874 63978 565494 64046
rect 564874 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 565494 63978
rect 564874 46350 565494 63922
rect 564874 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 565494 46350
rect 564874 46226 565494 46294
rect 564874 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 565494 46226
rect 564874 46102 565494 46170
rect 564874 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 565494 46102
rect 564874 45978 565494 46046
rect 564874 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 565494 45978
rect 564874 28350 565494 45922
rect 564874 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 565494 28350
rect 564874 28226 565494 28294
rect 564874 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 565494 28226
rect 564874 28102 565494 28170
rect 564874 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 565494 28102
rect 564874 27978 565494 28046
rect 564874 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 565494 27978
rect 564874 10350 565494 27922
rect 564874 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 565494 10350
rect 564874 10226 565494 10294
rect 564874 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 565494 10226
rect 564874 10102 565494 10170
rect 564874 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 565494 10102
rect 564874 9978 565494 10046
rect 564874 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 565494 9978
rect 564874 -1120 565494 9922
rect 564874 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 565494 -1120
rect 564874 -1244 565494 -1176
rect 564874 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 565494 -1244
rect 564874 -1368 565494 -1300
rect 564874 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 565494 -1368
rect 564874 -1492 565494 -1424
rect 564874 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 565494 -1492
rect 564874 -1644 565494 -1548
rect 579154 597212 579774 598268
rect 579154 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 579774 597212
rect 579154 597088 579774 597156
rect 579154 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 579774 597088
rect 579154 596964 579774 597032
rect 579154 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 579774 596964
rect 579154 596840 579774 596908
rect 579154 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 579774 596840
rect 579154 580350 579774 596784
rect 579154 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 579774 580350
rect 579154 580226 579774 580294
rect 579154 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 579774 580226
rect 579154 580102 579774 580170
rect 579154 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 579774 580102
rect 579154 579978 579774 580046
rect 579154 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 579774 579978
rect 579154 562350 579774 579922
rect 579154 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 579774 562350
rect 579154 562226 579774 562294
rect 579154 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 579774 562226
rect 579154 562102 579774 562170
rect 579154 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 579774 562102
rect 579154 561978 579774 562046
rect 579154 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 579774 561978
rect 579154 544350 579774 561922
rect 579154 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 579774 544350
rect 579154 544226 579774 544294
rect 579154 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 579774 544226
rect 579154 544102 579774 544170
rect 579154 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 579774 544102
rect 579154 543978 579774 544046
rect 579154 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 579774 543978
rect 579154 526350 579774 543922
rect 579154 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 579774 526350
rect 579154 526226 579774 526294
rect 579154 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 579774 526226
rect 579154 526102 579774 526170
rect 579154 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 579774 526102
rect 579154 525978 579774 526046
rect 579154 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 579774 525978
rect 579154 508350 579774 525922
rect 579154 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 579774 508350
rect 579154 508226 579774 508294
rect 579154 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 579774 508226
rect 579154 508102 579774 508170
rect 579154 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 579774 508102
rect 579154 507978 579774 508046
rect 579154 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 579774 507978
rect 579154 490350 579774 507922
rect 579154 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 579774 490350
rect 579154 490226 579774 490294
rect 579154 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 579774 490226
rect 579154 490102 579774 490170
rect 579154 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 579774 490102
rect 579154 489978 579774 490046
rect 579154 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 579774 489978
rect 579154 472350 579774 489922
rect 579154 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 579774 472350
rect 579154 472226 579774 472294
rect 579154 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 579774 472226
rect 579154 472102 579774 472170
rect 579154 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 579774 472102
rect 579154 471978 579774 472046
rect 579154 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 579774 471978
rect 579154 454350 579774 471922
rect 579154 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 579774 454350
rect 579154 454226 579774 454294
rect 579154 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 579774 454226
rect 579154 454102 579774 454170
rect 579154 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 579774 454102
rect 579154 453978 579774 454046
rect 579154 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 579774 453978
rect 579154 436350 579774 453922
rect 579154 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 579774 436350
rect 579154 436226 579774 436294
rect 579154 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 579774 436226
rect 579154 436102 579774 436170
rect 579154 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 579774 436102
rect 579154 435978 579774 436046
rect 579154 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 579774 435978
rect 579154 418350 579774 435922
rect 579154 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 579774 418350
rect 579154 418226 579774 418294
rect 579154 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 579774 418226
rect 579154 418102 579774 418170
rect 579154 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 579774 418102
rect 579154 417978 579774 418046
rect 579154 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 579774 417978
rect 579154 400350 579774 417922
rect 579154 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 579774 400350
rect 579154 400226 579774 400294
rect 579154 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 579774 400226
rect 579154 400102 579774 400170
rect 579154 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 579774 400102
rect 579154 399978 579774 400046
rect 579154 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 579774 399978
rect 579154 382350 579774 399922
rect 579154 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 579774 382350
rect 579154 382226 579774 382294
rect 579154 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 579774 382226
rect 579154 382102 579774 382170
rect 579154 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 579774 382102
rect 579154 381978 579774 382046
rect 579154 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 579774 381978
rect 579154 364350 579774 381922
rect 579154 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 579774 364350
rect 579154 364226 579774 364294
rect 579154 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 579774 364226
rect 579154 364102 579774 364170
rect 579154 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 579774 364102
rect 579154 363978 579774 364046
rect 579154 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 579774 363978
rect 579154 346350 579774 363922
rect 579154 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 579774 346350
rect 579154 346226 579774 346294
rect 579154 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 579774 346226
rect 579154 346102 579774 346170
rect 579154 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 579774 346102
rect 579154 345978 579774 346046
rect 579154 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 579774 345978
rect 579154 328350 579774 345922
rect 579154 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 579774 328350
rect 579154 328226 579774 328294
rect 579154 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 579774 328226
rect 579154 328102 579774 328170
rect 579154 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 579774 328102
rect 579154 327978 579774 328046
rect 579154 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 579774 327978
rect 579154 310350 579774 327922
rect 579154 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 579774 310350
rect 579154 310226 579774 310294
rect 579154 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 579774 310226
rect 579154 310102 579774 310170
rect 579154 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 579774 310102
rect 579154 309978 579774 310046
rect 579154 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 579774 309978
rect 579154 292350 579774 309922
rect 579154 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 579774 292350
rect 579154 292226 579774 292294
rect 579154 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 579774 292226
rect 579154 292102 579774 292170
rect 579154 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 579774 292102
rect 579154 291978 579774 292046
rect 579154 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 579774 291978
rect 579154 274350 579774 291922
rect 579154 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 579774 274350
rect 579154 274226 579774 274294
rect 579154 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 579774 274226
rect 579154 274102 579774 274170
rect 579154 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 579774 274102
rect 579154 273978 579774 274046
rect 579154 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 579774 273978
rect 579154 256350 579774 273922
rect 579154 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 579774 256350
rect 579154 256226 579774 256294
rect 579154 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 579774 256226
rect 579154 256102 579774 256170
rect 579154 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 579774 256102
rect 579154 255978 579774 256046
rect 579154 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 579774 255978
rect 579154 238350 579774 255922
rect 579154 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 579774 238350
rect 579154 238226 579774 238294
rect 579154 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 579774 238226
rect 579154 238102 579774 238170
rect 579154 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 579774 238102
rect 579154 237978 579774 238046
rect 579154 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 579774 237978
rect 579154 220350 579774 237922
rect 579154 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 579774 220350
rect 579154 220226 579774 220294
rect 579154 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 579774 220226
rect 579154 220102 579774 220170
rect 579154 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 579774 220102
rect 579154 219978 579774 220046
rect 579154 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 579774 219978
rect 579154 202350 579774 219922
rect 579154 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 579774 202350
rect 579154 202226 579774 202294
rect 579154 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 579774 202226
rect 579154 202102 579774 202170
rect 579154 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 579774 202102
rect 579154 201978 579774 202046
rect 579154 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 579774 201978
rect 579154 184350 579774 201922
rect 579154 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 579774 184350
rect 579154 184226 579774 184294
rect 579154 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 579774 184226
rect 579154 184102 579774 184170
rect 579154 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 579774 184102
rect 579154 183978 579774 184046
rect 579154 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 579774 183978
rect 579154 166350 579774 183922
rect 579154 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 579774 166350
rect 579154 166226 579774 166294
rect 579154 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 579774 166226
rect 579154 166102 579774 166170
rect 579154 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 579774 166102
rect 579154 165978 579774 166046
rect 579154 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 579774 165978
rect 579154 148350 579774 165922
rect 579154 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 579774 148350
rect 579154 148226 579774 148294
rect 579154 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 579774 148226
rect 579154 148102 579774 148170
rect 579154 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 579774 148102
rect 579154 147978 579774 148046
rect 579154 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 579774 147978
rect 579154 130350 579774 147922
rect 579154 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 579774 130350
rect 579154 130226 579774 130294
rect 579154 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 579774 130226
rect 579154 130102 579774 130170
rect 579154 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 579774 130102
rect 579154 129978 579774 130046
rect 579154 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 579774 129978
rect 579154 112350 579774 129922
rect 579154 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 579774 112350
rect 579154 112226 579774 112294
rect 579154 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 579774 112226
rect 579154 112102 579774 112170
rect 579154 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 579774 112102
rect 579154 111978 579774 112046
rect 579154 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 579774 111978
rect 579154 94350 579774 111922
rect 579154 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 579774 94350
rect 579154 94226 579774 94294
rect 579154 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 579774 94226
rect 579154 94102 579774 94170
rect 579154 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 579774 94102
rect 579154 93978 579774 94046
rect 579154 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 579774 93978
rect 579154 76350 579774 93922
rect 579154 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 579774 76350
rect 579154 76226 579774 76294
rect 579154 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 579774 76226
rect 579154 76102 579774 76170
rect 579154 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 579774 76102
rect 579154 75978 579774 76046
rect 579154 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 579774 75978
rect 579154 58350 579774 75922
rect 579154 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 579774 58350
rect 579154 58226 579774 58294
rect 579154 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 579774 58226
rect 579154 58102 579774 58170
rect 579154 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 579774 58102
rect 579154 57978 579774 58046
rect 579154 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 579774 57978
rect 579154 40350 579774 57922
rect 579154 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 579774 40350
rect 579154 40226 579774 40294
rect 579154 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 579774 40226
rect 579154 40102 579774 40170
rect 579154 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 579774 40102
rect 579154 39978 579774 40046
rect 579154 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 579774 39978
rect 579154 22350 579774 39922
rect 579154 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 579774 22350
rect 579154 22226 579774 22294
rect 579154 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 579774 22226
rect 579154 22102 579774 22170
rect 579154 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 579774 22102
rect 579154 21978 579774 22046
rect 579154 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 579774 21978
rect 579154 4350 579774 21922
rect 579154 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 579774 4350
rect 579154 4226 579774 4294
rect 579154 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 579774 4226
rect 579154 4102 579774 4170
rect 579154 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 579774 4102
rect 579154 3978 579774 4046
rect 579154 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 579774 3978
rect 579154 -160 579774 3922
rect 579154 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 579774 -160
rect 579154 -284 579774 -216
rect 579154 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 579774 -284
rect 579154 -408 579774 -340
rect 579154 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 579774 -408
rect 579154 -532 579774 -464
rect 579154 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 579774 -532
rect 579154 -1644 579774 -588
rect 582874 598172 583494 598268
rect 582874 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 583494 598172
rect 582874 598048 583494 598116
rect 582874 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 583494 598048
rect 582874 597924 583494 597992
rect 582874 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 583494 597924
rect 582874 597800 583494 597868
rect 582874 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 583494 597800
rect 582874 586350 583494 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 582874 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 583494 586350
rect 582874 586226 583494 586294
rect 582874 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 583494 586226
rect 582874 586102 583494 586170
rect 582874 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 583494 586102
rect 582874 585978 583494 586046
rect 582874 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 583494 585978
rect 582874 568350 583494 585922
rect 582874 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 583494 568350
rect 582874 568226 583494 568294
rect 582874 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 583494 568226
rect 582874 568102 583494 568170
rect 582874 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 583494 568102
rect 582874 567978 583494 568046
rect 582874 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 583494 567978
rect 582874 550350 583494 567922
rect 582874 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 583494 550350
rect 582874 550226 583494 550294
rect 582874 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 583494 550226
rect 582874 550102 583494 550170
rect 582874 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 583494 550102
rect 582874 549978 583494 550046
rect 582874 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 583494 549978
rect 582874 532350 583494 549922
rect 582874 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 583494 532350
rect 582874 532226 583494 532294
rect 582874 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 583494 532226
rect 582874 532102 583494 532170
rect 582874 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 583494 532102
rect 582874 531978 583494 532046
rect 582874 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 583494 531978
rect 582874 514350 583494 531922
rect 582874 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 583494 514350
rect 582874 514226 583494 514294
rect 582874 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 583494 514226
rect 582874 514102 583494 514170
rect 582874 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 583494 514102
rect 582874 513978 583494 514046
rect 582874 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 583494 513978
rect 582874 496350 583494 513922
rect 582874 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 583494 496350
rect 582874 496226 583494 496294
rect 582874 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 583494 496226
rect 582874 496102 583494 496170
rect 582874 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 583494 496102
rect 582874 495978 583494 496046
rect 582874 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 583494 495978
rect 582874 478350 583494 495922
rect 582874 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 583494 478350
rect 582874 478226 583494 478294
rect 582874 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 583494 478226
rect 582874 478102 583494 478170
rect 582874 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 583494 478102
rect 582874 477978 583494 478046
rect 582874 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 583494 477978
rect 582874 460350 583494 477922
rect 582874 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 583494 460350
rect 582874 460226 583494 460294
rect 582874 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 583494 460226
rect 582874 460102 583494 460170
rect 582874 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 583494 460102
rect 582874 459978 583494 460046
rect 582874 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 583494 459978
rect 582874 442350 583494 459922
rect 582874 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 583494 442350
rect 582874 442226 583494 442294
rect 582874 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 583494 442226
rect 582874 442102 583494 442170
rect 582874 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 583494 442102
rect 582874 441978 583494 442046
rect 582874 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 583494 441978
rect 582874 424350 583494 441922
rect 582874 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 583494 424350
rect 582874 424226 583494 424294
rect 582874 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 583494 424226
rect 582874 424102 583494 424170
rect 582874 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 583494 424102
rect 582874 423978 583494 424046
rect 582874 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 583494 423978
rect 582874 406350 583494 423922
rect 582874 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 583494 406350
rect 582874 406226 583494 406294
rect 582874 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 583494 406226
rect 582874 406102 583494 406170
rect 582874 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 583494 406102
rect 582874 405978 583494 406046
rect 582874 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 583494 405978
rect 582874 388350 583494 405922
rect 582874 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 583494 388350
rect 582874 388226 583494 388294
rect 582874 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 583494 388226
rect 582874 388102 583494 388170
rect 582874 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 583494 388102
rect 582874 387978 583494 388046
rect 582874 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 583494 387978
rect 582874 370350 583494 387922
rect 582874 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 583494 370350
rect 582874 370226 583494 370294
rect 582874 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 583494 370226
rect 582874 370102 583494 370170
rect 582874 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 583494 370102
rect 582874 369978 583494 370046
rect 582874 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 583494 369978
rect 582874 352350 583494 369922
rect 582874 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 583494 352350
rect 582874 352226 583494 352294
rect 582874 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 583494 352226
rect 582874 352102 583494 352170
rect 582874 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 583494 352102
rect 582874 351978 583494 352046
rect 582874 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 583494 351978
rect 582874 334350 583494 351922
rect 582874 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 583494 334350
rect 582874 334226 583494 334294
rect 582874 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 583494 334226
rect 582874 334102 583494 334170
rect 582874 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 583494 334102
rect 582874 333978 583494 334046
rect 582874 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 583494 333978
rect 582874 316350 583494 333922
rect 582874 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 583494 316350
rect 582874 316226 583494 316294
rect 582874 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 583494 316226
rect 582874 316102 583494 316170
rect 582874 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 583494 316102
rect 582874 315978 583494 316046
rect 582874 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 583494 315978
rect 582874 298350 583494 315922
rect 582874 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 583494 298350
rect 582874 298226 583494 298294
rect 582874 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 583494 298226
rect 582874 298102 583494 298170
rect 582874 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 583494 298102
rect 582874 297978 583494 298046
rect 582874 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 583494 297978
rect 582874 280350 583494 297922
rect 582874 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 583494 280350
rect 582874 280226 583494 280294
rect 582874 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 583494 280226
rect 582874 280102 583494 280170
rect 582874 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 583494 280102
rect 582874 279978 583494 280046
rect 582874 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 583494 279978
rect 582874 262350 583494 279922
rect 582874 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 583494 262350
rect 582874 262226 583494 262294
rect 582874 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 583494 262226
rect 582874 262102 583494 262170
rect 582874 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 583494 262102
rect 582874 261978 583494 262046
rect 582874 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 583494 261978
rect 582874 244350 583494 261922
rect 582874 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 583494 244350
rect 582874 244226 583494 244294
rect 582874 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 583494 244226
rect 582874 244102 583494 244170
rect 582874 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 583494 244102
rect 582874 243978 583494 244046
rect 582874 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 583494 243978
rect 582874 226350 583494 243922
rect 582874 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 583494 226350
rect 582874 226226 583494 226294
rect 582874 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 583494 226226
rect 582874 226102 583494 226170
rect 582874 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 583494 226102
rect 582874 225978 583494 226046
rect 582874 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 583494 225978
rect 582874 208350 583494 225922
rect 582874 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 583494 208350
rect 582874 208226 583494 208294
rect 582874 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 583494 208226
rect 582874 208102 583494 208170
rect 582874 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 583494 208102
rect 582874 207978 583494 208046
rect 582874 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 583494 207978
rect 582874 190350 583494 207922
rect 582874 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 583494 190350
rect 582874 190226 583494 190294
rect 582874 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 583494 190226
rect 582874 190102 583494 190170
rect 582874 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 583494 190102
rect 582874 189978 583494 190046
rect 582874 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 583494 189978
rect 582874 172350 583494 189922
rect 582874 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 583494 172350
rect 582874 172226 583494 172294
rect 582874 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 583494 172226
rect 582874 172102 583494 172170
rect 582874 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 583494 172102
rect 582874 171978 583494 172046
rect 582874 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 583494 171978
rect 582874 154350 583494 171922
rect 582874 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 583494 154350
rect 582874 154226 583494 154294
rect 582874 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 583494 154226
rect 582874 154102 583494 154170
rect 582874 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 583494 154102
rect 582874 153978 583494 154046
rect 582874 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 583494 153978
rect 582874 136350 583494 153922
rect 582874 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 583494 136350
rect 582874 136226 583494 136294
rect 582874 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 583494 136226
rect 582874 136102 583494 136170
rect 582874 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 583494 136102
rect 582874 135978 583494 136046
rect 582874 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 583494 135978
rect 582874 118350 583494 135922
rect 582874 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 583494 118350
rect 582874 118226 583494 118294
rect 582874 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 583494 118226
rect 582874 118102 583494 118170
rect 582874 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 583494 118102
rect 582874 117978 583494 118046
rect 582874 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 583494 117978
rect 582874 100350 583494 117922
rect 582874 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 583494 100350
rect 582874 100226 583494 100294
rect 582874 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 583494 100226
rect 582874 100102 583494 100170
rect 582874 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 583494 100102
rect 582874 99978 583494 100046
rect 582874 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 583494 99978
rect 582874 82350 583494 99922
rect 582874 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 583494 82350
rect 582874 82226 583494 82294
rect 582874 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 583494 82226
rect 582874 82102 583494 82170
rect 582874 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 583494 82102
rect 582874 81978 583494 82046
rect 582874 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 583494 81978
rect 582874 64350 583494 81922
rect 582874 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 583494 64350
rect 582874 64226 583494 64294
rect 582874 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 583494 64226
rect 582874 64102 583494 64170
rect 582874 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 583494 64102
rect 582874 63978 583494 64046
rect 582874 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 583494 63978
rect 582874 46350 583494 63922
rect 582874 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 583494 46350
rect 582874 46226 583494 46294
rect 582874 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 583494 46226
rect 582874 46102 583494 46170
rect 582874 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 583494 46102
rect 582874 45978 583494 46046
rect 582874 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 583494 45978
rect 582874 28350 583494 45922
rect 582874 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 583494 28350
rect 582874 28226 583494 28294
rect 582874 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 583494 28226
rect 582874 28102 583494 28170
rect 582874 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 583494 28102
rect 582874 27978 583494 28046
rect 582874 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 583494 27978
rect 582874 10350 583494 27922
rect 582874 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 583494 10350
rect 582874 10226 583494 10294
rect 582874 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 583494 10226
rect 582874 10102 583494 10170
rect 582874 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 583494 10102
rect 582874 9978 583494 10046
rect 582874 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 583494 9978
rect 582874 -1120 583494 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 582874 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 583494 -1120
rect 582874 -1244 583494 -1176
rect 582874 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 583494 -1244
rect 582874 -1368 583494 -1300
rect 582874 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 583494 -1368
rect 582874 -1492 583494 -1424
rect 582874 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 583494 -1492
rect 582874 -1644 583494 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 3250 597156 3306 597212
rect 3374 597156 3430 597212
rect 3498 597156 3554 597212
rect 3622 597156 3678 597212
rect 3250 597032 3306 597088
rect 3374 597032 3430 597088
rect 3498 597032 3554 597088
rect 3622 597032 3678 597088
rect 3250 596908 3306 596964
rect 3374 596908 3430 596964
rect 3498 596908 3554 596964
rect 3622 596908 3678 596964
rect 3250 596784 3306 596840
rect 3374 596784 3430 596840
rect 3498 596784 3554 596840
rect 3622 596784 3678 596840
rect 3250 580294 3306 580350
rect 3374 580294 3430 580350
rect 3498 580294 3554 580350
rect 3622 580294 3678 580350
rect 3250 580170 3306 580226
rect 3374 580170 3430 580226
rect 3498 580170 3554 580226
rect 3622 580170 3678 580226
rect 3250 580046 3306 580102
rect 3374 580046 3430 580102
rect 3498 580046 3554 580102
rect 3622 580046 3678 580102
rect 3250 579922 3306 579978
rect 3374 579922 3430 579978
rect 3498 579922 3554 579978
rect 3622 579922 3678 579978
rect 3250 562294 3306 562350
rect 3374 562294 3430 562350
rect 3498 562294 3554 562350
rect 3622 562294 3678 562350
rect 3250 562170 3306 562226
rect 3374 562170 3430 562226
rect 3498 562170 3554 562226
rect 3622 562170 3678 562226
rect 3250 562046 3306 562102
rect 3374 562046 3430 562102
rect 3498 562046 3554 562102
rect 3622 562046 3678 562102
rect 3250 561922 3306 561978
rect 3374 561922 3430 561978
rect 3498 561922 3554 561978
rect 3622 561922 3678 561978
rect 3250 544294 3306 544350
rect 3374 544294 3430 544350
rect 3498 544294 3554 544350
rect 3622 544294 3678 544350
rect 3250 544170 3306 544226
rect 3374 544170 3430 544226
rect 3498 544170 3554 544226
rect 3622 544170 3678 544226
rect 3250 544046 3306 544102
rect 3374 544046 3430 544102
rect 3498 544046 3554 544102
rect 3622 544046 3678 544102
rect 3250 543922 3306 543978
rect 3374 543922 3430 543978
rect 3498 543922 3554 543978
rect 3622 543922 3678 543978
rect 3250 526294 3306 526350
rect 3374 526294 3430 526350
rect 3498 526294 3554 526350
rect 3622 526294 3678 526350
rect 3250 526170 3306 526226
rect 3374 526170 3430 526226
rect 3498 526170 3554 526226
rect 3622 526170 3678 526226
rect 3250 526046 3306 526102
rect 3374 526046 3430 526102
rect 3498 526046 3554 526102
rect 3622 526046 3678 526102
rect 3250 525922 3306 525978
rect 3374 525922 3430 525978
rect 3498 525922 3554 525978
rect 3622 525922 3678 525978
rect 3250 508294 3306 508350
rect 3374 508294 3430 508350
rect 3498 508294 3554 508350
rect 3622 508294 3678 508350
rect 3250 508170 3306 508226
rect 3374 508170 3430 508226
rect 3498 508170 3554 508226
rect 3622 508170 3678 508226
rect 3250 508046 3306 508102
rect 3374 508046 3430 508102
rect 3498 508046 3554 508102
rect 3622 508046 3678 508102
rect 3250 507922 3306 507978
rect 3374 507922 3430 507978
rect 3498 507922 3554 507978
rect 3622 507922 3678 507978
rect 3250 490294 3306 490350
rect 3374 490294 3430 490350
rect 3498 490294 3554 490350
rect 3622 490294 3678 490350
rect 3250 490170 3306 490226
rect 3374 490170 3430 490226
rect 3498 490170 3554 490226
rect 3622 490170 3678 490226
rect 3250 490046 3306 490102
rect 3374 490046 3430 490102
rect 3498 490046 3554 490102
rect 3622 490046 3678 490102
rect 3250 489922 3306 489978
rect 3374 489922 3430 489978
rect 3498 489922 3554 489978
rect 3622 489922 3678 489978
rect 3250 472294 3306 472350
rect 3374 472294 3430 472350
rect 3498 472294 3554 472350
rect 3622 472294 3678 472350
rect 3250 472170 3306 472226
rect 3374 472170 3430 472226
rect 3498 472170 3554 472226
rect 3622 472170 3678 472226
rect 3250 472046 3306 472102
rect 3374 472046 3430 472102
rect 3498 472046 3554 472102
rect 3622 472046 3678 472102
rect 3250 471922 3306 471978
rect 3374 471922 3430 471978
rect 3498 471922 3554 471978
rect 3622 471922 3678 471978
rect 3250 454294 3306 454350
rect 3374 454294 3430 454350
rect 3498 454294 3554 454350
rect 3622 454294 3678 454350
rect 3250 454170 3306 454226
rect 3374 454170 3430 454226
rect 3498 454170 3554 454226
rect 3622 454170 3678 454226
rect 3250 454046 3306 454102
rect 3374 454046 3430 454102
rect 3498 454046 3554 454102
rect 3622 454046 3678 454102
rect 3250 453922 3306 453978
rect 3374 453922 3430 453978
rect 3498 453922 3554 453978
rect 3622 453922 3678 453978
rect 3250 436294 3306 436350
rect 3374 436294 3430 436350
rect 3498 436294 3554 436350
rect 3622 436294 3678 436350
rect 3250 436170 3306 436226
rect 3374 436170 3430 436226
rect 3498 436170 3554 436226
rect 3622 436170 3678 436226
rect 3250 436046 3306 436102
rect 3374 436046 3430 436102
rect 3498 436046 3554 436102
rect 3622 436046 3678 436102
rect 3250 435922 3306 435978
rect 3374 435922 3430 435978
rect 3498 435922 3554 435978
rect 3622 435922 3678 435978
rect 3250 418294 3306 418350
rect 3374 418294 3430 418350
rect 3498 418294 3554 418350
rect 3622 418294 3678 418350
rect 3250 418170 3306 418226
rect 3374 418170 3430 418226
rect 3498 418170 3554 418226
rect 3622 418170 3678 418226
rect 3250 418046 3306 418102
rect 3374 418046 3430 418102
rect 3498 418046 3554 418102
rect 3622 418046 3678 418102
rect 3250 417922 3306 417978
rect 3374 417922 3430 417978
rect 3498 417922 3554 417978
rect 3622 417922 3678 417978
rect 3250 400294 3306 400350
rect 3374 400294 3430 400350
rect 3498 400294 3554 400350
rect 3622 400294 3678 400350
rect 3250 400170 3306 400226
rect 3374 400170 3430 400226
rect 3498 400170 3554 400226
rect 3622 400170 3678 400226
rect 3250 400046 3306 400102
rect 3374 400046 3430 400102
rect 3498 400046 3554 400102
rect 3622 400046 3678 400102
rect 3250 399922 3306 399978
rect 3374 399922 3430 399978
rect 3498 399922 3554 399978
rect 3622 399922 3678 399978
rect 3250 382294 3306 382350
rect 3374 382294 3430 382350
rect 3498 382294 3554 382350
rect 3622 382294 3678 382350
rect 3250 382170 3306 382226
rect 3374 382170 3430 382226
rect 3498 382170 3554 382226
rect 3622 382170 3678 382226
rect 3250 382046 3306 382102
rect 3374 382046 3430 382102
rect 3498 382046 3554 382102
rect 3622 382046 3678 382102
rect 3250 381922 3306 381978
rect 3374 381922 3430 381978
rect 3498 381922 3554 381978
rect 3622 381922 3678 381978
rect 3250 364294 3306 364350
rect 3374 364294 3430 364350
rect 3498 364294 3554 364350
rect 3622 364294 3678 364350
rect 3250 364170 3306 364226
rect 3374 364170 3430 364226
rect 3498 364170 3554 364226
rect 3622 364170 3678 364226
rect 3250 364046 3306 364102
rect 3374 364046 3430 364102
rect 3498 364046 3554 364102
rect 3622 364046 3678 364102
rect 3250 363922 3306 363978
rect 3374 363922 3430 363978
rect 3498 363922 3554 363978
rect 3622 363922 3678 363978
rect 3250 346294 3306 346350
rect 3374 346294 3430 346350
rect 3498 346294 3554 346350
rect 3622 346294 3678 346350
rect 3250 346170 3306 346226
rect 3374 346170 3430 346226
rect 3498 346170 3554 346226
rect 3622 346170 3678 346226
rect 3250 346046 3306 346102
rect 3374 346046 3430 346102
rect 3498 346046 3554 346102
rect 3622 346046 3678 346102
rect 3250 345922 3306 345978
rect 3374 345922 3430 345978
rect 3498 345922 3554 345978
rect 3622 345922 3678 345978
rect 3250 328294 3306 328350
rect 3374 328294 3430 328350
rect 3498 328294 3554 328350
rect 3622 328294 3678 328350
rect 3250 328170 3306 328226
rect 3374 328170 3430 328226
rect 3498 328170 3554 328226
rect 3622 328170 3678 328226
rect 3250 328046 3306 328102
rect 3374 328046 3430 328102
rect 3498 328046 3554 328102
rect 3622 328046 3678 328102
rect 3250 327922 3306 327978
rect 3374 327922 3430 327978
rect 3498 327922 3554 327978
rect 3622 327922 3678 327978
rect 3250 310294 3306 310350
rect 3374 310294 3430 310350
rect 3498 310294 3554 310350
rect 3622 310294 3678 310350
rect 3250 310170 3306 310226
rect 3374 310170 3430 310226
rect 3498 310170 3554 310226
rect 3622 310170 3678 310226
rect 3250 310046 3306 310102
rect 3374 310046 3430 310102
rect 3498 310046 3554 310102
rect 3622 310046 3678 310102
rect 3250 309922 3306 309978
rect 3374 309922 3430 309978
rect 3498 309922 3554 309978
rect 3622 309922 3678 309978
rect 3250 292294 3306 292350
rect 3374 292294 3430 292350
rect 3498 292294 3554 292350
rect 3622 292294 3678 292350
rect 3250 292170 3306 292226
rect 3374 292170 3430 292226
rect 3498 292170 3554 292226
rect 3622 292170 3678 292226
rect 3250 292046 3306 292102
rect 3374 292046 3430 292102
rect 3498 292046 3554 292102
rect 3622 292046 3678 292102
rect 3250 291922 3306 291978
rect 3374 291922 3430 291978
rect 3498 291922 3554 291978
rect 3622 291922 3678 291978
rect 3250 274294 3306 274350
rect 3374 274294 3430 274350
rect 3498 274294 3554 274350
rect 3622 274294 3678 274350
rect 3250 274170 3306 274226
rect 3374 274170 3430 274226
rect 3498 274170 3554 274226
rect 3622 274170 3678 274226
rect 3250 274046 3306 274102
rect 3374 274046 3430 274102
rect 3498 274046 3554 274102
rect 3622 274046 3678 274102
rect 3250 273922 3306 273978
rect 3374 273922 3430 273978
rect 3498 273922 3554 273978
rect 3622 273922 3678 273978
rect 3250 256294 3306 256350
rect 3374 256294 3430 256350
rect 3498 256294 3554 256350
rect 3622 256294 3678 256350
rect 3250 256170 3306 256226
rect 3374 256170 3430 256226
rect 3498 256170 3554 256226
rect 3622 256170 3678 256226
rect 3250 256046 3306 256102
rect 3374 256046 3430 256102
rect 3498 256046 3554 256102
rect 3622 256046 3678 256102
rect 3250 255922 3306 255978
rect 3374 255922 3430 255978
rect 3498 255922 3554 255978
rect 3622 255922 3678 255978
rect 3250 238294 3306 238350
rect 3374 238294 3430 238350
rect 3498 238294 3554 238350
rect 3622 238294 3678 238350
rect 3250 238170 3306 238226
rect 3374 238170 3430 238226
rect 3498 238170 3554 238226
rect 3622 238170 3678 238226
rect 3250 238046 3306 238102
rect 3374 238046 3430 238102
rect 3498 238046 3554 238102
rect 3622 238046 3678 238102
rect 3250 237922 3306 237978
rect 3374 237922 3430 237978
rect 3498 237922 3554 237978
rect 3622 237922 3678 237978
rect 3250 220294 3306 220350
rect 3374 220294 3430 220350
rect 3498 220294 3554 220350
rect 3622 220294 3678 220350
rect 3250 220170 3306 220226
rect 3374 220170 3430 220226
rect 3498 220170 3554 220226
rect 3622 220170 3678 220226
rect 3250 220046 3306 220102
rect 3374 220046 3430 220102
rect 3498 220046 3554 220102
rect 3622 220046 3678 220102
rect 3250 219922 3306 219978
rect 3374 219922 3430 219978
rect 3498 219922 3554 219978
rect 3622 219922 3678 219978
rect 3250 202294 3306 202350
rect 3374 202294 3430 202350
rect 3498 202294 3554 202350
rect 3622 202294 3678 202350
rect 3250 202170 3306 202226
rect 3374 202170 3430 202226
rect 3498 202170 3554 202226
rect 3622 202170 3678 202226
rect 3250 202046 3306 202102
rect 3374 202046 3430 202102
rect 3498 202046 3554 202102
rect 3622 202046 3678 202102
rect 3250 201922 3306 201978
rect 3374 201922 3430 201978
rect 3498 201922 3554 201978
rect 3622 201922 3678 201978
rect 3250 184294 3306 184350
rect 3374 184294 3430 184350
rect 3498 184294 3554 184350
rect 3622 184294 3678 184350
rect 3250 184170 3306 184226
rect 3374 184170 3430 184226
rect 3498 184170 3554 184226
rect 3622 184170 3678 184226
rect 3250 184046 3306 184102
rect 3374 184046 3430 184102
rect 3498 184046 3554 184102
rect 3622 184046 3678 184102
rect 3250 183922 3306 183978
rect 3374 183922 3430 183978
rect 3498 183922 3554 183978
rect 3622 183922 3678 183978
rect 3250 166294 3306 166350
rect 3374 166294 3430 166350
rect 3498 166294 3554 166350
rect 3622 166294 3678 166350
rect 3250 166170 3306 166226
rect 3374 166170 3430 166226
rect 3498 166170 3554 166226
rect 3622 166170 3678 166226
rect 3250 166046 3306 166102
rect 3374 166046 3430 166102
rect 3498 166046 3554 166102
rect 3622 166046 3678 166102
rect 3250 165922 3306 165978
rect 3374 165922 3430 165978
rect 3498 165922 3554 165978
rect 3622 165922 3678 165978
rect 3250 148294 3306 148350
rect 3374 148294 3430 148350
rect 3498 148294 3554 148350
rect 3622 148294 3678 148350
rect 3250 148170 3306 148226
rect 3374 148170 3430 148226
rect 3498 148170 3554 148226
rect 3622 148170 3678 148226
rect 3250 148046 3306 148102
rect 3374 148046 3430 148102
rect 3498 148046 3554 148102
rect 3622 148046 3678 148102
rect 3250 147922 3306 147978
rect 3374 147922 3430 147978
rect 3498 147922 3554 147978
rect 3622 147922 3678 147978
rect 3250 130294 3306 130350
rect 3374 130294 3430 130350
rect 3498 130294 3554 130350
rect 3622 130294 3678 130350
rect 3250 130170 3306 130226
rect 3374 130170 3430 130226
rect 3498 130170 3554 130226
rect 3622 130170 3678 130226
rect 3250 130046 3306 130102
rect 3374 130046 3430 130102
rect 3498 130046 3554 130102
rect 3622 130046 3678 130102
rect 3250 129922 3306 129978
rect 3374 129922 3430 129978
rect 3498 129922 3554 129978
rect 3622 129922 3678 129978
rect 3250 112294 3306 112350
rect 3374 112294 3430 112350
rect 3498 112294 3554 112350
rect 3622 112294 3678 112350
rect 3250 112170 3306 112226
rect 3374 112170 3430 112226
rect 3498 112170 3554 112226
rect 3622 112170 3678 112226
rect 3250 112046 3306 112102
rect 3374 112046 3430 112102
rect 3498 112046 3554 112102
rect 3622 112046 3678 112102
rect 3250 111922 3306 111978
rect 3374 111922 3430 111978
rect 3498 111922 3554 111978
rect 3622 111922 3678 111978
rect 3250 94294 3306 94350
rect 3374 94294 3430 94350
rect 3498 94294 3554 94350
rect 3622 94294 3678 94350
rect 3250 94170 3306 94226
rect 3374 94170 3430 94226
rect 3498 94170 3554 94226
rect 3622 94170 3678 94226
rect 3250 94046 3306 94102
rect 3374 94046 3430 94102
rect 3498 94046 3554 94102
rect 3622 94046 3678 94102
rect 3250 93922 3306 93978
rect 3374 93922 3430 93978
rect 3498 93922 3554 93978
rect 3622 93922 3678 93978
rect 3250 76294 3306 76350
rect 3374 76294 3430 76350
rect 3498 76294 3554 76350
rect 3622 76294 3678 76350
rect 3250 76170 3306 76226
rect 3374 76170 3430 76226
rect 3498 76170 3554 76226
rect 3622 76170 3678 76226
rect 3250 76046 3306 76102
rect 3374 76046 3430 76102
rect 3498 76046 3554 76102
rect 3622 76046 3678 76102
rect 3250 75922 3306 75978
rect 3374 75922 3430 75978
rect 3498 75922 3554 75978
rect 3622 75922 3678 75978
rect 3250 58294 3306 58350
rect 3374 58294 3430 58350
rect 3498 58294 3554 58350
rect 3622 58294 3678 58350
rect 3250 58170 3306 58226
rect 3374 58170 3430 58226
rect 3498 58170 3554 58226
rect 3622 58170 3678 58226
rect 3250 58046 3306 58102
rect 3374 58046 3430 58102
rect 3498 58046 3554 58102
rect 3622 58046 3678 58102
rect 3250 57922 3306 57978
rect 3374 57922 3430 57978
rect 3498 57922 3554 57978
rect 3622 57922 3678 57978
rect 3250 40294 3306 40350
rect 3374 40294 3430 40350
rect 3498 40294 3554 40350
rect 3622 40294 3678 40350
rect 3250 40170 3306 40226
rect 3374 40170 3430 40226
rect 3498 40170 3554 40226
rect 3622 40170 3678 40226
rect 3250 40046 3306 40102
rect 3374 40046 3430 40102
rect 3498 40046 3554 40102
rect 3622 40046 3678 40102
rect 3250 39922 3306 39978
rect 3374 39922 3430 39978
rect 3498 39922 3554 39978
rect 3622 39922 3678 39978
rect 3250 22294 3306 22350
rect 3374 22294 3430 22350
rect 3498 22294 3554 22350
rect 3622 22294 3678 22350
rect 3250 22170 3306 22226
rect 3374 22170 3430 22226
rect 3498 22170 3554 22226
rect 3622 22170 3678 22226
rect 3250 22046 3306 22102
rect 3374 22046 3430 22102
rect 3498 22046 3554 22102
rect 3622 22046 3678 22102
rect 3250 21922 3306 21978
rect 3374 21922 3430 21978
rect 3498 21922 3554 21978
rect 3622 21922 3678 21978
rect 3250 4294 3306 4350
rect 3374 4294 3430 4350
rect 3498 4294 3554 4350
rect 3622 4294 3678 4350
rect 3250 4170 3306 4226
rect 3374 4170 3430 4226
rect 3498 4170 3554 4226
rect 3622 4170 3678 4226
rect 3250 4046 3306 4102
rect 3374 4046 3430 4102
rect 3498 4046 3554 4102
rect 3622 4046 3678 4102
rect 3250 3922 3306 3978
rect 3374 3922 3430 3978
rect 3498 3922 3554 3978
rect 3622 3922 3678 3978
rect 3250 -216 3306 -160
rect 3374 -216 3430 -160
rect 3498 -216 3554 -160
rect 3622 -216 3678 -160
rect 3250 -340 3306 -284
rect 3374 -340 3430 -284
rect 3498 -340 3554 -284
rect 3622 -340 3678 -284
rect 3250 -464 3306 -408
rect 3374 -464 3430 -408
rect 3498 -464 3554 -408
rect 3622 -464 3678 -408
rect 3250 -588 3306 -532
rect 3374 -588 3430 -532
rect 3498 -588 3554 -532
rect 3622 -588 3678 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 6970 598116 7026 598172
rect 7094 598116 7150 598172
rect 7218 598116 7274 598172
rect 7342 598116 7398 598172
rect 6970 597992 7026 598048
rect 7094 597992 7150 598048
rect 7218 597992 7274 598048
rect 7342 597992 7398 598048
rect 6970 597868 7026 597924
rect 7094 597868 7150 597924
rect 7218 597868 7274 597924
rect 7342 597868 7398 597924
rect 6970 597744 7026 597800
rect 7094 597744 7150 597800
rect 7218 597744 7274 597800
rect 7342 597744 7398 597800
rect 6970 586294 7026 586350
rect 7094 586294 7150 586350
rect 7218 586294 7274 586350
rect 7342 586294 7398 586350
rect 6970 586170 7026 586226
rect 7094 586170 7150 586226
rect 7218 586170 7274 586226
rect 7342 586170 7398 586226
rect 6970 586046 7026 586102
rect 7094 586046 7150 586102
rect 7218 586046 7274 586102
rect 7342 586046 7398 586102
rect 6970 585922 7026 585978
rect 7094 585922 7150 585978
rect 7218 585922 7274 585978
rect 7342 585922 7398 585978
rect 6970 568294 7026 568350
rect 7094 568294 7150 568350
rect 7218 568294 7274 568350
rect 7342 568294 7398 568350
rect 6970 568170 7026 568226
rect 7094 568170 7150 568226
rect 7218 568170 7274 568226
rect 7342 568170 7398 568226
rect 6970 568046 7026 568102
rect 7094 568046 7150 568102
rect 7218 568046 7274 568102
rect 7342 568046 7398 568102
rect 6970 567922 7026 567978
rect 7094 567922 7150 567978
rect 7218 567922 7274 567978
rect 7342 567922 7398 567978
rect 6970 550294 7026 550350
rect 7094 550294 7150 550350
rect 7218 550294 7274 550350
rect 7342 550294 7398 550350
rect 6970 550170 7026 550226
rect 7094 550170 7150 550226
rect 7218 550170 7274 550226
rect 7342 550170 7398 550226
rect 6970 550046 7026 550102
rect 7094 550046 7150 550102
rect 7218 550046 7274 550102
rect 7342 550046 7398 550102
rect 6970 549922 7026 549978
rect 7094 549922 7150 549978
rect 7218 549922 7274 549978
rect 7342 549922 7398 549978
rect 6970 532294 7026 532350
rect 7094 532294 7150 532350
rect 7218 532294 7274 532350
rect 7342 532294 7398 532350
rect 6970 532170 7026 532226
rect 7094 532170 7150 532226
rect 7218 532170 7274 532226
rect 7342 532170 7398 532226
rect 6970 532046 7026 532102
rect 7094 532046 7150 532102
rect 7218 532046 7274 532102
rect 7342 532046 7398 532102
rect 6970 531922 7026 531978
rect 7094 531922 7150 531978
rect 7218 531922 7274 531978
rect 7342 531922 7398 531978
rect 6970 514294 7026 514350
rect 7094 514294 7150 514350
rect 7218 514294 7274 514350
rect 7342 514294 7398 514350
rect 6970 514170 7026 514226
rect 7094 514170 7150 514226
rect 7218 514170 7274 514226
rect 7342 514170 7398 514226
rect 6970 514046 7026 514102
rect 7094 514046 7150 514102
rect 7218 514046 7274 514102
rect 7342 514046 7398 514102
rect 6970 513922 7026 513978
rect 7094 513922 7150 513978
rect 7218 513922 7274 513978
rect 7342 513922 7398 513978
rect 6970 496294 7026 496350
rect 7094 496294 7150 496350
rect 7218 496294 7274 496350
rect 7342 496294 7398 496350
rect 6970 496170 7026 496226
rect 7094 496170 7150 496226
rect 7218 496170 7274 496226
rect 7342 496170 7398 496226
rect 6970 496046 7026 496102
rect 7094 496046 7150 496102
rect 7218 496046 7274 496102
rect 7342 496046 7398 496102
rect 6970 495922 7026 495978
rect 7094 495922 7150 495978
rect 7218 495922 7274 495978
rect 7342 495922 7398 495978
rect 6970 478294 7026 478350
rect 7094 478294 7150 478350
rect 7218 478294 7274 478350
rect 7342 478294 7398 478350
rect 6970 478170 7026 478226
rect 7094 478170 7150 478226
rect 7218 478170 7274 478226
rect 7342 478170 7398 478226
rect 6970 478046 7026 478102
rect 7094 478046 7150 478102
rect 7218 478046 7274 478102
rect 7342 478046 7398 478102
rect 6970 477922 7026 477978
rect 7094 477922 7150 477978
rect 7218 477922 7274 477978
rect 7342 477922 7398 477978
rect 6970 460294 7026 460350
rect 7094 460294 7150 460350
rect 7218 460294 7274 460350
rect 7342 460294 7398 460350
rect 6970 460170 7026 460226
rect 7094 460170 7150 460226
rect 7218 460170 7274 460226
rect 7342 460170 7398 460226
rect 6970 460046 7026 460102
rect 7094 460046 7150 460102
rect 7218 460046 7274 460102
rect 7342 460046 7398 460102
rect 6970 459922 7026 459978
rect 7094 459922 7150 459978
rect 7218 459922 7274 459978
rect 7342 459922 7398 459978
rect 6970 442294 7026 442350
rect 7094 442294 7150 442350
rect 7218 442294 7274 442350
rect 7342 442294 7398 442350
rect 6970 442170 7026 442226
rect 7094 442170 7150 442226
rect 7218 442170 7274 442226
rect 7342 442170 7398 442226
rect 6970 442046 7026 442102
rect 7094 442046 7150 442102
rect 7218 442046 7274 442102
rect 7342 442046 7398 442102
rect 6970 441922 7026 441978
rect 7094 441922 7150 441978
rect 7218 441922 7274 441978
rect 7342 441922 7398 441978
rect 6970 424294 7026 424350
rect 7094 424294 7150 424350
rect 7218 424294 7274 424350
rect 7342 424294 7398 424350
rect 6970 424170 7026 424226
rect 7094 424170 7150 424226
rect 7218 424170 7274 424226
rect 7342 424170 7398 424226
rect 6970 424046 7026 424102
rect 7094 424046 7150 424102
rect 7218 424046 7274 424102
rect 7342 424046 7398 424102
rect 6970 423922 7026 423978
rect 7094 423922 7150 423978
rect 7218 423922 7274 423978
rect 7342 423922 7398 423978
rect 6970 406294 7026 406350
rect 7094 406294 7150 406350
rect 7218 406294 7274 406350
rect 7342 406294 7398 406350
rect 6970 406170 7026 406226
rect 7094 406170 7150 406226
rect 7218 406170 7274 406226
rect 7342 406170 7398 406226
rect 6970 406046 7026 406102
rect 7094 406046 7150 406102
rect 7218 406046 7274 406102
rect 7342 406046 7398 406102
rect 6970 405922 7026 405978
rect 7094 405922 7150 405978
rect 7218 405922 7274 405978
rect 7342 405922 7398 405978
rect 6970 388294 7026 388350
rect 7094 388294 7150 388350
rect 7218 388294 7274 388350
rect 7342 388294 7398 388350
rect 6970 388170 7026 388226
rect 7094 388170 7150 388226
rect 7218 388170 7274 388226
rect 7342 388170 7398 388226
rect 6970 388046 7026 388102
rect 7094 388046 7150 388102
rect 7218 388046 7274 388102
rect 7342 388046 7398 388102
rect 6970 387922 7026 387978
rect 7094 387922 7150 387978
rect 7218 387922 7274 387978
rect 7342 387922 7398 387978
rect 6970 370294 7026 370350
rect 7094 370294 7150 370350
rect 7218 370294 7274 370350
rect 7342 370294 7398 370350
rect 6970 370170 7026 370226
rect 7094 370170 7150 370226
rect 7218 370170 7274 370226
rect 7342 370170 7398 370226
rect 6970 370046 7026 370102
rect 7094 370046 7150 370102
rect 7218 370046 7274 370102
rect 7342 370046 7398 370102
rect 6970 369922 7026 369978
rect 7094 369922 7150 369978
rect 7218 369922 7274 369978
rect 7342 369922 7398 369978
rect 6970 352294 7026 352350
rect 7094 352294 7150 352350
rect 7218 352294 7274 352350
rect 7342 352294 7398 352350
rect 6970 352170 7026 352226
rect 7094 352170 7150 352226
rect 7218 352170 7274 352226
rect 7342 352170 7398 352226
rect 6970 352046 7026 352102
rect 7094 352046 7150 352102
rect 7218 352046 7274 352102
rect 7342 352046 7398 352102
rect 6970 351922 7026 351978
rect 7094 351922 7150 351978
rect 7218 351922 7274 351978
rect 7342 351922 7398 351978
rect 6970 334294 7026 334350
rect 7094 334294 7150 334350
rect 7218 334294 7274 334350
rect 7342 334294 7398 334350
rect 6970 334170 7026 334226
rect 7094 334170 7150 334226
rect 7218 334170 7274 334226
rect 7342 334170 7398 334226
rect 6970 334046 7026 334102
rect 7094 334046 7150 334102
rect 7218 334046 7274 334102
rect 7342 334046 7398 334102
rect 6970 333922 7026 333978
rect 7094 333922 7150 333978
rect 7218 333922 7274 333978
rect 7342 333922 7398 333978
rect 6970 316294 7026 316350
rect 7094 316294 7150 316350
rect 7218 316294 7274 316350
rect 7342 316294 7398 316350
rect 6970 316170 7026 316226
rect 7094 316170 7150 316226
rect 7218 316170 7274 316226
rect 7342 316170 7398 316226
rect 6970 316046 7026 316102
rect 7094 316046 7150 316102
rect 7218 316046 7274 316102
rect 7342 316046 7398 316102
rect 6970 315922 7026 315978
rect 7094 315922 7150 315978
rect 7218 315922 7274 315978
rect 7342 315922 7398 315978
rect 6970 298294 7026 298350
rect 7094 298294 7150 298350
rect 7218 298294 7274 298350
rect 7342 298294 7398 298350
rect 6970 298170 7026 298226
rect 7094 298170 7150 298226
rect 7218 298170 7274 298226
rect 7342 298170 7398 298226
rect 6970 298046 7026 298102
rect 7094 298046 7150 298102
rect 7218 298046 7274 298102
rect 7342 298046 7398 298102
rect 6970 297922 7026 297978
rect 7094 297922 7150 297978
rect 7218 297922 7274 297978
rect 7342 297922 7398 297978
rect 6970 280294 7026 280350
rect 7094 280294 7150 280350
rect 7218 280294 7274 280350
rect 7342 280294 7398 280350
rect 6970 280170 7026 280226
rect 7094 280170 7150 280226
rect 7218 280170 7274 280226
rect 7342 280170 7398 280226
rect 6970 280046 7026 280102
rect 7094 280046 7150 280102
rect 7218 280046 7274 280102
rect 7342 280046 7398 280102
rect 6970 279922 7026 279978
rect 7094 279922 7150 279978
rect 7218 279922 7274 279978
rect 7342 279922 7398 279978
rect 6970 262294 7026 262350
rect 7094 262294 7150 262350
rect 7218 262294 7274 262350
rect 7342 262294 7398 262350
rect 6970 262170 7026 262226
rect 7094 262170 7150 262226
rect 7218 262170 7274 262226
rect 7342 262170 7398 262226
rect 6970 262046 7026 262102
rect 7094 262046 7150 262102
rect 7218 262046 7274 262102
rect 7342 262046 7398 262102
rect 6970 261922 7026 261978
rect 7094 261922 7150 261978
rect 7218 261922 7274 261978
rect 7342 261922 7398 261978
rect 6970 244294 7026 244350
rect 7094 244294 7150 244350
rect 7218 244294 7274 244350
rect 7342 244294 7398 244350
rect 6970 244170 7026 244226
rect 7094 244170 7150 244226
rect 7218 244170 7274 244226
rect 7342 244170 7398 244226
rect 6970 244046 7026 244102
rect 7094 244046 7150 244102
rect 7218 244046 7274 244102
rect 7342 244046 7398 244102
rect 6970 243922 7026 243978
rect 7094 243922 7150 243978
rect 7218 243922 7274 243978
rect 7342 243922 7398 243978
rect 6970 226294 7026 226350
rect 7094 226294 7150 226350
rect 7218 226294 7274 226350
rect 7342 226294 7398 226350
rect 6970 226170 7026 226226
rect 7094 226170 7150 226226
rect 7218 226170 7274 226226
rect 7342 226170 7398 226226
rect 6970 226046 7026 226102
rect 7094 226046 7150 226102
rect 7218 226046 7274 226102
rect 7342 226046 7398 226102
rect 6970 225922 7026 225978
rect 7094 225922 7150 225978
rect 7218 225922 7274 225978
rect 7342 225922 7398 225978
rect 6970 208294 7026 208350
rect 7094 208294 7150 208350
rect 7218 208294 7274 208350
rect 7342 208294 7398 208350
rect 6970 208170 7026 208226
rect 7094 208170 7150 208226
rect 7218 208170 7274 208226
rect 7342 208170 7398 208226
rect 6970 208046 7026 208102
rect 7094 208046 7150 208102
rect 7218 208046 7274 208102
rect 7342 208046 7398 208102
rect 6970 207922 7026 207978
rect 7094 207922 7150 207978
rect 7218 207922 7274 207978
rect 7342 207922 7398 207978
rect 6970 190294 7026 190350
rect 7094 190294 7150 190350
rect 7218 190294 7274 190350
rect 7342 190294 7398 190350
rect 6970 190170 7026 190226
rect 7094 190170 7150 190226
rect 7218 190170 7274 190226
rect 7342 190170 7398 190226
rect 6970 190046 7026 190102
rect 7094 190046 7150 190102
rect 7218 190046 7274 190102
rect 7342 190046 7398 190102
rect 6970 189922 7026 189978
rect 7094 189922 7150 189978
rect 7218 189922 7274 189978
rect 7342 189922 7398 189978
rect 6970 172294 7026 172350
rect 7094 172294 7150 172350
rect 7218 172294 7274 172350
rect 7342 172294 7398 172350
rect 6970 172170 7026 172226
rect 7094 172170 7150 172226
rect 7218 172170 7274 172226
rect 7342 172170 7398 172226
rect 6970 172046 7026 172102
rect 7094 172046 7150 172102
rect 7218 172046 7274 172102
rect 7342 172046 7398 172102
rect 6970 171922 7026 171978
rect 7094 171922 7150 171978
rect 7218 171922 7274 171978
rect 7342 171922 7398 171978
rect 6970 154294 7026 154350
rect 7094 154294 7150 154350
rect 7218 154294 7274 154350
rect 7342 154294 7398 154350
rect 6970 154170 7026 154226
rect 7094 154170 7150 154226
rect 7218 154170 7274 154226
rect 7342 154170 7398 154226
rect 6970 154046 7026 154102
rect 7094 154046 7150 154102
rect 7218 154046 7274 154102
rect 7342 154046 7398 154102
rect 6970 153922 7026 153978
rect 7094 153922 7150 153978
rect 7218 153922 7274 153978
rect 7342 153922 7398 153978
rect 6970 136294 7026 136350
rect 7094 136294 7150 136350
rect 7218 136294 7274 136350
rect 7342 136294 7398 136350
rect 6970 136170 7026 136226
rect 7094 136170 7150 136226
rect 7218 136170 7274 136226
rect 7342 136170 7398 136226
rect 6970 136046 7026 136102
rect 7094 136046 7150 136102
rect 7218 136046 7274 136102
rect 7342 136046 7398 136102
rect 6970 135922 7026 135978
rect 7094 135922 7150 135978
rect 7218 135922 7274 135978
rect 7342 135922 7398 135978
rect 6970 118294 7026 118350
rect 7094 118294 7150 118350
rect 7218 118294 7274 118350
rect 7342 118294 7398 118350
rect 6970 118170 7026 118226
rect 7094 118170 7150 118226
rect 7218 118170 7274 118226
rect 7342 118170 7398 118226
rect 6970 118046 7026 118102
rect 7094 118046 7150 118102
rect 7218 118046 7274 118102
rect 7342 118046 7398 118102
rect 6970 117922 7026 117978
rect 7094 117922 7150 117978
rect 7218 117922 7274 117978
rect 7342 117922 7398 117978
rect 6970 100294 7026 100350
rect 7094 100294 7150 100350
rect 7218 100294 7274 100350
rect 7342 100294 7398 100350
rect 6970 100170 7026 100226
rect 7094 100170 7150 100226
rect 7218 100170 7274 100226
rect 7342 100170 7398 100226
rect 6970 100046 7026 100102
rect 7094 100046 7150 100102
rect 7218 100046 7274 100102
rect 7342 100046 7398 100102
rect 6970 99922 7026 99978
rect 7094 99922 7150 99978
rect 7218 99922 7274 99978
rect 7342 99922 7398 99978
rect 6970 82294 7026 82350
rect 7094 82294 7150 82350
rect 7218 82294 7274 82350
rect 7342 82294 7398 82350
rect 6970 82170 7026 82226
rect 7094 82170 7150 82226
rect 7218 82170 7274 82226
rect 7342 82170 7398 82226
rect 6970 82046 7026 82102
rect 7094 82046 7150 82102
rect 7218 82046 7274 82102
rect 7342 82046 7398 82102
rect 6970 81922 7026 81978
rect 7094 81922 7150 81978
rect 7218 81922 7274 81978
rect 7342 81922 7398 81978
rect 6970 64294 7026 64350
rect 7094 64294 7150 64350
rect 7218 64294 7274 64350
rect 7342 64294 7398 64350
rect 6970 64170 7026 64226
rect 7094 64170 7150 64226
rect 7218 64170 7274 64226
rect 7342 64170 7398 64226
rect 6970 64046 7026 64102
rect 7094 64046 7150 64102
rect 7218 64046 7274 64102
rect 7342 64046 7398 64102
rect 6970 63922 7026 63978
rect 7094 63922 7150 63978
rect 7218 63922 7274 63978
rect 7342 63922 7398 63978
rect 6970 46294 7026 46350
rect 7094 46294 7150 46350
rect 7218 46294 7274 46350
rect 7342 46294 7398 46350
rect 6970 46170 7026 46226
rect 7094 46170 7150 46226
rect 7218 46170 7274 46226
rect 7342 46170 7398 46226
rect 6970 46046 7026 46102
rect 7094 46046 7150 46102
rect 7218 46046 7274 46102
rect 7342 46046 7398 46102
rect 6970 45922 7026 45978
rect 7094 45922 7150 45978
rect 7218 45922 7274 45978
rect 7342 45922 7398 45978
rect 6970 28294 7026 28350
rect 7094 28294 7150 28350
rect 7218 28294 7274 28350
rect 7342 28294 7398 28350
rect 6970 28170 7026 28226
rect 7094 28170 7150 28226
rect 7218 28170 7274 28226
rect 7342 28170 7398 28226
rect 6970 28046 7026 28102
rect 7094 28046 7150 28102
rect 7218 28046 7274 28102
rect 7342 28046 7398 28102
rect 6970 27922 7026 27978
rect 7094 27922 7150 27978
rect 7218 27922 7274 27978
rect 7342 27922 7398 27978
rect 6970 10294 7026 10350
rect 7094 10294 7150 10350
rect 7218 10294 7274 10350
rect 7342 10294 7398 10350
rect 6970 10170 7026 10226
rect 7094 10170 7150 10226
rect 7218 10170 7274 10226
rect 7342 10170 7398 10226
rect 6970 10046 7026 10102
rect 7094 10046 7150 10102
rect 7218 10046 7274 10102
rect 7342 10046 7398 10102
rect 6970 9922 7026 9978
rect 7094 9922 7150 9978
rect 7218 9922 7274 9978
rect 7342 9922 7398 9978
rect 6970 -1176 7026 -1120
rect 7094 -1176 7150 -1120
rect 7218 -1176 7274 -1120
rect 7342 -1176 7398 -1120
rect 6970 -1300 7026 -1244
rect 7094 -1300 7150 -1244
rect 7218 -1300 7274 -1244
rect 7342 -1300 7398 -1244
rect 6970 -1424 7026 -1368
rect 7094 -1424 7150 -1368
rect 7218 -1424 7274 -1368
rect 7342 -1424 7398 -1368
rect 6970 -1548 7026 -1492
rect 7094 -1548 7150 -1492
rect 7218 -1548 7274 -1492
rect 7342 -1548 7398 -1492
rect 21250 597156 21306 597212
rect 21374 597156 21430 597212
rect 21498 597156 21554 597212
rect 21622 597156 21678 597212
rect 21250 597032 21306 597088
rect 21374 597032 21430 597088
rect 21498 597032 21554 597088
rect 21622 597032 21678 597088
rect 21250 596908 21306 596964
rect 21374 596908 21430 596964
rect 21498 596908 21554 596964
rect 21622 596908 21678 596964
rect 21250 596784 21306 596840
rect 21374 596784 21430 596840
rect 21498 596784 21554 596840
rect 21622 596784 21678 596840
rect 21250 580294 21306 580350
rect 21374 580294 21430 580350
rect 21498 580294 21554 580350
rect 21622 580294 21678 580350
rect 21250 580170 21306 580226
rect 21374 580170 21430 580226
rect 21498 580170 21554 580226
rect 21622 580170 21678 580226
rect 21250 580046 21306 580102
rect 21374 580046 21430 580102
rect 21498 580046 21554 580102
rect 21622 580046 21678 580102
rect 21250 579922 21306 579978
rect 21374 579922 21430 579978
rect 21498 579922 21554 579978
rect 21622 579922 21678 579978
rect 21250 562294 21306 562350
rect 21374 562294 21430 562350
rect 21498 562294 21554 562350
rect 21622 562294 21678 562350
rect 21250 562170 21306 562226
rect 21374 562170 21430 562226
rect 21498 562170 21554 562226
rect 21622 562170 21678 562226
rect 21250 562046 21306 562102
rect 21374 562046 21430 562102
rect 21498 562046 21554 562102
rect 21622 562046 21678 562102
rect 21250 561922 21306 561978
rect 21374 561922 21430 561978
rect 21498 561922 21554 561978
rect 21622 561922 21678 561978
rect 21250 544294 21306 544350
rect 21374 544294 21430 544350
rect 21498 544294 21554 544350
rect 21622 544294 21678 544350
rect 21250 544170 21306 544226
rect 21374 544170 21430 544226
rect 21498 544170 21554 544226
rect 21622 544170 21678 544226
rect 21250 544046 21306 544102
rect 21374 544046 21430 544102
rect 21498 544046 21554 544102
rect 21622 544046 21678 544102
rect 21250 543922 21306 543978
rect 21374 543922 21430 543978
rect 21498 543922 21554 543978
rect 21622 543922 21678 543978
rect 21250 526294 21306 526350
rect 21374 526294 21430 526350
rect 21498 526294 21554 526350
rect 21622 526294 21678 526350
rect 21250 526170 21306 526226
rect 21374 526170 21430 526226
rect 21498 526170 21554 526226
rect 21622 526170 21678 526226
rect 21250 526046 21306 526102
rect 21374 526046 21430 526102
rect 21498 526046 21554 526102
rect 21622 526046 21678 526102
rect 21250 525922 21306 525978
rect 21374 525922 21430 525978
rect 21498 525922 21554 525978
rect 21622 525922 21678 525978
rect 21250 508294 21306 508350
rect 21374 508294 21430 508350
rect 21498 508294 21554 508350
rect 21622 508294 21678 508350
rect 21250 508170 21306 508226
rect 21374 508170 21430 508226
rect 21498 508170 21554 508226
rect 21622 508170 21678 508226
rect 21250 508046 21306 508102
rect 21374 508046 21430 508102
rect 21498 508046 21554 508102
rect 21622 508046 21678 508102
rect 21250 507922 21306 507978
rect 21374 507922 21430 507978
rect 21498 507922 21554 507978
rect 21622 507922 21678 507978
rect 21250 490294 21306 490350
rect 21374 490294 21430 490350
rect 21498 490294 21554 490350
rect 21622 490294 21678 490350
rect 21250 490170 21306 490226
rect 21374 490170 21430 490226
rect 21498 490170 21554 490226
rect 21622 490170 21678 490226
rect 21250 490046 21306 490102
rect 21374 490046 21430 490102
rect 21498 490046 21554 490102
rect 21622 490046 21678 490102
rect 21250 489922 21306 489978
rect 21374 489922 21430 489978
rect 21498 489922 21554 489978
rect 21622 489922 21678 489978
rect 21250 472294 21306 472350
rect 21374 472294 21430 472350
rect 21498 472294 21554 472350
rect 21622 472294 21678 472350
rect 21250 472170 21306 472226
rect 21374 472170 21430 472226
rect 21498 472170 21554 472226
rect 21622 472170 21678 472226
rect 21250 472046 21306 472102
rect 21374 472046 21430 472102
rect 21498 472046 21554 472102
rect 21622 472046 21678 472102
rect 21250 471922 21306 471978
rect 21374 471922 21430 471978
rect 21498 471922 21554 471978
rect 21622 471922 21678 471978
rect 21250 454294 21306 454350
rect 21374 454294 21430 454350
rect 21498 454294 21554 454350
rect 21622 454294 21678 454350
rect 21250 454170 21306 454226
rect 21374 454170 21430 454226
rect 21498 454170 21554 454226
rect 21622 454170 21678 454226
rect 21250 454046 21306 454102
rect 21374 454046 21430 454102
rect 21498 454046 21554 454102
rect 21622 454046 21678 454102
rect 21250 453922 21306 453978
rect 21374 453922 21430 453978
rect 21498 453922 21554 453978
rect 21622 453922 21678 453978
rect 21250 436294 21306 436350
rect 21374 436294 21430 436350
rect 21498 436294 21554 436350
rect 21622 436294 21678 436350
rect 21250 436170 21306 436226
rect 21374 436170 21430 436226
rect 21498 436170 21554 436226
rect 21622 436170 21678 436226
rect 21250 436046 21306 436102
rect 21374 436046 21430 436102
rect 21498 436046 21554 436102
rect 21622 436046 21678 436102
rect 21250 435922 21306 435978
rect 21374 435922 21430 435978
rect 21498 435922 21554 435978
rect 21622 435922 21678 435978
rect 21250 418294 21306 418350
rect 21374 418294 21430 418350
rect 21498 418294 21554 418350
rect 21622 418294 21678 418350
rect 21250 418170 21306 418226
rect 21374 418170 21430 418226
rect 21498 418170 21554 418226
rect 21622 418170 21678 418226
rect 21250 418046 21306 418102
rect 21374 418046 21430 418102
rect 21498 418046 21554 418102
rect 21622 418046 21678 418102
rect 21250 417922 21306 417978
rect 21374 417922 21430 417978
rect 21498 417922 21554 417978
rect 21622 417922 21678 417978
rect 21250 400294 21306 400350
rect 21374 400294 21430 400350
rect 21498 400294 21554 400350
rect 21622 400294 21678 400350
rect 21250 400170 21306 400226
rect 21374 400170 21430 400226
rect 21498 400170 21554 400226
rect 21622 400170 21678 400226
rect 21250 400046 21306 400102
rect 21374 400046 21430 400102
rect 21498 400046 21554 400102
rect 21622 400046 21678 400102
rect 21250 399922 21306 399978
rect 21374 399922 21430 399978
rect 21498 399922 21554 399978
rect 21622 399922 21678 399978
rect 21250 382294 21306 382350
rect 21374 382294 21430 382350
rect 21498 382294 21554 382350
rect 21622 382294 21678 382350
rect 21250 382170 21306 382226
rect 21374 382170 21430 382226
rect 21498 382170 21554 382226
rect 21622 382170 21678 382226
rect 21250 382046 21306 382102
rect 21374 382046 21430 382102
rect 21498 382046 21554 382102
rect 21622 382046 21678 382102
rect 21250 381922 21306 381978
rect 21374 381922 21430 381978
rect 21498 381922 21554 381978
rect 21622 381922 21678 381978
rect 21250 364294 21306 364350
rect 21374 364294 21430 364350
rect 21498 364294 21554 364350
rect 21622 364294 21678 364350
rect 21250 364170 21306 364226
rect 21374 364170 21430 364226
rect 21498 364170 21554 364226
rect 21622 364170 21678 364226
rect 21250 364046 21306 364102
rect 21374 364046 21430 364102
rect 21498 364046 21554 364102
rect 21622 364046 21678 364102
rect 21250 363922 21306 363978
rect 21374 363922 21430 363978
rect 21498 363922 21554 363978
rect 21622 363922 21678 363978
rect 21250 346294 21306 346350
rect 21374 346294 21430 346350
rect 21498 346294 21554 346350
rect 21622 346294 21678 346350
rect 21250 346170 21306 346226
rect 21374 346170 21430 346226
rect 21498 346170 21554 346226
rect 21622 346170 21678 346226
rect 21250 346046 21306 346102
rect 21374 346046 21430 346102
rect 21498 346046 21554 346102
rect 21622 346046 21678 346102
rect 21250 345922 21306 345978
rect 21374 345922 21430 345978
rect 21498 345922 21554 345978
rect 21622 345922 21678 345978
rect 21250 328294 21306 328350
rect 21374 328294 21430 328350
rect 21498 328294 21554 328350
rect 21622 328294 21678 328350
rect 21250 328170 21306 328226
rect 21374 328170 21430 328226
rect 21498 328170 21554 328226
rect 21622 328170 21678 328226
rect 21250 328046 21306 328102
rect 21374 328046 21430 328102
rect 21498 328046 21554 328102
rect 21622 328046 21678 328102
rect 21250 327922 21306 327978
rect 21374 327922 21430 327978
rect 21498 327922 21554 327978
rect 21622 327922 21678 327978
rect 21250 310294 21306 310350
rect 21374 310294 21430 310350
rect 21498 310294 21554 310350
rect 21622 310294 21678 310350
rect 21250 310170 21306 310226
rect 21374 310170 21430 310226
rect 21498 310170 21554 310226
rect 21622 310170 21678 310226
rect 21250 310046 21306 310102
rect 21374 310046 21430 310102
rect 21498 310046 21554 310102
rect 21622 310046 21678 310102
rect 21250 309922 21306 309978
rect 21374 309922 21430 309978
rect 21498 309922 21554 309978
rect 21622 309922 21678 309978
rect 21250 292294 21306 292350
rect 21374 292294 21430 292350
rect 21498 292294 21554 292350
rect 21622 292294 21678 292350
rect 21250 292170 21306 292226
rect 21374 292170 21430 292226
rect 21498 292170 21554 292226
rect 21622 292170 21678 292226
rect 21250 292046 21306 292102
rect 21374 292046 21430 292102
rect 21498 292046 21554 292102
rect 21622 292046 21678 292102
rect 21250 291922 21306 291978
rect 21374 291922 21430 291978
rect 21498 291922 21554 291978
rect 21622 291922 21678 291978
rect 21250 274294 21306 274350
rect 21374 274294 21430 274350
rect 21498 274294 21554 274350
rect 21622 274294 21678 274350
rect 21250 274170 21306 274226
rect 21374 274170 21430 274226
rect 21498 274170 21554 274226
rect 21622 274170 21678 274226
rect 21250 274046 21306 274102
rect 21374 274046 21430 274102
rect 21498 274046 21554 274102
rect 21622 274046 21678 274102
rect 21250 273922 21306 273978
rect 21374 273922 21430 273978
rect 21498 273922 21554 273978
rect 21622 273922 21678 273978
rect 21250 256294 21306 256350
rect 21374 256294 21430 256350
rect 21498 256294 21554 256350
rect 21622 256294 21678 256350
rect 21250 256170 21306 256226
rect 21374 256170 21430 256226
rect 21498 256170 21554 256226
rect 21622 256170 21678 256226
rect 21250 256046 21306 256102
rect 21374 256046 21430 256102
rect 21498 256046 21554 256102
rect 21622 256046 21678 256102
rect 21250 255922 21306 255978
rect 21374 255922 21430 255978
rect 21498 255922 21554 255978
rect 21622 255922 21678 255978
rect 21250 238294 21306 238350
rect 21374 238294 21430 238350
rect 21498 238294 21554 238350
rect 21622 238294 21678 238350
rect 21250 238170 21306 238226
rect 21374 238170 21430 238226
rect 21498 238170 21554 238226
rect 21622 238170 21678 238226
rect 21250 238046 21306 238102
rect 21374 238046 21430 238102
rect 21498 238046 21554 238102
rect 21622 238046 21678 238102
rect 21250 237922 21306 237978
rect 21374 237922 21430 237978
rect 21498 237922 21554 237978
rect 21622 237922 21678 237978
rect 21250 220294 21306 220350
rect 21374 220294 21430 220350
rect 21498 220294 21554 220350
rect 21622 220294 21678 220350
rect 21250 220170 21306 220226
rect 21374 220170 21430 220226
rect 21498 220170 21554 220226
rect 21622 220170 21678 220226
rect 21250 220046 21306 220102
rect 21374 220046 21430 220102
rect 21498 220046 21554 220102
rect 21622 220046 21678 220102
rect 21250 219922 21306 219978
rect 21374 219922 21430 219978
rect 21498 219922 21554 219978
rect 21622 219922 21678 219978
rect 21250 202294 21306 202350
rect 21374 202294 21430 202350
rect 21498 202294 21554 202350
rect 21622 202294 21678 202350
rect 21250 202170 21306 202226
rect 21374 202170 21430 202226
rect 21498 202170 21554 202226
rect 21622 202170 21678 202226
rect 21250 202046 21306 202102
rect 21374 202046 21430 202102
rect 21498 202046 21554 202102
rect 21622 202046 21678 202102
rect 21250 201922 21306 201978
rect 21374 201922 21430 201978
rect 21498 201922 21554 201978
rect 21622 201922 21678 201978
rect 21250 184294 21306 184350
rect 21374 184294 21430 184350
rect 21498 184294 21554 184350
rect 21622 184294 21678 184350
rect 21250 184170 21306 184226
rect 21374 184170 21430 184226
rect 21498 184170 21554 184226
rect 21622 184170 21678 184226
rect 21250 184046 21306 184102
rect 21374 184046 21430 184102
rect 21498 184046 21554 184102
rect 21622 184046 21678 184102
rect 21250 183922 21306 183978
rect 21374 183922 21430 183978
rect 21498 183922 21554 183978
rect 21622 183922 21678 183978
rect 21250 166294 21306 166350
rect 21374 166294 21430 166350
rect 21498 166294 21554 166350
rect 21622 166294 21678 166350
rect 21250 166170 21306 166226
rect 21374 166170 21430 166226
rect 21498 166170 21554 166226
rect 21622 166170 21678 166226
rect 21250 166046 21306 166102
rect 21374 166046 21430 166102
rect 21498 166046 21554 166102
rect 21622 166046 21678 166102
rect 21250 165922 21306 165978
rect 21374 165922 21430 165978
rect 21498 165922 21554 165978
rect 21622 165922 21678 165978
rect 21250 148294 21306 148350
rect 21374 148294 21430 148350
rect 21498 148294 21554 148350
rect 21622 148294 21678 148350
rect 21250 148170 21306 148226
rect 21374 148170 21430 148226
rect 21498 148170 21554 148226
rect 21622 148170 21678 148226
rect 21250 148046 21306 148102
rect 21374 148046 21430 148102
rect 21498 148046 21554 148102
rect 21622 148046 21678 148102
rect 21250 147922 21306 147978
rect 21374 147922 21430 147978
rect 21498 147922 21554 147978
rect 21622 147922 21678 147978
rect 21250 130294 21306 130350
rect 21374 130294 21430 130350
rect 21498 130294 21554 130350
rect 21622 130294 21678 130350
rect 21250 130170 21306 130226
rect 21374 130170 21430 130226
rect 21498 130170 21554 130226
rect 21622 130170 21678 130226
rect 21250 130046 21306 130102
rect 21374 130046 21430 130102
rect 21498 130046 21554 130102
rect 21622 130046 21678 130102
rect 21250 129922 21306 129978
rect 21374 129922 21430 129978
rect 21498 129922 21554 129978
rect 21622 129922 21678 129978
rect 21250 112294 21306 112350
rect 21374 112294 21430 112350
rect 21498 112294 21554 112350
rect 21622 112294 21678 112350
rect 21250 112170 21306 112226
rect 21374 112170 21430 112226
rect 21498 112170 21554 112226
rect 21622 112170 21678 112226
rect 21250 112046 21306 112102
rect 21374 112046 21430 112102
rect 21498 112046 21554 112102
rect 21622 112046 21678 112102
rect 21250 111922 21306 111978
rect 21374 111922 21430 111978
rect 21498 111922 21554 111978
rect 21622 111922 21678 111978
rect 21250 94294 21306 94350
rect 21374 94294 21430 94350
rect 21498 94294 21554 94350
rect 21622 94294 21678 94350
rect 21250 94170 21306 94226
rect 21374 94170 21430 94226
rect 21498 94170 21554 94226
rect 21622 94170 21678 94226
rect 21250 94046 21306 94102
rect 21374 94046 21430 94102
rect 21498 94046 21554 94102
rect 21622 94046 21678 94102
rect 21250 93922 21306 93978
rect 21374 93922 21430 93978
rect 21498 93922 21554 93978
rect 21622 93922 21678 93978
rect 21250 76294 21306 76350
rect 21374 76294 21430 76350
rect 21498 76294 21554 76350
rect 21622 76294 21678 76350
rect 21250 76170 21306 76226
rect 21374 76170 21430 76226
rect 21498 76170 21554 76226
rect 21622 76170 21678 76226
rect 21250 76046 21306 76102
rect 21374 76046 21430 76102
rect 21498 76046 21554 76102
rect 21622 76046 21678 76102
rect 21250 75922 21306 75978
rect 21374 75922 21430 75978
rect 21498 75922 21554 75978
rect 21622 75922 21678 75978
rect 21250 58294 21306 58350
rect 21374 58294 21430 58350
rect 21498 58294 21554 58350
rect 21622 58294 21678 58350
rect 21250 58170 21306 58226
rect 21374 58170 21430 58226
rect 21498 58170 21554 58226
rect 21622 58170 21678 58226
rect 21250 58046 21306 58102
rect 21374 58046 21430 58102
rect 21498 58046 21554 58102
rect 21622 58046 21678 58102
rect 21250 57922 21306 57978
rect 21374 57922 21430 57978
rect 21498 57922 21554 57978
rect 21622 57922 21678 57978
rect 21250 40294 21306 40350
rect 21374 40294 21430 40350
rect 21498 40294 21554 40350
rect 21622 40294 21678 40350
rect 21250 40170 21306 40226
rect 21374 40170 21430 40226
rect 21498 40170 21554 40226
rect 21622 40170 21678 40226
rect 21250 40046 21306 40102
rect 21374 40046 21430 40102
rect 21498 40046 21554 40102
rect 21622 40046 21678 40102
rect 21250 39922 21306 39978
rect 21374 39922 21430 39978
rect 21498 39922 21554 39978
rect 21622 39922 21678 39978
rect 21250 22294 21306 22350
rect 21374 22294 21430 22350
rect 21498 22294 21554 22350
rect 21622 22294 21678 22350
rect 21250 22170 21306 22226
rect 21374 22170 21430 22226
rect 21498 22170 21554 22226
rect 21622 22170 21678 22226
rect 21250 22046 21306 22102
rect 21374 22046 21430 22102
rect 21498 22046 21554 22102
rect 21622 22046 21678 22102
rect 21250 21922 21306 21978
rect 21374 21922 21430 21978
rect 21498 21922 21554 21978
rect 21622 21922 21678 21978
rect 21250 4294 21306 4350
rect 21374 4294 21430 4350
rect 21498 4294 21554 4350
rect 21622 4294 21678 4350
rect 21250 4170 21306 4226
rect 21374 4170 21430 4226
rect 21498 4170 21554 4226
rect 21622 4170 21678 4226
rect 21250 4046 21306 4102
rect 21374 4046 21430 4102
rect 21498 4046 21554 4102
rect 21622 4046 21678 4102
rect 21250 3922 21306 3978
rect 21374 3922 21430 3978
rect 21498 3922 21554 3978
rect 21622 3922 21678 3978
rect 21250 -216 21306 -160
rect 21374 -216 21430 -160
rect 21498 -216 21554 -160
rect 21622 -216 21678 -160
rect 21250 -340 21306 -284
rect 21374 -340 21430 -284
rect 21498 -340 21554 -284
rect 21622 -340 21678 -284
rect 21250 -464 21306 -408
rect 21374 -464 21430 -408
rect 21498 -464 21554 -408
rect 21622 -464 21678 -408
rect 21250 -588 21306 -532
rect 21374 -588 21430 -532
rect 21498 -588 21554 -532
rect 21622 -588 21678 -532
rect 24970 598116 25026 598172
rect 25094 598116 25150 598172
rect 25218 598116 25274 598172
rect 25342 598116 25398 598172
rect 24970 597992 25026 598048
rect 25094 597992 25150 598048
rect 25218 597992 25274 598048
rect 25342 597992 25398 598048
rect 24970 597868 25026 597924
rect 25094 597868 25150 597924
rect 25218 597868 25274 597924
rect 25342 597868 25398 597924
rect 24970 597744 25026 597800
rect 25094 597744 25150 597800
rect 25218 597744 25274 597800
rect 25342 597744 25398 597800
rect 24970 586294 25026 586350
rect 25094 586294 25150 586350
rect 25218 586294 25274 586350
rect 25342 586294 25398 586350
rect 24970 586170 25026 586226
rect 25094 586170 25150 586226
rect 25218 586170 25274 586226
rect 25342 586170 25398 586226
rect 24970 586046 25026 586102
rect 25094 586046 25150 586102
rect 25218 586046 25274 586102
rect 25342 586046 25398 586102
rect 24970 585922 25026 585978
rect 25094 585922 25150 585978
rect 25218 585922 25274 585978
rect 25342 585922 25398 585978
rect 24970 568294 25026 568350
rect 25094 568294 25150 568350
rect 25218 568294 25274 568350
rect 25342 568294 25398 568350
rect 24970 568170 25026 568226
rect 25094 568170 25150 568226
rect 25218 568170 25274 568226
rect 25342 568170 25398 568226
rect 24970 568046 25026 568102
rect 25094 568046 25150 568102
rect 25218 568046 25274 568102
rect 25342 568046 25398 568102
rect 24970 567922 25026 567978
rect 25094 567922 25150 567978
rect 25218 567922 25274 567978
rect 25342 567922 25398 567978
rect 24970 550294 25026 550350
rect 25094 550294 25150 550350
rect 25218 550294 25274 550350
rect 25342 550294 25398 550350
rect 24970 550170 25026 550226
rect 25094 550170 25150 550226
rect 25218 550170 25274 550226
rect 25342 550170 25398 550226
rect 24970 550046 25026 550102
rect 25094 550046 25150 550102
rect 25218 550046 25274 550102
rect 25342 550046 25398 550102
rect 24970 549922 25026 549978
rect 25094 549922 25150 549978
rect 25218 549922 25274 549978
rect 25342 549922 25398 549978
rect 24970 532294 25026 532350
rect 25094 532294 25150 532350
rect 25218 532294 25274 532350
rect 25342 532294 25398 532350
rect 24970 532170 25026 532226
rect 25094 532170 25150 532226
rect 25218 532170 25274 532226
rect 25342 532170 25398 532226
rect 24970 532046 25026 532102
rect 25094 532046 25150 532102
rect 25218 532046 25274 532102
rect 25342 532046 25398 532102
rect 24970 531922 25026 531978
rect 25094 531922 25150 531978
rect 25218 531922 25274 531978
rect 25342 531922 25398 531978
rect 24970 514294 25026 514350
rect 25094 514294 25150 514350
rect 25218 514294 25274 514350
rect 25342 514294 25398 514350
rect 24970 514170 25026 514226
rect 25094 514170 25150 514226
rect 25218 514170 25274 514226
rect 25342 514170 25398 514226
rect 24970 514046 25026 514102
rect 25094 514046 25150 514102
rect 25218 514046 25274 514102
rect 25342 514046 25398 514102
rect 24970 513922 25026 513978
rect 25094 513922 25150 513978
rect 25218 513922 25274 513978
rect 25342 513922 25398 513978
rect 24970 496294 25026 496350
rect 25094 496294 25150 496350
rect 25218 496294 25274 496350
rect 25342 496294 25398 496350
rect 24970 496170 25026 496226
rect 25094 496170 25150 496226
rect 25218 496170 25274 496226
rect 25342 496170 25398 496226
rect 24970 496046 25026 496102
rect 25094 496046 25150 496102
rect 25218 496046 25274 496102
rect 25342 496046 25398 496102
rect 24970 495922 25026 495978
rect 25094 495922 25150 495978
rect 25218 495922 25274 495978
rect 25342 495922 25398 495978
rect 24970 478294 25026 478350
rect 25094 478294 25150 478350
rect 25218 478294 25274 478350
rect 25342 478294 25398 478350
rect 24970 478170 25026 478226
rect 25094 478170 25150 478226
rect 25218 478170 25274 478226
rect 25342 478170 25398 478226
rect 24970 478046 25026 478102
rect 25094 478046 25150 478102
rect 25218 478046 25274 478102
rect 25342 478046 25398 478102
rect 24970 477922 25026 477978
rect 25094 477922 25150 477978
rect 25218 477922 25274 477978
rect 25342 477922 25398 477978
rect 24970 460294 25026 460350
rect 25094 460294 25150 460350
rect 25218 460294 25274 460350
rect 25342 460294 25398 460350
rect 24970 460170 25026 460226
rect 25094 460170 25150 460226
rect 25218 460170 25274 460226
rect 25342 460170 25398 460226
rect 24970 460046 25026 460102
rect 25094 460046 25150 460102
rect 25218 460046 25274 460102
rect 25342 460046 25398 460102
rect 24970 459922 25026 459978
rect 25094 459922 25150 459978
rect 25218 459922 25274 459978
rect 25342 459922 25398 459978
rect 24970 442294 25026 442350
rect 25094 442294 25150 442350
rect 25218 442294 25274 442350
rect 25342 442294 25398 442350
rect 24970 442170 25026 442226
rect 25094 442170 25150 442226
rect 25218 442170 25274 442226
rect 25342 442170 25398 442226
rect 24970 442046 25026 442102
rect 25094 442046 25150 442102
rect 25218 442046 25274 442102
rect 25342 442046 25398 442102
rect 24970 441922 25026 441978
rect 25094 441922 25150 441978
rect 25218 441922 25274 441978
rect 25342 441922 25398 441978
rect 24970 424294 25026 424350
rect 25094 424294 25150 424350
rect 25218 424294 25274 424350
rect 25342 424294 25398 424350
rect 24970 424170 25026 424226
rect 25094 424170 25150 424226
rect 25218 424170 25274 424226
rect 25342 424170 25398 424226
rect 24970 424046 25026 424102
rect 25094 424046 25150 424102
rect 25218 424046 25274 424102
rect 25342 424046 25398 424102
rect 24970 423922 25026 423978
rect 25094 423922 25150 423978
rect 25218 423922 25274 423978
rect 25342 423922 25398 423978
rect 24970 406294 25026 406350
rect 25094 406294 25150 406350
rect 25218 406294 25274 406350
rect 25342 406294 25398 406350
rect 24970 406170 25026 406226
rect 25094 406170 25150 406226
rect 25218 406170 25274 406226
rect 25342 406170 25398 406226
rect 24970 406046 25026 406102
rect 25094 406046 25150 406102
rect 25218 406046 25274 406102
rect 25342 406046 25398 406102
rect 24970 405922 25026 405978
rect 25094 405922 25150 405978
rect 25218 405922 25274 405978
rect 25342 405922 25398 405978
rect 24970 388294 25026 388350
rect 25094 388294 25150 388350
rect 25218 388294 25274 388350
rect 25342 388294 25398 388350
rect 24970 388170 25026 388226
rect 25094 388170 25150 388226
rect 25218 388170 25274 388226
rect 25342 388170 25398 388226
rect 24970 388046 25026 388102
rect 25094 388046 25150 388102
rect 25218 388046 25274 388102
rect 25342 388046 25398 388102
rect 24970 387922 25026 387978
rect 25094 387922 25150 387978
rect 25218 387922 25274 387978
rect 25342 387922 25398 387978
rect 24970 370294 25026 370350
rect 25094 370294 25150 370350
rect 25218 370294 25274 370350
rect 25342 370294 25398 370350
rect 24970 370170 25026 370226
rect 25094 370170 25150 370226
rect 25218 370170 25274 370226
rect 25342 370170 25398 370226
rect 24970 370046 25026 370102
rect 25094 370046 25150 370102
rect 25218 370046 25274 370102
rect 25342 370046 25398 370102
rect 24970 369922 25026 369978
rect 25094 369922 25150 369978
rect 25218 369922 25274 369978
rect 25342 369922 25398 369978
rect 24970 352294 25026 352350
rect 25094 352294 25150 352350
rect 25218 352294 25274 352350
rect 25342 352294 25398 352350
rect 24970 352170 25026 352226
rect 25094 352170 25150 352226
rect 25218 352170 25274 352226
rect 25342 352170 25398 352226
rect 24970 352046 25026 352102
rect 25094 352046 25150 352102
rect 25218 352046 25274 352102
rect 25342 352046 25398 352102
rect 24970 351922 25026 351978
rect 25094 351922 25150 351978
rect 25218 351922 25274 351978
rect 25342 351922 25398 351978
rect 24970 334294 25026 334350
rect 25094 334294 25150 334350
rect 25218 334294 25274 334350
rect 25342 334294 25398 334350
rect 24970 334170 25026 334226
rect 25094 334170 25150 334226
rect 25218 334170 25274 334226
rect 25342 334170 25398 334226
rect 24970 334046 25026 334102
rect 25094 334046 25150 334102
rect 25218 334046 25274 334102
rect 25342 334046 25398 334102
rect 24970 333922 25026 333978
rect 25094 333922 25150 333978
rect 25218 333922 25274 333978
rect 25342 333922 25398 333978
rect 24970 316294 25026 316350
rect 25094 316294 25150 316350
rect 25218 316294 25274 316350
rect 25342 316294 25398 316350
rect 24970 316170 25026 316226
rect 25094 316170 25150 316226
rect 25218 316170 25274 316226
rect 25342 316170 25398 316226
rect 24970 316046 25026 316102
rect 25094 316046 25150 316102
rect 25218 316046 25274 316102
rect 25342 316046 25398 316102
rect 24970 315922 25026 315978
rect 25094 315922 25150 315978
rect 25218 315922 25274 315978
rect 25342 315922 25398 315978
rect 24970 298294 25026 298350
rect 25094 298294 25150 298350
rect 25218 298294 25274 298350
rect 25342 298294 25398 298350
rect 24970 298170 25026 298226
rect 25094 298170 25150 298226
rect 25218 298170 25274 298226
rect 25342 298170 25398 298226
rect 24970 298046 25026 298102
rect 25094 298046 25150 298102
rect 25218 298046 25274 298102
rect 25342 298046 25398 298102
rect 24970 297922 25026 297978
rect 25094 297922 25150 297978
rect 25218 297922 25274 297978
rect 25342 297922 25398 297978
rect 24970 280294 25026 280350
rect 25094 280294 25150 280350
rect 25218 280294 25274 280350
rect 25342 280294 25398 280350
rect 24970 280170 25026 280226
rect 25094 280170 25150 280226
rect 25218 280170 25274 280226
rect 25342 280170 25398 280226
rect 24970 280046 25026 280102
rect 25094 280046 25150 280102
rect 25218 280046 25274 280102
rect 25342 280046 25398 280102
rect 24970 279922 25026 279978
rect 25094 279922 25150 279978
rect 25218 279922 25274 279978
rect 25342 279922 25398 279978
rect 24970 262294 25026 262350
rect 25094 262294 25150 262350
rect 25218 262294 25274 262350
rect 25342 262294 25398 262350
rect 24970 262170 25026 262226
rect 25094 262170 25150 262226
rect 25218 262170 25274 262226
rect 25342 262170 25398 262226
rect 24970 262046 25026 262102
rect 25094 262046 25150 262102
rect 25218 262046 25274 262102
rect 25342 262046 25398 262102
rect 24970 261922 25026 261978
rect 25094 261922 25150 261978
rect 25218 261922 25274 261978
rect 25342 261922 25398 261978
rect 24970 244294 25026 244350
rect 25094 244294 25150 244350
rect 25218 244294 25274 244350
rect 25342 244294 25398 244350
rect 24970 244170 25026 244226
rect 25094 244170 25150 244226
rect 25218 244170 25274 244226
rect 25342 244170 25398 244226
rect 24970 244046 25026 244102
rect 25094 244046 25150 244102
rect 25218 244046 25274 244102
rect 25342 244046 25398 244102
rect 24970 243922 25026 243978
rect 25094 243922 25150 243978
rect 25218 243922 25274 243978
rect 25342 243922 25398 243978
rect 24970 226294 25026 226350
rect 25094 226294 25150 226350
rect 25218 226294 25274 226350
rect 25342 226294 25398 226350
rect 24970 226170 25026 226226
rect 25094 226170 25150 226226
rect 25218 226170 25274 226226
rect 25342 226170 25398 226226
rect 24970 226046 25026 226102
rect 25094 226046 25150 226102
rect 25218 226046 25274 226102
rect 25342 226046 25398 226102
rect 24970 225922 25026 225978
rect 25094 225922 25150 225978
rect 25218 225922 25274 225978
rect 25342 225922 25398 225978
rect 24970 208294 25026 208350
rect 25094 208294 25150 208350
rect 25218 208294 25274 208350
rect 25342 208294 25398 208350
rect 24970 208170 25026 208226
rect 25094 208170 25150 208226
rect 25218 208170 25274 208226
rect 25342 208170 25398 208226
rect 24970 208046 25026 208102
rect 25094 208046 25150 208102
rect 25218 208046 25274 208102
rect 25342 208046 25398 208102
rect 24970 207922 25026 207978
rect 25094 207922 25150 207978
rect 25218 207922 25274 207978
rect 25342 207922 25398 207978
rect 24970 190294 25026 190350
rect 25094 190294 25150 190350
rect 25218 190294 25274 190350
rect 25342 190294 25398 190350
rect 24970 190170 25026 190226
rect 25094 190170 25150 190226
rect 25218 190170 25274 190226
rect 25342 190170 25398 190226
rect 24970 190046 25026 190102
rect 25094 190046 25150 190102
rect 25218 190046 25274 190102
rect 25342 190046 25398 190102
rect 24970 189922 25026 189978
rect 25094 189922 25150 189978
rect 25218 189922 25274 189978
rect 25342 189922 25398 189978
rect 24970 172294 25026 172350
rect 25094 172294 25150 172350
rect 25218 172294 25274 172350
rect 25342 172294 25398 172350
rect 24970 172170 25026 172226
rect 25094 172170 25150 172226
rect 25218 172170 25274 172226
rect 25342 172170 25398 172226
rect 24970 172046 25026 172102
rect 25094 172046 25150 172102
rect 25218 172046 25274 172102
rect 25342 172046 25398 172102
rect 24970 171922 25026 171978
rect 25094 171922 25150 171978
rect 25218 171922 25274 171978
rect 25342 171922 25398 171978
rect 24970 154294 25026 154350
rect 25094 154294 25150 154350
rect 25218 154294 25274 154350
rect 25342 154294 25398 154350
rect 24970 154170 25026 154226
rect 25094 154170 25150 154226
rect 25218 154170 25274 154226
rect 25342 154170 25398 154226
rect 24970 154046 25026 154102
rect 25094 154046 25150 154102
rect 25218 154046 25274 154102
rect 25342 154046 25398 154102
rect 24970 153922 25026 153978
rect 25094 153922 25150 153978
rect 25218 153922 25274 153978
rect 25342 153922 25398 153978
rect 24970 136294 25026 136350
rect 25094 136294 25150 136350
rect 25218 136294 25274 136350
rect 25342 136294 25398 136350
rect 24970 136170 25026 136226
rect 25094 136170 25150 136226
rect 25218 136170 25274 136226
rect 25342 136170 25398 136226
rect 24970 136046 25026 136102
rect 25094 136046 25150 136102
rect 25218 136046 25274 136102
rect 25342 136046 25398 136102
rect 24970 135922 25026 135978
rect 25094 135922 25150 135978
rect 25218 135922 25274 135978
rect 25342 135922 25398 135978
rect 24970 118294 25026 118350
rect 25094 118294 25150 118350
rect 25218 118294 25274 118350
rect 25342 118294 25398 118350
rect 24970 118170 25026 118226
rect 25094 118170 25150 118226
rect 25218 118170 25274 118226
rect 25342 118170 25398 118226
rect 24970 118046 25026 118102
rect 25094 118046 25150 118102
rect 25218 118046 25274 118102
rect 25342 118046 25398 118102
rect 24970 117922 25026 117978
rect 25094 117922 25150 117978
rect 25218 117922 25274 117978
rect 25342 117922 25398 117978
rect 24970 100294 25026 100350
rect 25094 100294 25150 100350
rect 25218 100294 25274 100350
rect 25342 100294 25398 100350
rect 24970 100170 25026 100226
rect 25094 100170 25150 100226
rect 25218 100170 25274 100226
rect 25342 100170 25398 100226
rect 24970 100046 25026 100102
rect 25094 100046 25150 100102
rect 25218 100046 25274 100102
rect 25342 100046 25398 100102
rect 24970 99922 25026 99978
rect 25094 99922 25150 99978
rect 25218 99922 25274 99978
rect 25342 99922 25398 99978
rect 24970 82294 25026 82350
rect 25094 82294 25150 82350
rect 25218 82294 25274 82350
rect 25342 82294 25398 82350
rect 24970 82170 25026 82226
rect 25094 82170 25150 82226
rect 25218 82170 25274 82226
rect 25342 82170 25398 82226
rect 24970 82046 25026 82102
rect 25094 82046 25150 82102
rect 25218 82046 25274 82102
rect 25342 82046 25398 82102
rect 24970 81922 25026 81978
rect 25094 81922 25150 81978
rect 25218 81922 25274 81978
rect 25342 81922 25398 81978
rect 24970 64294 25026 64350
rect 25094 64294 25150 64350
rect 25218 64294 25274 64350
rect 25342 64294 25398 64350
rect 24970 64170 25026 64226
rect 25094 64170 25150 64226
rect 25218 64170 25274 64226
rect 25342 64170 25398 64226
rect 24970 64046 25026 64102
rect 25094 64046 25150 64102
rect 25218 64046 25274 64102
rect 25342 64046 25398 64102
rect 24970 63922 25026 63978
rect 25094 63922 25150 63978
rect 25218 63922 25274 63978
rect 25342 63922 25398 63978
rect 24970 46294 25026 46350
rect 25094 46294 25150 46350
rect 25218 46294 25274 46350
rect 25342 46294 25398 46350
rect 24970 46170 25026 46226
rect 25094 46170 25150 46226
rect 25218 46170 25274 46226
rect 25342 46170 25398 46226
rect 24970 46046 25026 46102
rect 25094 46046 25150 46102
rect 25218 46046 25274 46102
rect 25342 46046 25398 46102
rect 24970 45922 25026 45978
rect 25094 45922 25150 45978
rect 25218 45922 25274 45978
rect 25342 45922 25398 45978
rect 24970 28294 25026 28350
rect 25094 28294 25150 28350
rect 25218 28294 25274 28350
rect 25342 28294 25398 28350
rect 24970 28170 25026 28226
rect 25094 28170 25150 28226
rect 25218 28170 25274 28226
rect 25342 28170 25398 28226
rect 24970 28046 25026 28102
rect 25094 28046 25150 28102
rect 25218 28046 25274 28102
rect 25342 28046 25398 28102
rect 24970 27922 25026 27978
rect 25094 27922 25150 27978
rect 25218 27922 25274 27978
rect 25342 27922 25398 27978
rect 24970 10294 25026 10350
rect 25094 10294 25150 10350
rect 25218 10294 25274 10350
rect 25342 10294 25398 10350
rect 24970 10170 25026 10226
rect 25094 10170 25150 10226
rect 25218 10170 25274 10226
rect 25342 10170 25398 10226
rect 24970 10046 25026 10102
rect 25094 10046 25150 10102
rect 25218 10046 25274 10102
rect 25342 10046 25398 10102
rect 24970 9922 25026 9978
rect 25094 9922 25150 9978
rect 25218 9922 25274 9978
rect 25342 9922 25398 9978
rect 24970 -1176 25026 -1120
rect 25094 -1176 25150 -1120
rect 25218 -1176 25274 -1120
rect 25342 -1176 25398 -1120
rect 24970 -1300 25026 -1244
rect 25094 -1300 25150 -1244
rect 25218 -1300 25274 -1244
rect 25342 -1300 25398 -1244
rect 24970 -1424 25026 -1368
rect 25094 -1424 25150 -1368
rect 25218 -1424 25274 -1368
rect 25342 -1424 25398 -1368
rect 24970 -1548 25026 -1492
rect 25094 -1548 25150 -1492
rect 25218 -1548 25274 -1492
rect 25342 -1548 25398 -1492
rect 39250 597156 39306 597212
rect 39374 597156 39430 597212
rect 39498 597156 39554 597212
rect 39622 597156 39678 597212
rect 39250 597032 39306 597088
rect 39374 597032 39430 597088
rect 39498 597032 39554 597088
rect 39622 597032 39678 597088
rect 39250 596908 39306 596964
rect 39374 596908 39430 596964
rect 39498 596908 39554 596964
rect 39622 596908 39678 596964
rect 39250 596784 39306 596840
rect 39374 596784 39430 596840
rect 39498 596784 39554 596840
rect 39622 596784 39678 596840
rect 39250 580294 39306 580350
rect 39374 580294 39430 580350
rect 39498 580294 39554 580350
rect 39622 580294 39678 580350
rect 39250 580170 39306 580226
rect 39374 580170 39430 580226
rect 39498 580170 39554 580226
rect 39622 580170 39678 580226
rect 39250 580046 39306 580102
rect 39374 580046 39430 580102
rect 39498 580046 39554 580102
rect 39622 580046 39678 580102
rect 39250 579922 39306 579978
rect 39374 579922 39430 579978
rect 39498 579922 39554 579978
rect 39622 579922 39678 579978
rect 39250 562294 39306 562350
rect 39374 562294 39430 562350
rect 39498 562294 39554 562350
rect 39622 562294 39678 562350
rect 39250 562170 39306 562226
rect 39374 562170 39430 562226
rect 39498 562170 39554 562226
rect 39622 562170 39678 562226
rect 39250 562046 39306 562102
rect 39374 562046 39430 562102
rect 39498 562046 39554 562102
rect 39622 562046 39678 562102
rect 39250 561922 39306 561978
rect 39374 561922 39430 561978
rect 39498 561922 39554 561978
rect 39622 561922 39678 561978
rect 39250 544294 39306 544350
rect 39374 544294 39430 544350
rect 39498 544294 39554 544350
rect 39622 544294 39678 544350
rect 39250 544170 39306 544226
rect 39374 544170 39430 544226
rect 39498 544170 39554 544226
rect 39622 544170 39678 544226
rect 39250 544046 39306 544102
rect 39374 544046 39430 544102
rect 39498 544046 39554 544102
rect 39622 544046 39678 544102
rect 39250 543922 39306 543978
rect 39374 543922 39430 543978
rect 39498 543922 39554 543978
rect 39622 543922 39678 543978
rect 39250 526294 39306 526350
rect 39374 526294 39430 526350
rect 39498 526294 39554 526350
rect 39622 526294 39678 526350
rect 39250 526170 39306 526226
rect 39374 526170 39430 526226
rect 39498 526170 39554 526226
rect 39622 526170 39678 526226
rect 39250 526046 39306 526102
rect 39374 526046 39430 526102
rect 39498 526046 39554 526102
rect 39622 526046 39678 526102
rect 39250 525922 39306 525978
rect 39374 525922 39430 525978
rect 39498 525922 39554 525978
rect 39622 525922 39678 525978
rect 39250 508294 39306 508350
rect 39374 508294 39430 508350
rect 39498 508294 39554 508350
rect 39622 508294 39678 508350
rect 39250 508170 39306 508226
rect 39374 508170 39430 508226
rect 39498 508170 39554 508226
rect 39622 508170 39678 508226
rect 39250 508046 39306 508102
rect 39374 508046 39430 508102
rect 39498 508046 39554 508102
rect 39622 508046 39678 508102
rect 39250 507922 39306 507978
rect 39374 507922 39430 507978
rect 39498 507922 39554 507978
rect 39622 507922 39678 507978
rect 39250 490294 39306 490350
rect 39374 490294 39430 490350
rect 39498 490294 39554 490350
rect 39622 490294 39678 490350
rect 39250 490170 39306 490226
rect 39374 490170 39430 490226
rect 39498 490170 39554 490226
rect 39622 490170 39678 490226
rect 39250 490046 39306 490102
rect 39374 490046 39430 490102
rect 39498 490046 39554 490102
rect 39622 490046 39678 490102
rect 39250 489922 39306 489978
rect 39374 489922 39430 489978
rect 39498 489922 39554 489978
rect 39622 489922 39678 489978
rect 39250 472294 39306 472350
rect 39374 472294 39430 472350
rect 39498 472294 39554 472350
rect 39622 472294 39678 472350
rect 39250 472170 39306 472226
rect 39374 472170 39430 472226
rect 39498 472170 39554 472226
rect 39622 472170 39678 472226
rect 39250 472046 39306 472102
rect 39374 472046 39430 472102
rect 39498 472046 39554 472102
rect 39622 472046 39678 472102
rect 39250 471922 39306 471978
rect 39374 471922 39430 471978
rect 39498 471922 39554 471978
rect 39622 471922 39678 471978
rect 39250 454294 39306 454350
rect 39374 454294 39430 454350
rect 39498 454294 39554 454350
rect 39622 454294 39678 454350
rect 39250 454170 39306 454226
rect 39374 454170 39430 454226
rect 39498 454170 39554 454226
rect 39622 454170 39678 454226
rect 39250 454046 39306 454102
rect 39374 454046 39430 454102
rect 39498 454046 39554 454102
rect 39622 454046 39678 454102
rect 39250 453922 39306 453978
rect 39374 453922 39430 453978
rect 39498 453922 39554 453978
rect 39622 453922 39678 453978
rect 39250 436294 39306 436350
rect 39374 436294 39430 436350
rect 39498 436294 39554 436350
rect 39622 436294 39678 436350
rect 39250 436170 39306 436226
rect 39374 436170 39430 436226
rect 39498 436170 39554 436226
rect 39622 436170 39678 436226
rect 39250 436046 39306 436102
rect 39374 436046 39430 436102
rect 39498 436046 39554 436102
rect 39622 436046 39678 436102
rect 39250 435922 39306 435978
rect 39374 435922 39430 435978
rect 39498 435922 39554 435978
rect 39622 435922 39678 435978
rect 39250 418294 39306 418350
rect 39374 418294 39430 418350
rect 39498 418294 39554 418350
rect 39622 418294 39678 418350
rect 39250 418170 39306 418226
rect 39374 418170 39430 418226
rect 39498 418170 39554 418226
rect 39622 418170 39678 418226
rect 39250 418046 39306 418102
rect 39374 418046 39430 418102
rect 39498 418046 39554 418102
rect 39622 418046 39678 418102
rect 39250 417922 39306 417978
rect 39374 417922 39430 417978
rect 39498 417922 39554 417978
rect 39622 417922 39678 417978
rect 39250 400294 39306 400350
rect 39374 400294 39430 400350
rect 39498 400294 39554 400350
rect 39622 400294 39678 400350
rect 39250 400170 39306 400226
rect 39374 400170 39430 400226
rect 39498 400170 39554 400226
rect 39622 400170 39678 400226
rect 39250 400046 39306 400102
rect 39374 400046 39430 400102
rect 39498 400046 39554 400102
rect 39622 400046 39678 400102
rect 39250 399922 39306 399978
rect 39374 399922 39430 399978
rect 39498 399922 39554 399978
rect 39622 399922 39678 399978
rect 39250 382294 39306 382350
rect 39374 382294 39430 382350
rect 39498 382294 39554 382350
rect 39622 382294 39678 382350
rect 39250 382170 39306 382226
rect 39374 382170 39430 382226
rect 39498 382170 39554 382226
rect 39622 382170 39678 382226
rect 39250 382046 39306 382102
rect 39374 382046 39430 382102
rect 39498 382046 39554 382102
rect 39622 382046 39678 382102
rect 39250 381922 39306 381978
rect 39374 381922 39430 381978
rect 39498 381922 39554 381978
rect 39622 381922 39678 381978
rect 39250 364294 39306 364350
rect 39374 364294 39430 364350
rect 39498 364294 39554 364350
rect 39622 364294 39678 364350
rect 39250 364170 39306 364226
rect 39374 364170 39430 364226
rect 39498 364170 39554 364226
rect 39622 364170 39678 364226
rect 39250 364046 39306 364102
rect 39374 364046 39430 364102
rect 39498 364046 39554 364102
rect 39622 364046 39678 364102
rect 39250 363922 39306 363978
rect 39374 363922 39430 363978
rect 39498 363922 39554 363978
rect 39622 363922 39678 363978
rect 39250 346294 39306 346350
rect 39374 346294 39430 346350
rect 39498 346294 39554 346350
rect 39622 346294 39678 346350
rect 39250 346170 39306 346226
rect 39374 346170 39430 346226
rect 39498 346170 39554 346226
rect 39622 346170 39678 346226
rect 39250 346046 39306 346102
rect 39374 346046 39430 346102
rect 39498 346046 39554 346102
rect 39622 346046 39678 346102
rect 39250 345922 39306 345978
rect 39374 345922 39430 345978
rect 39498 345922 39554 345978
rect 39622 345922 39678 345978
rect 39250 328294 39306 328350
rect 39374 328294 39430 328350
rect 39498 328294 39554 328350
rect 39622 328294 39678 328350
rect 39250 328170 39306 328226
rect 39374 328170 39430 328226
rect 39498 328170 39554 328226
rect 39622 328170 39678 328226
rect 39250 328046 39306 328102
rect 39374 328046 39430 328102
rect 39498 328046 39554 328102
rect 39622 328046 39678 328102
rect 39250 327922 39306 327978
rect 39374 327922 39430 327978
rect 39498 327922 39554 327978
rect 39622 327922 39678 327978
rect 39250 310294 39306 310350
rect 39374 310294 39430 310350
rect 39498 310294 39554 310350
rect 39622 310294 39678 310350
rect 39250 310170 39306 310226
rect 39374 310170 39430 310226
rect 39498 310170 39554 310226
rect 39622 310170 39678 310226
rect 39250 310046 39306 310102
rect 39374 310046 39430 310102
rect 39498 310046 39554 310102
rect 39622 310046 39678 310102
rect 39250 309922 39306 309978
rect 39374 309922 39430 309978
rect 39498 309922 39554 309978
rect 39622 309922 39678 309978
rect 39250 292294 39306 292350
rect 39374 292294 39430 292350
rect 39498 292294 39554 292350
rect 39622 292294 39678 292350
rect 39250 292170 39306 292226
rect 39374 292170 39430 292226
rect 39498 292170 39554 292226
rect 39622 292170 39678 292226
rect 39250 292046 39306 292102
rect 39374 292046 39430 292102
rect 39498 292046 39554 292102
rect 39622 292046 39678 292102
rect 39250 291922 39306 291978
rect 39374 291922 39430 291978
rect 39498 291922 39554 291978
rect 39622 291922 39678 291978
rect 39250 274294 39306 274350
rect 39374 274294 39430 274350
rect 39498 274294 39554 274350
rect 39622 274294 39678 274350
rect 39250 274170 39306 274226
rect 39374 274170 39430 274226
rect 39498 274170 39554 274226
rect 39622 274170 39678 274226
rect 39250 274046 39306 274102
rect 39374 274046 39430 274102
rect 39498 274046 39554 274102
rect 39622 274046 39678 274102
rect 39250 273922 39306 273978
rect 39374 273922 39430 273978
rect 39498 273922 39554 273978
rect 39622 273922 39678 273978
rect 39250 256294 39306 256350
rect 39374 256294 39430 256350
rect 39498 256294 39554 256350
rect 39622 256294 39678 256350
rect 39250 256170 39306 256226
rect 39374 256170 39430 256226
rect 39498 256170 39554 256226
rect 39622 256170 39678 256226
rect 39250 256046 39306 256102
rect 39374 256046 39430 256102
rect 39498 256046 39554 256102
rect 39622 256046 39678 256102
rect 39250 255922 39306 255978
rect 39374 255922 39430 255978
rect 39498 255922 39554 255978
rect 39622 255922 39678 255978
rect 39250 238294 39306 238350
rect 39374 238294 39430 238350
rect 39498 238294 39554 238350
rect 39622 238294 39678 238350
rect 39250 238170 39306 238226
rect 39374 238170 39430 238226
rect 39498 238170 39554 238226
rect 39622 238170 39678 238226
rect 39250 238046 39306 238102
rect 39374 238046 39430 238102
rect 39498 238046 39554 238102
rect 39622 238046 39678 238102
rect 39250 237922 39306 237978
rect 39374 237922 39430 237978
rect 39498 237922 39554 237978
rect 39622 237922 39678 237978
rect 39250 220294 39306 220350
rect 39374 220294 39430 220350
rect 39498 220294 39554 220350
rect 39622 220294 39678 220350
rect 39250 220170 39306 220226
rect 39374 220170 39430 220226
rect 39498 220170 39554 220226
rect 39622 220170 39678 220226
rect 39250 220046 39306 220102
rect 39374 220046 39430 220102
rect 39498 220046 39554 220102
rect 39622 220046 39678 220102
rect 39250 219922 39306 219978
rect 39374 219922 39430 219978
rect 39498 219922 39554 219978
rect 39622 219922 39678 219978
rect 39250 202294 39306 202350
rect 39374 202294 39430 202350
rect 39498 202294 39554 202350
rect 39622 202294 39678 202350
rect 39250 202170 39306 202226
rect 39374 202170 39430 202226
rect 39498 202170 39554 202226
rect 39622 202170 39678 202226
rect 39250 202046 39306 202102
rect 39374 202046 39430 202102
rect 39498 202046 39554 202102
rect 39622 202046 39678 202102
rect 39250 201922 39306 201978
rect 39374 201922 39430 201978
rect 39498 201922 39554 201978
rect 39622 201922 39678 201978
rect 39250 184294 39306 184350
rect 39374 184294 39430 184350
rect 39498 184294 39554 184350
rect 39622 184294 39678 184350
rect 39250 184170 39306 184226
rect 39374 184170 39430 184226
rect 39498 184170 39554 184226
rect 39622 184170 39678 184226
rect 39250 184046 39306 184102
rect 39374 184046 39430 184102
rect 39498 184046 39554 184102
rect 39622 184046 39678 184102
rect 39250 183922 39306 183978
rect 39374 183922 39430 183978
rect 39498 183922 39554 183978
rect 39622 183922 39678 183978
rect 39250 166294 39306 166350
rect 39374 166294 39430 166350
rect 39498 166294 39554 166350
rect 39622 166294 39678 166350
rect 39250 166170 39306 166226
rect 39374 166170 39430 166226
rect 39498 166170 39554 166226
rect 39622 166170 39678 166226
rect 39250 166046 39306 166102
rect 39374 166046 39430 166102
rect 39498 166046 39554 166102
rect 39622 166046 39678 166102
rect 39250 165922 39306 165978
rect 39374 165922 39430 165978
rect 39498 165922 39554 165978
rect 39622 165922 39678 165978
rect 39250 148294 39306 148350
rect 39374 148294 39430 148350
rect 39498 148294 39554 148350
rect 39622 148294 39678 148350
rect 39250 148170 39306 148226
rect 39374 148170 39430 148226
rect 39498 148170 39554 148226
rect 39622 148170 39678 148226
rect 39250 148046 39306 148102
rect 39374 148046 39430 148102
rect 39498 148046 39554 148102
rect 39622 148046 39678 148102
rect 39250 147922 39306 147978
rect 39374 147922 39430 147978
rect 39498 147922 39554 147978
rect 39622 147922 39678 147978
rect 39250 130294 39306 130350
rect 39374 130294 39430 130350
rect 39498 130294 39554 130350
rect 39622 130294 39678 130350
rect 39250 130170 39306 130226
rect 39374 130170 39430 130226
rect 39498 130170 39554 130226
rect 39622 130170 39678 130226
rect 39250 130046 39306 130102
rect 39374 130046 39430 130102
rect 39498 130046 39554 130102
rect 39622 130046 39678 130102
rect 39250 129922 39306 129978
rect 39374 129922 39430 129978
rect 39498 129922 39554 129978
rect 39622 129922 39678 129978
rect 39250 112294 39306 112350
rect 39374 112294 39430 112350
rect 39498 112294 39554 112350
rect 39622 112294 39678 112350
rect 39250 112170 39306 112226
rect 39374 112170 39430 112226
rect 39498 112170 39554 112226
rect 39622 112170 39678 112226
rect 39250 112046 39306 112102
rect 39374 112046 39430 112102
rect 39498 112046 39554 112102
rect 39622 112046 39678 112102
rect 39250 111922 39306 111978
rect 39374 111922 39430 111978
rect 39498 111922 39554 111978
rect 39622 111922 39678 111978
rect 39250 94294 39306 94350
rect 39374 94294 39430 94350
rect 39498 94294 39554 94350
rect 39622 94294 39678 94350
rect 39250 94170 39306 94226
rect 39374 94170 39430 94226
rect 39498 94170 39554 94226
rect 39622 94170 39678 94226
rect 39250 94046 39306 94102
rect 39374 94046 39430 94102
rect 39498 94046 39554 94102
rect 39622 94046 39678 94102
rect 39250 93922 39306 93978
rect 39374 93922 39430 93978
rect 39498 93922 39554 93978
rect 39622 93922 39678 93978
rect 39250 76294 39306 76350
rect 39374 76294 39430 76350
rect 39498 76294 39554 76350
rect 39622 76294 39678 76350
rect 39250 76170 39306 76226
rect 39374 76170 39430 76226
rect 39498 76170 39554 76226
rect 39622 76170 39678 76226
rect 39250 76046 39306 76102
rect 39374 76046 39430 76102
rect 39498 76046 39554 76102
rect 39622 76046 39678 76102
rect 39250 75922 39306 75978
rect 39374 75922 39430 75978
rect 39498 75922 39554 75978
rect 39622 75922 39678 75978
rect 39250 58294 39306 58350
rect 39374 58294 39430 58350
rect 39498 58294 39554 58350
rect 39622 58294 39678 58350
rect 39250 58170 39306 58226
rect 39374 58170 39430 58226
rect 39498 58170 39554 58226
rect 39622 58170 39678 58226
rect 39250 58046 39306 58102
rect 39374 58046 39430 58102
rect 39498 58046 39554 58102
rect 39622 58046 39678 58102
rect 39250 57922 39306 57978
rect 39374 57922 39430 57978
rect 39498 57922 39554 57978
rect 39622 57922 39678 57978
rect 39250 40294 39306 40350
rect 39374 40294 39430 40350
rect 39498 40294 39554 40350
rect 39622 40294 39678 40350
rect 39250 40170 39306 40226
rect 39374 40170 39430 40226
rect 39498 40170 39554 40226
rect 39622 40170 39678 40226
rect 39250 40046 39306 40102
rect 39374 40046 39430 40102
rect 39498 40046 39554 40102
rect 39622 40046 39678 40102
rect 39250 39922 39306 39978
rect 39374 39922 39430 39978
rect 39498 39922 39554 39978
rect 39622 39922 39678 39978
rect 39250 22294 39306 22350
rect 39374 22294 39430 22350
rect 39498 22294 39554 22350
rect 39622 22294 39678 22350
rect 39250 22170 39306 22226
rect 39374 22170 39430 22226
rect 39498 22170 39554 22226
rect 39622 22170 39678 22226
rect 39250 22046 39306 22102
rect 39374 22046 39430 22102
rect 39498 22046 39554 22102
rect 39622 22046 39678 22102
rect 39250 21922 39306 21978
rect 39374 21922 39430 21978
rect 39498 21922 39554 21978
rect 39622 21922 39678 21978
rect 39250 4294 39306 4350
rect 39374 4294 39430 4350
rect 39498 4294 39554 4350
rect 39622 4294 39678 4350
rect 39250 4170 39306 4226
rect 39374 4170 39430 4226
rect 39498 4170 39554 4226
rect 39622 4170 39678 4226
rect 39250 4046 39306 4102
rect 39374 4046 39430 4102
rect 39498 4046 39554 4102
rect 39622 4046 39678 4102
rect 39250 3922 39306 3978
rect 39374 3922 39430 3978
rect 39498 3922 39554 3978
rect 39622 3922 39678 3978
rect 39250 -216 39306 -160
rect 39374 -216 39430 -160
rect 39498 -216 39554 -160
rect 39622 -216 39678 -160
rect 39250 -340 39306 -284
rect 39374 -340 39430 -284
rect 39498 -340 39554 -284
rect 39622 -340 39678 -284
rect 39250 -464 39306 -408
rect 39374 -464 39430 -408
rect 39498 -464 39554 -408
rect 39622 -464 39678 -408
rect 39250 -588 39306 -532
rect 39374 -588 39430 -532
rect 39498 -588 39554 -532
rect 39622 -588 39678 -532
rect 42970 598116 43026 598172
rect 43094 598116 43150 598172
rect 43218 598116 43274 598172
rect 43342 598116 43398 598172
rect 42970 597992 43026 598048
rect 43094 597992 43150 598048
rect 43218 597992 43274 598048
rect 43342 597992 43398 598048
rect 42970 597868 43026 597924
rect 43094 597868 43150 597924
rect 43218 597868 43274 597924
rect 43342 597868 43398 597924
rect 42970 597744 43026 597800
rect 43094 597744 43150 597800
rect 43218 597744 43274 597800
rect 43342 597744 43398 597800
rect 42970 586294 43026 586350
rect 43094 586294 43150 586350
rect 43218 586294 43274 586350
rect 43342 586294 43398 586350
rect 42970 586170 43026 586226
rect 43094 586170 43150 586226
rect 43218 586170 43274 586226
rect 43342 586170 43398 586226
rect 42970 586046 43026 586102
rect 43094 586046 43150 586102
rect 43218 586046 43274 586102
rect 43342 586046 43398 586102
rect 42970 585922 43026 585978
rect 43094 585922 43150 585978
rect 43218 585922 43274 585978
rect 43342 585922 43398 585978
rect 42970 568294 43026 568350
rect 43094 568294 43150 568350
rect 43218 568294 43274 568350
rect 43342 568294 43398 568350
rect 42970 568170 43026 568226
rect 43094 568170 43150 568226
rect 43218 568170 43274 568226
rect 43342 568170 43398 568226
rect 42970 568046 43026 568102
rect 43094 568046 43150 568102
rect 43218 568046 43274 568102
rect 43342 568046 43398 568102
rect 42970 567922 43026 567978
rect 43094 567922 43150 567978
rect 43218 567922 43274 567978
rect 43342 567922 43398 567978
rect 42970 550294 43026 550350
rect 43094 550294 43150 550350
rect 43218 550294 43274 550350
rect 43342 550294 43398 550350
rect 42970 550170 43026 550226
rect 43094 550170 43150 550226
rect 43218 550170 43274 550226
rect 43342 550170 43398 550226
rect 42970 550046 43026 550102
rect 43094 550046 43150 550102
rect 43218 550046 43274 550102
rect 43342 550046 43398 550102
rect 42970 549922 43026 549978
rect 43094 549922 43150 549978
rect 43218 549922 43274 549978
rect 43342 549922 43398 549978
rect 42970 532294 43026 532350
rect 43094 532294 43150 532350
rect 43218 532294 43274 532350
rect 43342 532294 43398 532350
rect 42970 532170 43026 532226
rect 43094 532170 43150 532226
rect 43218 532170 43274 532226
rect 43342 532170 43398 532226
rect 42970 532046 43026 532102
rect 43094 532046 43150 532102
rect 43218 532046 43274 532102
rect 43342 532046 43398 532102
rect 42970 531922 43026 531978
rect 43094 531922 43150 531978
rect 43218 531922 43274 531978
rect 43342 531922 43398 531978
rect 42970 514294 43026 514350
rect 43094 514294 43150 514350
rect 43218 514294 43274 514350
rect 43342 514294 43398 514350
rect 42970 514170 43026 514226
rect 43094 514170 43150 514226
rect 43218 514170 43274 514226
rect 43342 514170 43398 514226
rect 42970 514046 43026 514102
rect 43094 514046 43150 514102
rect 43218 514046 43274 514102
rect 43342 514046 43398 514102
rect 42970 513922 43026 513978
rect 43094 513922 43150 513978
rect 43218 513922 43274 513978
rect 43342 513922 43398 513978
rect 42970 496294 43026 496350
rect 43094 496294 43150 496350
rect 43218 496294 43274 496350
rect 43342 496294 43398 496350
rect 42970 496170 43026 496226
rect 43094 496170 43150 496226
rect 43218 496170 43274 496226
rect 43342 496170 43398 496226
rect 42970 496046 43026 496102
rect 43094 496046 43150 496102
rect 43218 496046 43274 496102
rect 43342 496046 43398 496102
rect 42970 495922 43026 495978
rect 43094 495922 43150 495978
rect 43218 495922 43274 495978
rect 43342 495922 43398 495978
rect 42970 478294 43026 478350
rect 43094 478294 43150 478350
rect 43218 478294 43274 478350
rect 43342 478294 43398 478350
rect 42970 478170 43026 478226
rect 43094 478170 43150 478226
rect 43218 478170 43274 478226
rect 43342 478170 43398 478226
rect 42970 478046 43026 478102
rect 43094 478046 43150 478102
rect 43218 478046 43274 478102
rect 43342 478046 43398 478102
rect 42970 477922 43026 477978
rect 43094 477922 43150 477978
rect 43218 477922 43274 477978
rect 43342 477922 43398 477978
rect 42970 460294 43026 460350
rect 43094 460294 43150 460350
rect 43218 460294 43274 460350
rect 43342 460294 43398 460350
rect 42970 460170 43026 460226
rect 43094 460170 43150 460226
rect 43218 460170 43274 460226
rect 43342 460170 43398 460226
rect 42970 460046 43026 460102
rect 43094 460046 43150 460102
rect 43218 460046 43274 460102
rect 43342 460046 43398 460102
rect 42970 459922 43026 459978
rect 43094 459922 43150 459978
rect 43218 459922 43274 459978
rect 43342 459922 43398 459978
rect 42970 442294 43026 442350
rect 43094 442294 43150 442350
rect 43218 442294 43274 442350
rect 43342 442294 43398 442350
rect 42970 442170 43026 442226
rect 43094 442170 43150 442226
rect 43218 442170 43274 442226
rect 43342 442170 43398 442226
rect 42970 442046 43026 442102
rect 43094 442046 43150 442102
rect 43218 442046 43274 442102
rect 43342 442046 43398 442102
rect 42970 441922 43026 441978
rect 43094 441922 43150 441978
rect 43218 441922 43274 441978
rect 43342 441922 43398 441978
rect 42970 424294 43026 424350
rect 43094 424294 43150 424350
rect 43218 424294 43274 424350
rect 43342 424294 43398 424350
rect 42970 424170 43026 424226
rect 43094 424170 43150 424226
rect 43218 424170 43274 424226
rect 43342 424170 43398 424226
rect 42970 424046 43026 424102
rect 43094 424046 43150 424102
rect 43218 424046 43274 424102
rect 43342 424046 43398 424102
rect 42970 423922 43026 423978
rect 43094 423922 43150 423978
rect 43218 423922 43274 423978
rect 43342 423922 43398 423978
rect 42970 406294 43026 406350
rect 43094 406294 43150 406350
rect 43218 406294 43274 406350
rect 43342 406294 43398 406350
rect 42970 406170 43026 406226
rect 43094 406170 43150 406226
rect 43218 406170 43274 406226
rect 43342 406170 43398 406226
rect 42970 406046 43026 406102
rect 43094 406046 43150 406102
rect 43218 406046 43274 406102
rect 43342 406046 43398 406102
rect 42970 405922 43026 405978
rect 43094 405922 43150 405978
rect 43218 405922 43274 405978
rect 43342 405922 43398 405978
rect 42970 388294 43026 388350
rect 43094 388294 43150 388350
rect 43218 388294 43274 388350
rect 43342 388294 43398 388350
rect 42970 388170 43026 388226
rect 43094 388170 43150 388226
rect 43218 388170 43274 388226
rect 43342 388170 43398 388226
rect 42970 388046 43026 388102
rect 43094 388046 43150 388102
rect 43218 388046 43274 388102
rect 43342 388046 43398 388102
rect 42970 387922 43026 387978
rect 43094 387922 43150 387978
rect 43218 387922 43274 387978
rect 43342 387922 43398 387978
rect 42970 370294 43026 370350
rect 43094 370294 43150 370350
rect 43218 370294 43274 370350
rect 43342 370294 43398 370350
rect 42970 370170 43026 370226
rect 43094 370170 43150 370226
rect 43218 370170 43274 370226
rect 43342 370170 43398 370226
rect 42970 370046 43026 370102
rect 43094 370046 43150 370102
rect 43218 370046 43274 370102
rect 43342 370046 43398 370102
rect 42970 369922 43026 369978
rect 43094 369922 43150 369978
rect 43218 369922 43274 369978
rect 43342 369922 43398 369978
rect 42970 352294 43026 352350
rect 43094 352294 43150 352350
rect 43218 352294 43274 352350
rect 43342 352294 43398 352350
rect 42970 352170 43026 352226
rect 43094 352170 43150 352226
rect 43218 352170 43274 352226
rect 43342 352170 43398 352226
rect 42970 352046 43026 352102
rect 43094 352046 43150 352102
rect 43218 352046 43274 352102
rect 43342 352046 43398 352102
rect 42970 351922 43026 351978
rect 43094 351922 43150 351978
rect 43218 351922 43274 351978
rect 43342 351922 43398 351978
rect 42970 334294 43026 334350
rect 43094 334294 43150 334350
rect 43218 334294 43274 334350
rect 43342 334294 43398 334350
rect 42970 334170 43026 334226
rect 43094 334170 43150 334226
rect 43218 334170 43274 334226
rect 43342 334170 43398 334226
rect 42970 334046 43026 334102
rect 43094 334046 43150 334102
rect 43218 334046 43274 334102
rect 43342 334046 43398 334102
rect 42970 333922 43026 333978
rect 43094 333922 43150 333978
rect 43218 333922 43274 333978
rect 43342 333922 43398 333978
rect 42970 316294 43026 316350
rect 43094 316294 43150 316350
rect 43218 316294 43274 316350
rect 43342 316294 43398 316350
rect 42970 316170 43026 316226
rect 43094 316170 43150 316226
rect 43218 316170 43274 316226
rect 43342 316170 43398 316226
rect 42970 316046 43026 316102
rect 43094 316046 43150 316102
rect 43218 316046 43274 316102
rect 43342 316046 43398 316102
rect 42970 315922 43026 315978
rect 43094 315922 43150 315978
rect 43218 315922 43274 315978
rect 43342 315922 43398 315978
rect 42970 298294 43026 298350
rect 43094 298294 43150 298350
rect 43218 298294 43274 298350
rect 43342 298294 43398 298350
rect 42970 298170 43026 298226
rect 43094 298170 43150 298226
rect 43218 298170 43274 298226
rect 43342 298170 43398 298226
rect 42970 298046 43026 298102
rect 43094 298046 43150 298102
rect 43218 298046 43274 298102
rect 43342 298046 43398 298102
rect 42970 297922 43026 297978
rect 43094 297922 43150 297978
rect 43218 297922 43274 297978
rect 43342 297922 43398 297978
rect 42970 280294 43026 280350
rect 43094 280294 43150 280350
rect 43218 280294 43274 280350
rect 43342 280294 43398 280350
rect 42970 280170 43026 280226
rect 43094 280170 43150 280226
rect 43218 280170 43274 280226
rect 43342 280170 43398 280226
rect 42970 280046 43026 280102
rect 43094 280046 43150 280102
rect 43218 280046 43274 280102
rect 43342 280046 43398 280102
rect 42970 279922 43026 279978
rect 43094 279922 43150 279978
rect 43218 279922 43274 279978
rect 43342 279922 43398 279978
rect 42970 262294 43026 262350
rect 43094 262294 43150 262350
rect 43218 262294 43274 262350
rect 43342 262294 43398 262350
rect 42970 262170 43026 262226
rect 43094 262170 43150 262226
rect 43218 262170 43274 262226
rect 43342 262170 43398 262226
rect 42970 262046 43026 262102
rect 43094 262046 43150 262102
rect 43218 262046 43274 262102
rect 43342 262046 43398 262102
rect 42970 261922 43026 261978
rect 43094 261922 43150 261978
rect 43218 261922 43274 261978
rect 43342 261922 43398 261978
rect 42970 244294 43026 244350
rect 43094 244294 43150 244350
rect 43218 244294 43274 244350
rect 43342 244294 43398 244350
rect 42970 244170 43026 244226
rect 43094 244170 43150 244226
rect 43218 244170 43274 244226
rect 43342 244170 43398 244226
rect 42970 244046 43026 244102
rect 43094 244046 43150 244102
rect 43218 244046 43274 244102
rect 43342 244046 43398 244102
rect 42970 243922 43026 243978
rect 43094 243922 43150 243978
rect 43218 243922 43274 243978
rect 43342 243922 43398 243978
rect 42970 226294 43026 226350
rect 43094 226294 43150 226350
rect 43218 226294 43274 226350
rect 43342 226294 43398 226350
rect 42970 226170 43026 226226
rect 43094 226170 43150 226226
rect 43218 226170 43274 226226
rect 43342 226170 43398 226226
rect 42970 226046 43026 226102
rect 43094 226046 43150 226102
rect 43218 226046 43274 226102
rect 43342 226046 43398 226102
rect 42970 225922 43026 225978
rect 43094 225922 43150 225978
rect 43218 225922 43274 225978
rect 43342 225922 43398 225978
rect 42970 208294 43026 208350
rect 43094 208294 43150 208350
rect 43218 208294 43274 208350
rect 43342 208294 43398 208350
rect 42970 208170 43026 208226
rect 43094 208170 43150 208226
rect 43218 208170 43274 208226
rect 43342 208170 43398 208226
rect 42970 208046 43026 208102
rect 43094 208046 43150 208102
rect 43218 208046 43274 208102
rect 43342 208046 43398 208102
rect 42970 207922 43026 207978
rect 43094 207922 43150 207978
rect 43218 207922 43274 207978
rect 43342 207922 43398 207978
rect 42970 190294 43026 190350
rect 43094 190294 43150 190350
rect 43218 190294 43274 190350
rect 43342 190294 43398 190350
rect 42970 190170 43026 190226
rect 43094 190170 43150 190226
rect 43218 190170 43274 190226
rect 43342 190170 43398 190226
rect 42970 190046 43026 190102
rect 43094 190046 43150 190102
rect 43218 190046 43274 190102
rect 43342 190046 43398 190102
rect 42970 189922 43026 189978
rect 43094 189922 43150 189978
rect 43218 189922 43274 189978
rect 43342 189922 43398 189978
rect 42970 172294 43026 172350
rect 43094 172294 43150 172350
rect 43218 172294 43274 172350
rect 43342 172294 43398 172350
rect 42970 172170 43026 172226
rect 43094 172170 43150 172226
rect 43218 172170 43274 172226
rect 43342 172170 43398 172226
rect 42970 172046 43026 172102
rect 43094 172046 43150 172102
rect 43218 172046 43274 172102
rect 43342 172046 43398 172102
rect 42970 171922 43026 171978
rect 43094 171922 43150 171978
rect 43218 171922 43274 171978
rect 43342 171922 43398 171978
rect 42970 154294 43026 154350
rect 43094 154294 43150 154350
rect 43218 154294 43274 154350
rect 43342 154294 43398 154350
rect 42970 154170 43026 154226
rect 43094 154170 43150 154226
rect 43218 154170 43274 154226
rect 43342 154170 43398 154226
rect 42970 154046 43026 154102
rect 43094 154046 43150 154102
rect 43218 154046 43274 154102
rect 43342 154046 43398 154102
rect 42970 153922 43026 153978
rect 43094 153922 43150 153978
rect 43218 153922 43274 153978
rect 43342 153922 43398 153978
rect 42970 136294 43026 136350
rect 43094 136294 43150 136350
rect 43218 136294 43274 136350
rect 43342 136294 43398 136350
rect 42970 136170 43026 136226
rect 43094 136170 43150 136226
rect 43218 136170 43274 136226
rect 43342 136170 43398 136226
rect 42970 136046 43026 136102
rect 43094 136046 43150 136102
rect 43218 136046 43274 136102
rect 43342 136046 43398 136102
rect 42970 135922 43026 135978
rect 43094 135922 43150 135978
rect 43218 135922 43274 135978
rect 43342 135922 43398 135978
rect 42970 118294 43026 118350
rect 43094 118294 43150 118350
rect 43218 118294 43274 118350
rect 43342 118294 43398 118350
rect 42970 118170 43026 118226
rect 43094 118170 43150 118226
rect 43218 118170 43274 118226
rect 43342 118170 43398 118226
rect 42970 118046 43026 118102
rect 43094 118046 43150 118102
rect 43218 118046 43274 118102
rect 43342 118046 43398 118102
rect 42970 117922 43026 117978
rect 43094 117922 43150 117978
rect 43218 117922 43274 117978
rect 43342 117922 43398 117978
rect 42970 100294 43026 100350
rect 43094 100294 43150 100350
rect 43218 100294 43274 100350
rect 43342 100294 43398 100350
rect 42970 100170 43026 100226
rect 43094 100170 43150 100226
rect 43218 100170 43274 100226
rect 43342 100170 43398 100226
rect 42970 100046 43026 100102
rect 43094 100046 43150 100102
rect 43218 100046 43274 100102
rect 43342 100046 43398 100102
rect 42970 99922 43026 99978
rect 43094 99922 43150 99978
rect 43218 99922 43274 99978
rect 43342 99922 43398 99978
rect 42970 82294 43026 82350
rect 43094 82294 43150 82350
rect 43218 82294 43274 82350
rect 43342 82294 43398 82350
rect 42970 82170 43026 82226
rect 43094 82170 43150 82226
rect 43218 82170 43274 82226
rect 43342 82170 43398 82226
rect 42970 82046 43026 82102
rect 43094 82046 43150 82102
rect 43218 82046 43274 82102
rect 43342 82046 43398 82102
rect 42970 81922 43026 81978
rect 43094 81922 43150 81978
rect 43218 81922 43274 81978
rect 43342 81922 43398 81978
rect 42970 64294 43026 64350
rect 43094 64294 43150 64350
rect 43218 64294 43274 64350
rect 43342 64294 43398 64350
rect 42970 64170 43026 64226
rect 43094 64170 43150 64226
rect 43218 64170 43274 64226
rect 43342 64170 43398 64226
rect 42970 64046 43026 64102
rect 43094 64046 43150 64102
rect 43218 64046 43274 64102
rect 43342 64046 43398 64102
rect 42970 63922 43026 63978
rect 43094 63922 43150 63978
rect 43218 63922 43274 63978
rect 43342 63922 43398 63978
rect 42970 46294 43026 46350
rect 43094 46294 43150 46350
rect 43218 46294 43274 46350
rect 43342 46294 43398 46350
rect 42970 46170 43026 46226
rect 43094 46170 43150 46226
rect 43218 46170 43274 46226
rect 43342 46170 43398 46226
rect 42970 46046 43026 46102
rect 43094 46046 43150 46102
rect 43218 46046 43274 46102
rect 43342 46046 43398 46102
rect 42970 45922 43026 45978
rect 43094 45922 43150 45978
rect 43218 45922 43274 45978
rect 43342 45922 43398 45978
rect 42970 28294 43026 28350
rect 43094 28294 43150 28350
rect 43218 28294 43274 28350
rect 43342 28294 43398 28350
rect 42970 28170 43026 28226
rect 43094 28170 43150 28226
rect 43218 28170 43274 28226
rect 43342 28170 43398 28226
rect 42970 28046 43026 28102
rect 43094 28046 43150 28102
rect 43218 28046 43274 28102
rect 43342 28046 43398 28102
rect 42970 27922 43026 27978
rect 43094 27922 43150 27978
rect 43218 27922 43274 27978
rect 43342 27922 43398 27978
rect 42970 10294 43026 10350
rect 43094 10294 43150 10350
rect 43218 10294 43274 10350
rect 43342 10294 43398 10350
rect 42970 10170 43026 10226
rect 43094 10170 43150 10226
rect 43218 10170 43274 10226
rect 43342 10170 43398 10226
rect 42970 10046 43026 10102
rect 43094 10046 43150 10102
rect 43218 10046 43274 10102
rect 43342 10046 43398 10102
rect 42970 9922 43026 9978
rect 43094 9922 43150 9978
rect 43218 9922 43274 9978
rect 43342 9922 43398 9978
rect 42970 -1176 43026 -1120
rect 43094 -1176 43150 -1120
rect 43218 -1176 43274 -1120
rect 43342 -1176 43398 -1120
rect 42970 -1300 43026 -1244
rect 43094 -1300 43150 -1244
rect 43218 -1300 43274 -1244
rect 43342 -1300 43398 -1244
rect 42970 -1424 43026 -1368
rect 43094 -1424 43150 -1368
rect 43218 -1424 43274 -1368
rect 43342 -1424 43398 -1368
rect 42970 -1548 43026 -1492
rect 43094 -1548 43150 -1492
rect 43218 -1548 43274 -1492
rect 43342 -1548 43398 -1492
rect 57250 597156 57306 597212
rect 57374 597156 57430 597212
rect 57498 597156 57554 597212
rect 57622 597156 57678 597212
rect 57250 597032 57306 597088
rect 57374 597032 57430 597088
rect 57498 597032 57554 597088
rect 57622 597032 57678 597088
rect 57250 596908 57306 596964
rect 57374 596908 57430 596964
rect 57498 596908 57554 596964
rect 57622 596908 57678 596964
rect 57250 596784 57306 596840
rect 57374 596784 57430 596840
rect 57498 596784 57554 596840
rect 57622 596784 57678 596840
rect 57250 580294 57306 580350
rect 57374 580294 57430 580350
rect 57498 580294 57554 580350
rect 57622 580294 57678 580350
rect 57250 580170 57306 580226
rect 57374 580170 57430 580226
rect 57498 580170 57554 580226
rect 57622 580170 57678 580226
rect 57250 580046 57306 580102
rect 57374 580046 57430 580102
rect 57498 580046 57554 580102
rect 57622 580046 57678 580102
rect 57250 579922 57306 579978
rect 57374 579922 57430 579978
rect 57498 579922 57554 579978
rect 57622 579922 57678 579978
rect 57250 562294 57306 562350
rect 57374 562294 57430 562350
rect 57498 562294 57554 562350
rect 57622 562294 57678 562350
rect 57250 562170 57306 562226
rect 57374 562170 57430 562226
rect 57498 562170 57554 562226
rect 57622 562170 57678 562226
rect 57250 562046 57306 562102
rect 57374 562046 57430 562102
rect 57498 562046 57554 562102
rect 57622 562046 57678 562102
rect 57250 561922 57306 561978
rect 57374 561922 57430 561978
rect 57498 561922 57554 561978
rect 57622 561922 57678 561978
rect 57250 544294 57306 544350
rect 57374 544294 57430 544350
rect 57498 544294 57554 544350
rect 57622 544294 57678 544350
rect 57250 544170 57306 544226
rect 57374 544170 57430 544226
rect 57498 544170 57554 544226
rect 57622 544170 57678 544226
rect 57250 544046 57306 544102
rect 57374 544046 57430 544102
rect 57498 544046 57554 544102
rect 57622 544046 57678 544102
rect 57250 543922 57306 543978
rect 57374 543922 57430 543978
rect 57498 543922 57554 543978
rect 57622 543922 57678 543978
rect 57250 526294 57306 526350
rect 57374 526294 57430 526350
rect 57498 526294 57554 526350
rect 57622 526294 57678 526350
rect 57250 526170 57306 526226
rect 57374 526170 57430 526226
rect 57498 526170 57554 526226
rect 57622 526170 57678 526226
rect 57250 526046 57306 526102
rect 57374 526046 57430 526102
rect 57498 526046 57554 526102
rect 57622 526046 57678 526102
rect 57250 525922 57306 525978
rect 57374 525922 57430 525978
rect 57498 525922 57554 525978
rect 57622 525922 57678 525978
rect 57250 508294 57306 508350
rect 57374 508294 57430 508350
rect 57498 508294 57554 508350
rect 57622 508294 57678 508350
rect 57250 508170 57306 508226
rect 57374 508170 57430 508226
rect 57498 508170 57554 508226
rect 57622 508170 57678 508226
rect 57250 508046 57306 508102
rect 57374 508046 57430 508102
rect 57498 508046 57554 508102
rect 57622 508046 57678 508102
rect 57250 507922 57306 507978
rect 57374 507922 57430 507978
rect 57498 507922 57554 507978
rect 57622 507922 57678 507978
rect 57250 490294 57306 490350
rect 57374 490294 57430 490350
rect 57498 490294 57554 490350
rect 57622 490294 57678 490350
rect 57250 490170 57306 490226
rect 57374 490170 57430 490226
rect 57498 490170 57554 490226
rect 57622 490170 57678 490226
rect 57250 490046 57306 490102
rect 57374 490046 57430 490102
rect 57498 490046 57554 490102
rect 57622 490046 57678 490102
rect 57250 489922 57306 489978
rect 57374 489922 57430 489978
rect 57498 489922 57554 489978
rect 57622 489922 57678 489978
rect 57250 472294 57306 472350
rect 57374 472294 57430 472350
rect 57498 472294 57554 472350
rect 57622 472294 57678 472350
rect 57250 472170 57306 472226
rect 57374 472170 57430 472226
rect 57498 472170 57554 472226
rect 57622 472170 57678 472226
rect 57250 472046 57306 472102
rect 57374 472046 57430 472102
rect 57498 472046 57554 472102
rect 57622 472046 57678 472102
rect 57250 471922 57306 471978
rect 57374 471922 57430 471978
rect 57498 471922 57554 471978
rect 57622 471922 57678 471978
rect 57250 454294 57306 454350
rect 57374 454294 57430 454350
rect 57498 454294 57554 454350
rect 57622 454294 57678 454350
rect 57250 454170 57306 454226
rect 57374 454170 57430 454226
rect 57498 454170 57554 454226
rect 57622 454170 57678 454226
rect 57250 454046 57306 454102
rect 57374 454046 57430 454102
rect 57498 454046 57554 454102
rect 57622 454046 57678 454102
rect 57250 453922 57306 453978
rect 57374 453922 57430 453978
rect 57498 453922 57554 453978
rect 57622 453922 57678 453978
rect 57250 436294 57306 436350
rect 57374 436294 57430 436350
rect 57498 436294 57554 436350
rect 57622 436294 57678 436350
rect 57250 436170 57306 436226
rect 57374 436170 57430 436226
rect 57498 436170 57554 436226
rect 57622 436170 57678 436226
rect 57250 436046 57306 436102
rect 57374 436046 57430 436102
rect 57498 436046 57554 436102
rect 57622 436046 57678 436102
rect 57250 435922 57306 435978
rect 57374 435922 57430 435978
rect 57498 435922 57554 435978
rect 57622 435922 57678 435978
rect 57250 418294 57306 418350
rect 57374 418294 57430 418350
rect 57498 418294 57554 418350
rect 57622 418294 57678 418350
rect 57250 418170 57306 418226
rect 57374 418170 57430 418226
rect 57498 418170 57554 418226
rect 57622 418170 57678 418226
rect 57250 418046 57306 418102
rect 57374 418046 57430 418102
rect 57498 418046 57554 418102
rect 57622 418046 57678 418102
rect 57250 417922 57306 417978
rect 57374 417922 57430 417978
rect 57498 417922 57554 417978
rect 57622 417922 57678 417978
rect 57250 400294 57306 400350
rect 57374 400294 57430 400350
rect 57498 400294 57554 400350
rect 57622 400294 57678 400350
rect 57250 400170 57306 400226
rect 57374 400170 57430 400226
rect 57498 400170 57554 400226
rect 57622 400170 57678 400226
rect 57250 400046 57306 400102
rect 57374 400046 57430 400102
rect 57498 400046 57554 400102
rect 57622 400046 57678 400102
rect 57250 399922 57306 399978
rect 57374 399922 57430 399978
rect 57498 399922 57554 399978
rect 57622 399922 57678 399978
rect 57250 382294 57306 382350
rect 57374 382294 57430 382350
rect 57498 382294 57554 382350
rect 57622 382294 57678 382350
rect 57250 382170 57306 382226
rect 57374 382170 57430 382226
rect 57498 382170 57554 382226
rect 57622 382170 57678 382226
rect 57250 382046 57306 382102
rect 57374 382046 57430 382102
rect 57498 382046 57554 382102
rect 57622 382046 57678 382102
rect 57250 381922 57306 381978
rect 57374 381922 57430 381978
rect 57498 381922 57554 381978
rect 57622 381922 57678 381978
rect 57250 364294 57306 364350
rect 57374 364294 57430 364350
rect 57498 364294 57554 364350
rect 57622 364294 57678 364350
rect 57250 364170 57306 364226
rect 57374 364170 57430 364226
rect 57498 364170 57554 364226
rect 57622 364170 57678 364226
rect 57250 364046 57306 364102
rect 57374 364046 57430 364102
rect 57498 364046 57554 364102
rect 57622 364046 57678 364102
rect 57250 363922 57306 363978
rect 57374 363922 57430 363978
rect 57498 363922 57554 363978
rect 57622 363922 57678 363978
rect 57250 346294 57306 346350
rect 57374 346294 57430 346350
rect 57498 346294 57554 346350
rect 57622 346294 57678 346350
rect 57250 346170 57306 346226
rect 57374 346170 57430 346226
rect 57498 346170 57554 346226
rect 57622 346170 57678 346226
rect 57250 346046 57306 346102
rect 57374 346046 57430 346102
rect 57498 346046 57554 346102
rect 57622 346046 57678 346102
rect 57250 345922 57306 345978
rect 57374 345922 57430 345978
rect 57498 345922 57554 345978
rect 57622 345922 57678 345978
rect 57250 328294 57306 328350
rect 57374 328294 57430 328350
rect 57498 328294 57554 328350
rect 57622 328294 57678 328350
rect 57250 328170 57306 328226
rect 57374 328170 57430 328226
rect 57498 328170 57554 328226
rect 57622 328170 57678 328226
rect 57250 328046 57306 328102
rect 57374 328046 57430 328102
rect 57498 328046 57554 328102
rect 57622 328046 57678 328102
rect 57250 327922 57306 327978
rect 57374 327922 57430 327978
rect 57498 327922 57554 327978
rect 57622 327922 57678 327978
rect 57250 310294 57306 310350
rect 57374 310294 57430 310350
rect 57498 310294 57554 310350
rect 57622 310294 57678 310350
rect 57250 310170 57306 310226
rect 57374 310170 57430 310226
rect 57498 310170 57554 310226
rect 57622 310170 57678 310226
rect 57250 310046 57306 310102
rect 57374 310046 57430 310102
rect 57498 310046 57554 310102
rect 57622 310046 57678 310102
rect 57250 309922 57306 309978
rect 57374 309922 57430 309978
rect 57498 309922 57554 309978
rect 57622 309922 57678 309978
rect 57250 292294 57306 292350
rect 57374 292294 57430 292350
rect 57498 292294 57554 292350
rect 57622 292294 57678 292350
rect 57250 292170 57306 292226
rect 57374 292170 57430 292226
rect 57498 292170 57554 292226
rect 57622 292170 57678 292226
rect 57250 292046 57306 292102
rect 57374 292046 57430 292102
rect 57498 292046 57554 292102
rect 57622 292046 57678 292102
rect 57250 291922 57306 291978
rect 57374 291922 57430 291978
rect 57498 291922 57554 291978
rect 57622 291922 57678 291978
rect 57250 274294 57306 274350
rect 57374 274294 57430 274350
rect 57498 274294 57554 274350
rect 57622 274294 57678 274350
rect 57250 274170 57306 274226
rect 57374 274170 57430 274226
rect 57498 274170 57554 274226
rect 57622 274170 57678 274226
rect 57250 274046 57306 274102
rect 57374 274046 57430 274102
rect 57498 274046 57554 274102
rect 57622 274046 57678 274102
rect 57250 273922 57306 273978
rect 57374 273922 57430 273978
rect 57498 273922 57554 273978
rect 57622 273922 57678 273978
rect 57250 256294 57306 256350
rect 57374 256294 57430 256350
rect 57498 256294 57554 256350
rect 57622 256294 57678 256350
rect 57250 256170 57306 256226
rect 57374 256170 57430 256226
rect 57498 256170 57554 256226
rect 57622 256170 57678 256226
rect 57250 256046 57306 256102
rect 57374 256046 57430 256102
rect 57498 256046 57554 256102
rect 57622 256046 57678 256102
rect 57250 255922 57306 255978
rect 57374 255922 57430 255978
rect 57498 255922 57554 255978
rect 57622 255922 57678 255978
rect 57250 238294 57306 238350
rect 57374 238294 57430 238350
rect 57498 238294 57554 238350
rect 57622 238294 57678 238350
rect 57250 238170 57306 238226
rect 57374 238170 57430 238226
rect 57498 238170 57554 238226
rect 57622 238170 57678 238226
rect 57250 238046 57306 238102
rect 57374 238046 57430 238102
rect 57498 238046 57554 238102
rect 57622 238046 57678 238102
rect 57250 237922 57306 237978
rect 57374 237922 57430 237978
rect 57498 237922 57554 237978
rect 57622 237922 57678 237978
rect 57250 220294 57306 220350
rect 57374 220294 57430 220350
rect 57498 220294 57554 220350
rect 57622 220294 57678 220350
rect 57250 220170 57306 220226
rect 57374 220170 57430 220226
rect 57498 220170 57554 220226
rect 57622 220170 57678 220226
rect 57250 220046 57306 220102
rect 57374 220046 57430 220102
rect 57498 220046 57554 220102
rect 57622 220046 57678 220102
rect 57250 219922 57306 219978
rect 57374 219922 57430 219978
rect 57498 219922 57554 219978
rect 57622 219922 57678 219978
rect 57250 202294 57306 202350
rect 57374 202294 57430 202350
rect 57498 202294 57554 202350
rect 57622 202294 57678 202350
rect 57250 202170 57306 202226
rect 57374 202170 57430 202226
rect 57498 202170 57554 202226
rect 57622 202170 57678 202226
rect 57250 202046 57306 202102
rect 57374 202046 57430 202102
rect 57498 202046 57554 202102
rect 57622 202046 57678 202102
rect 57250 201922 57306 201978
rect 57374 201922 57430 201978
rect 57498 201922 57554 201978
rect 57622 201922 57678 201978
rect 57250 184294 57306 184350
rect 57374 184294 57430 184350
rect 57498 184294 57554 184350
rect 57622 184294 57678 184350
rect 57250 184170 57306 184226
rect 57374 184170 57430 184226
rect 57498 184170 57554 184226
rect 57622 184170 57678 184226
rect 57250 184046 57306 184102
rect 57374 184046 57430 184102
rect 57498 184046 57554 184102
rect 57622 184046 57678 184102
rect 57250 183922 57306 183978
rect 57374 183922 57430 183978
rect 57498 183922 57554 183978
rect 57622 183922 57678 183978
rect 57250 166294 57306 166350
rect 57374 166294 57430 166350
rect 57498 166294 57554 166350
rect 57622 166294 57678 166350
rect 57250 166170 57306 166226
rect 57374 166170 57430 166226
rect 57498 166170 57554 166226
rect 57622 166170 57678 166226
rect 57250 166046 57306 166102
rect 57374 166046 57430 166102
rect 57498 166046 57554 166102
rect 57622 166046 57678 166102
rect 57250 165922 57306 165978
rect 57374 165922 57430 165978
rect 57498 165922 57554 165978
rect 57622 165922 57678 165978
rect 57250 148294 57306 148350
rect 57374 148294 57430 148350
rect 57498 148294 57554 148350
rect 57622 148294 57678 148350
rect 57250 148170 57306 148226
rect 57374 148170 57430 148226
rect 57498 148170 57554 148226
rect 57622 148170 57678 148226
rect 57250 148046 57306 148102
rect 57374 148046 57430 148102
rect 57498 148046 57554 148102
rect 57622 148046 57678 148102
rect 57250 147922 57306 147978
rect 57374 147922 57430 147978
rect 57498 147922 57554 147978
rect 57622 147922 57678 147978
rect 57250 130294 57306 130350
rect 57374 130294 57430 130350
rect 57498 130294 57554 130350
rect 57622 130294 57678 130350
rect 57250 130170 57306 130226
rect 57374 130170 57430 130226
rect 57498 130170 57554 130226
rect 57622 130170 57678 130226
rect 57250 130046 57306 130102
rect 57374 130046 57430 130102
rect 57498 130046 57554 130102
rect 57622 130046 57678 130102
rect 57250 129922 57306 129978
rect 57374 129922 57430 129978
rect 57498 129922 57554 129978
rect 57622 129922 57678 129978
rect 57250 112294 57306 112350
rect 57374 112294 57430 112350
rect 57498 112294 57554 112350
rect 57622 112294 57678 112350
rect 57250 112170 57306 112226
rect 57374 112170 57430 112226
rect 57498 112170 57554 112226
rect 57622 112170 57678 112226
rect 57250 112046 57306 112102
rect 57374 112046 57430 112102
rect 57498 112046 57554 112102
rect 57622 112046 57678 112102
rect 57250 111922 57306 111978
rect 57374 111922 57430 111978
rect 57498 111922 57554 111978
rect 57622 111922 57678 111978
rect 57250 94294 57306 94350
rect 57374 94294 57430 94350
rect 57498 94294 57554 94350
rect 57622 94294 57678 94350
rect 57250 94170 57306 94226
rect 57374 94170 57430 94226
rect 57498 94170 57554 94226
rect 57622 94170 57678 94226
rect 57250 94046 57306 94102
rect 57374 94046 57430 94102
rect 57498 94046 57554 94102
rect 57622 94046 57678 94102
rect 57250 93922 57306 93978
rect 57374 93922 57430 93978
rect 57498 93922 57554 93978
rect 57622 93922 57678 93978
rect 57250 76294 57306 76350
rect 57374 76294 57430 76350
rect 57498 76294 57554 76350
rect 57622 76294 57678 76350
rect 57250 76170 57306 76226
rect 57374 76170 57430 76226
rect 57498 76170 57554 76226
rect 57622 76170 57678 76226
rect 57250 76046 57306 76102
rect 57374 76046 57430 76102
rect 57498 76046 57554 76102
rect 57622 76046 57678 76102
rect 57250 75922 57306 75978
rect 57374 75922 57430 75978
rect 57498 75922 57554 75978
rect 57622 75922 57678 75978
rect 57250 58294 57306 58350
rect 57374 58294 57430 58350
rect 57498 58294 57554 58350
rect 57622 58294 57678 58350
rect 57250 58170 57306 58226
rect 57374 58170 57430 58226
rect 57498 58170 57554 58226
rect 57622 58170 57678 58226
rect 57250 58046 57306 58102
rect 57374 58046 57430 58102
rect 57498 58046 57554 58102
rect 57622 58046 57678 58102
rect 57250 57922 57306 57978
rect 57374 57922 57430 57978
rect 57498 57922 57554 57978
rect 57622 57922 57678 57978
rect 57250 40294 57306 40350
rect 57374 40294 57430 40350
rect 57498 40294 57554 40350
rect 57622 40294 57678 40350
rect 57250 40170 57306 40226
rect 57374 40170 57430 40226
rect 57498 40170 57554 40226
rect 57622 40170 57678 40226
rect 57250 40046 57306 40102
rect 57374 40046 57430 40102
rect 57498 40046 57554 40102
rect 57622 40046 57678 40102
rect 57250 39922 57306 39978
rect 57374 39922 57430 39978
rect 57498 39922 57554 39978
rect 57622 39922 57678 39978
rect 57250 22294 57306 22350
rect 57374 22294 57430 22350
rect 57498 22294 57554 22350
rect 57622 22294 57678 22350
rect 57250 22170 57306 22226
rect 57374 22170 57430 22226
rect 57498 22170 57554 22226
rect 57622 22170 57678 22226
rect 57250 22046 57306 22102
rect 57374 22046 57430 22102
rect 57498 22046 57554 22102
rect 57622 22046 57678 22102
rect 57250 21922 57306 21978
rect 57374 21922 57430 21978
rect 57498 21922 57554 21978
rect 57622 21922 57678 21978
rect 57250 4294 57306 4350
rect 57374 4294 57430 4350
rect 57498 4294 57554 4350
rect 57622 4294 57678 4350
rect 57250 4170 57306 4226
rect 57374 4170 57430 4226
rect 57498 4170 57554 4226
rect 57622 4170 57678 4226
rect 57250 4046 57306 4102
rect 57374 4046 57430 4102
rect 57498 4046 57554 4102
rect 57622 4046 57678 4102
rect 57250 3922 57306 3978
rect 57374 3922 57430 3978
rect 57498 3922 57554 3978
rect 57622 3922 57678 3978
rect 57250 -216 57306 -160
rect 57374 -216 57430 -160
rect 57498 -216 57554 -160
rect 57622 -216 57678 -160
rect 57250 -340 57306 -284
rect 57374 -340 57430 -284
rect 57498 -340 57554 -284
rect 57622 -340 57678 -284
rect 57250 -464 57306 -408
rect 57374 -464 57430 -408
rect 57498 -464 57554 -408
rect 57622 -464 57678 -408
rect 57250 -588 57306 -532
rect 57374 -588 57430 -532
rect 57498 -588 57554 -532
rect 57622 -588 57678 -532
rect 60970 598116 61026 598172
rect 61094 598116 61150 598172
rect 61218 598116 61274 598172
rect 61342 598116 61398 598172
rect 60970 597992 61026 598048
rect 61094 597992 61150 598048
rect 61218 597992 61274 598048
rect 61342 597992 61398 598048
rect 60970 597868 61026 597924
rect 61094 597868 61150 597924
rect 61218 597868 61274 597924
rect 61342 597868 61398 597924
rect 60970 597744 61026 597800
rect 61094 597744 61150 597800
rect 61218 597744 61274 597800
rect 61342 597744 61398 597800
rect 60970 586294 61026 586350
rect 61094 586294 61150 586350
rect 61218 586294 61274 586350
rect 61342 586294 61398 586350
rect 60970 586170 61026 586226
rect 61094 586170 61150 586226
rect 61218 586170 61274 586226
rect 61342 586170 61398 586226
rect 60970 586046 61026 586102
rect 61094 586046 61150 586102
rect 61218 586046 61274 586102
rect 61342 586046 61398 586102
rect 60970 585922 61026 585978
rect 61094 585922 61150 585978
rect 61218 585922 61274 585978
rect 61342 585922 61398 585978
rect 60970 568294 61026 568350
rect 61094 568294 61150 568350
rect 61218 568294 61274 568350
rect 61342 568294 61398 568350
rect 60970 568170 61026 568226
rect 61094 568170 61150 568226
rect 61218 568170 61274 568226
rect 61342 568170 61398 568226
rect 60970 568046 61026 568102
rect 61094 568046 61150 568102
rect 61218 568046 61274 568102
rect 61342 568046 61398 568102
rect 60970 567922 61026 567978
rect 61094 567922 61150 567978
rect 61218 567922 61274 567978
rect 61342 567922 61398 567978
rect 60970 550294 61026 550350
rect 61094 550294 61150 550350
rect 61218 550294 61274 550350
rect 61342 550294 61398 550350
rect 60970 550170 61026 550226
rect 61094 550170 61150 550226
rect 61218 550170 61274 550226
rect 61342 550170 61398 550226
rect 60970 550046 61026 550102
rect 61094 550046 61150 550102
rect 61218 550046 61274 550102
rect 61342 550046 61398 550102
rect 60970 549922 61026 549978
rect 61094 549922 61150 549978
rect 61218 549922 61274 549978
rect 61342 549922 61398 549978
rect 60970 532294 61026 532350
rect 61094 532294 61150 532350
rect 61218 532294 61274 532350
rect 61342 532294 61398 532350
rect 60970 532170 61026 532226
rect 61094 532170 61150 532226
rect 61218 532170 61274 532226
rect 61342 532170 61398 532226
rect 60970 532046 61026 532102
rect 61094 532046 61150 532102
rect 61218 532046 61274 532102
rect 61342 532046 61398 532102
rect 60970 531922 61026 531978
rect 61094 531922 61150 531978
rect 61218 531922 61274 531978
rect 61342 531922 61398 531978
rect 60970 514294 61026 514350
rect 61094 514294 61150 514350
rect 61218 514294 61274 514350
rect 61342 514294 61398 514350
rect 60970 514170 61026 514226
rect 61094 514170 61150 514226
rect 61218 514170 61274 514226
rect 61342 514170 61398 514226
rect 60970 514046 61026 514102
rect 61094 514046 61150 514102
rect 61218 514046 61274 514102
rect 61342 514046 61398 514102
rect 60970 513922 61026 513978
rect 61094 513922 61150 513978
rect 61218 513922 61274 513978
rect 61342 513922 61398 513978
rect 60970 496294 61026 496350
rect 61094 496294 61150 496350
rect 61218 496294 61274 496350
rect 61342 496294 61398 496350
rect 60970 496170 61026 496226
rect 61094 496170 61150 496226
rect 61218 496170 61274 496226
rect 61342 496170 61398 496226
rect 60970 496046 61026 496102
rect 61094 496046 61150 496102
rect 61218 496046 61274 496102
rect 61342 496046 61398 496102
rect 60970 495922 61026 495978
rect 61094 495922 61150 495978
rect 61218 495922 61274 495978
rect 61342 495922 61398 495978
rect 60970 478294 61026 478350
rect 61094 478294 61150 478350
rect 61218 478294 61274 478350
rect 61342 478294 61398 478350
rect 60970 478170 61026 478226
rect 61094 478170 61150 478226
rect 61218 478170 61274 478226
rect 61342 478170 61398 478226
rect 60970 478046 61026 478102
rect 61094 478046 61150 478102
rect 61218 478046 61274 478102
rect 61342 478046 61398 478102
rect 60970 477922 61026 477978
rect 61094 477922 61150 477978
rect 61218 477922 61274 477978
rect 61342 477922 61398 477978
rect 60970 460294 61026 460350
rect 61094 460294 61150 460350
rect 61218 460294 61274 460350
rect 61342 460294 61398 460350
rect 60970 460170 61026 460226
rect 61094 460170 61150 460226
rect 61218 460170 61274 460226
rect 61342 460170 61398 460226
rect 60970 460046 61026 460102
rect 61094 460046 61150 460102
rect 61218 460046 61274 460102
rect 61342 460046 61398 460102
rect 60970 459922 61026 459978
rect 61094 459922 61150 459978
rect 61218 459922 61274 459978
rect 61342 459922 61398 459978
rect 60970 442294 61026 442350
rect 61094 442294 61150 442350
rect 61218 442294 61274 442350
rect 61342 442294 61398 442350
rect 60970 442170 61026 442226
rect 61094 442170 61150 442226
rect 61218 442170 61274 442226
rect 61342 442170 61398 442226
rect 60970 442046 61026 442102
rect 61094 442046 61150 442102
rect 61218 442046 61274 442102
rect 61342 442046 61398 442102
rect 60970 441922 61026 441978
rect 61094 441922 61150 441978
rect 61218 441922 61274 441978
rect 61342 441922 61398 441978
rect 60970 424294 61026 424350
rect 61094 424294 61150 424350
rect 61218 424294 61274 424350
rect 61342 424294 61398 424350
rect 60970 424170 61026 424226
rect 61094 424170 61150 424226
rect 61218 424170 61274 424226
rect 61342 424170 61398 424226
rect 60970 424046 61026 424102
rect 61094 424046 61150 424102
rect 61218 424046 61274 424102
rect 61342 424046 61398 424102
rect 60970 423922 61026 423978
rect 61094 423922 61150 423978
rect 61218 423922 61274 423978
rect 61342 423922 61398 423978
rect 60970 406294 61026 406350
rect 61094 406294 61150 406350
rect 61218 406294 61274 406350
rect 61342 406294 61398 406350
rect 60970 406170 61026 406226
rect 61094 406170 61150 406226
rect 61218 406170 61274 406226
rect 61342 406170 61398 406226
rect 60970 406046 61026 406102
rect 61094 406046 61150 406102
rect 61218 406046 61274 406102
rect 61342 406046 61398 406102
rect 60970 405922 61026 405978
rect 61094 405922 61150 405978
rect 61218 405922 61274 405978
rect 61342 405922 61398 405978
rect 60970 388294 61026 388350
rect 61094 388294 61150 388350
rect 61218 388294 61274 388350
rect 61342 388294 61398 388350
rect 60970 388170 61026 388226
rect 61094 388170 61150 388226
rect 61218 388170 61274 388226
rect 61342 388170 61398 388226
rect 60970 388046 61026 388102
rect 61094 388046 61150 388102
rect 61218 388046 61274 388102
rect 61342 388046 61398 388102
rect 60970 387922 61026 387978
rect 61094 387922 61150 387978
rect 61218 387922 61274 387978
rect 61342 387922 61398 387978
rect 60970 370294 61026 370350
rect 61094 370294 61150 370350
rect 61218 370294 61274 370350
rect 61342 370294 61398 370350
rect 60970 370170 61026 370226
rect 61094 370170 61150 370226
rect 61218 370170 61274 370226
rect 61342 370170 61398 370226
rect 60970 370046 61026 370102
rect 61094 370046 61150 370102
rect 61218 370046 61274 370102
rect 61342 370046 61398 370102
rect 60970 369922 61026 369978
rect 61094 369922 61150 369978
rect 61218 369922 61274 369978
rect 61342 369922 61398 369978
rect 60970 352294 61026 352350
rect 61094 352294 61150 352350
rect 61218 352294 61274 352350
rect 61342 352294 61398 352350
rect 60970 352170 61026 352226
rect 61094 352170 61150 352226
rect 61218 352170 61274 352226
rect 61342 352170 61398 352226
rect 60970 352046 61026 352102
rect 61094 352046 61150 352102
rect 61218 352046 61274 352102
rect 61342 352046 61398 352102
rect 60970 351922 61026 351978
rect 61094 351922 61150 351978
rect 61218 351922 61274 351978
rect 61342 351922 61398 351978
rect 60970 334294 61026 334350
rect 61094 334294 61150 334350
rect 61218 334294 61274 334350
rect 61342 334294 61398 334350
rect 60970 334170 61026 334226
rect 61094 334170 61150 334226
rect 61218 334170 61274 334226
rect 61342 334170 61398 334226
rect 60970 334046 61026 334102
rect 61094 334046 61150 334102
rect 61218 334046 61274 334102
rect 61342 334046 61398 334102
rect 60970 333922 61026 333978
rect 61094 333922 61150 333978
rect 61218 333922 61274 333978
rect 61342 333922 61398 333978
rect 60970 316294 61026 316350
rect 61094 316294 61150 316350
rect 61218 316294 61274 316350
rect 61342 316294 61398 316350
rect 60970 316170 61026 316226
rect 61094 316170 61150 316226
rect 61218 316170 61274 316226
rect 61342 316170 61398 316226
rect 60970 316046 61026 316102
rect 61094 316046 61150 316102
rect 61218 316046 61274 316102
rect 61342 316046 61398 316102
rect 60970 315922 61026 315978
rect 61094 315922 61150 315978
rect 61218 315922 61274 315978
rect 61342 315922 61398 315978
rect 60970 298294 61026 298350
rect 61094 298294 61150 298350
rect 61218 298294 61274 298350
rect 61342 298294 61398 298350
rect 60970 298170 61026 298226
rect 61094 298170 61150 298226
rect 61218 298170 61274 298226
rect 61342 298170 61398 298226
rect 60970 298046 61026 298102
rect 61094 298046 61150 298102
rect 61218 298046 61274 298102
rect 61342 298046 61398 298102
rect 60970 297922 61026 297978
rect 61094 297922 61150 297978
rect 61218 297922 61274 297978
rect 61342 297922 61398 297978
rect 60970 280294 61026 280350
rect 61094 280294 61150 280350
rect 61218 280294 61274 280350
rect 61342 280294 61398 280350
rect 60970 280170 61026 280226
rect 61094 280170 61150 280226
rect 61218 280170 61274 280226
rect 61342 280170 61398 280226
rect 60970 280046 61026 280102
rect 61094 280046 61150 280102
rect 61218 280046 61274 280102
rect 61342 280046 61398 280102
rect 60970 279922 61026 279978
rect 61094 279922 61150 279978
rect 61218 279922 61274 279978
rect 61342 279922 61398 279978
rect 60970 262294 61026 262350
rect 61094 262294 61150 262350
rect 61218 262294 61274 262350
rect 61342 262294 61398 262350
rect 60970 262170 61026 262226
rect 61094 262170 61150 262226
rect 61218 262170 61274 262226
rect 61342 262170 61398 262226
rect 60970 262046 61026 262102
rect 61094 262046 61150 262102
rect 61218 262046 61274 262102
rect 61342 262046 61398 262102
rect 60970 261922 61026 261978
rect 61094 261922 61150 261978
rect 61218 261922 61274 261978
rect 61342 261922 61398 261978
rect 60970 244294 61026 244350
rect 61094 244294 61150 244350
rect 61218 244294 61274 244350
rect 61342 244294 61398 244350
rect 60970 244170 61026 244226
rect 61094 244170 61150 244226
rect 61218 244170 61274 244226
rect 61342 244170 61398 244226
rect 60970 244046 61026 244102
rect 61094 244046 61150 244102
rect 61218 244046 61274 244102
rect 61342 244046 61398 244102
rect 60970 243922 61026 243978
rect 61094 243922 61150 243978
rect 61218 243922 61274 243978
rect 61342 243922 61398 243978
rect 60970 226294 61026 226350
rect 61094 226294 61150 226350
rect 61218 226294 61274 226350
rect 61342 226294 61398 226350
rect 60970 226170 61026 226226
rect 61094 226170 61150 226226
rect 61218 226170 61274 226226
rect 61342 226170 61398 226226
rect 60970 226046 61026 226102
rect 61094 226046 61150 226102
rect 61218 226046 61274 226102
rect 61342 226046 61398 226102
rect 60970 225922 61026 225978
rect 61094 225922 61150 225978
rect 61218 225922 61274 225978
rect 61342 225922 61398 225978
rect 60970 208294 61026 208350
rect 61094 208294 61150 208350
rect 61218 208294 61274 208350
rect 61342 208294 61398 208350
rect 60970 208170 61026 208226
rect 61094 208170 61150 208226
rect 61218 208170 61274 208226
rect 61342 208170 61398 208226
rect 60970 208046 61026 208102
rect 61094 208046 61150 208102
rect 61218 208046 61274 208102
rect 61342 208046 61398 208102
rect 60970 207922 61026 207978
rect 61094 207922 61150 207978
rect 61218 207922 61274 207978
rect 61342 207922 61398 207978
rect 60970 190294 61026 190350
rect 61094 190294 61150 190350
rect 61218 190294 61274 190350
rect 61342 190294 61398 190350
rect 60970 190170 61026 190226
rect 61094 190170 61150 190226
rect 61218 190170 61274 190226
rect 61342 190170 61398 190226
rect 60970 190046 61026 190102
rect 61094 190046 61150 190102
rect 61218 190046 61274 190102
rect 61342 190046 61398 190102
rect 60970 189922 61026 189978
rect 61094 189922 61150 189978
rect 61218 189922 61274 189978
rect 61342 189922 61398 189978
rect 60970 172294 61026 172350
rect 61094 172294 61150 172350
rect 61218 172294 61274 172350
rect 61342 172294 61398 172350
rect 60970 172170 61026 172226
rect 61094 172170 61150 172226
rect 61218 172170 61274 172226
rect 61342 172170 61398 172226
rect 60970 172046 61026 172102
rect 61094 172046 61150 172102
rect 61218 172046 61274 172102
rect 61342 172046 61398 172102
rect 60970 171922 61026 171978
rect 61094 171922 61150 171978
rect 61218 171922 61274 171978
rect 61342 171922 61398 171978
rect 60970 154294 61026 154350
rect 61094 154294 61150 154350
rect 61218 154294 61274 154350
rect 61342 154294 61398 154350
rect 60970 154170 61026 154226
rect 61094 154170 61150 154226
rect 61218 154170 61274 154226
rect 61342 154170 61398 154226
rect 60970 154046 61026 154102
rect 61094 154046 61150 154102
rect 61218 154046 61274 154102
rect 61342 154046 61398 154102
rect 60970 153922 61026 153978
rect 61094 153922 61150 153978
rect 61218 153922 61274 153978
rect 61342 153922 61398 153978
rect 60970 136294 61026 136350
rect 61094 136294 61150 136350
rect 61218 136294 61274 136350
rect 61342 136294 61398 136350
rect 60970 136170 61026 136226
rect 61094 136170 61150 136226
rect 61218 136170 61274 136226
rect 61342 136170 61398 136226
rect 60970 136046 61026 136102
rect 61094 136046 61150 136102
rect 61218 136046 61274 136102
rect 61342 136046 61398 136102
rect 60970 135922 61026 135978
rect 61094 135922 61150 135978
rect 61218 135922 61274 135978
rect 61342 135922 61398 135978
rect 60970 118294 61026 118350
rect 61094 118294 61150 118350
rect 61218 118294 61274 118350
rect 61342 118294 61398 118350
rect 60970 118170 61026 118226
rect 61094 118170 61150 118226
rect 61218 118170 61274 118226
rect 61342 118170 61398 118226
rect 60970 118046 61026 118102
rect 61094 118046 61150 118102
rect 61218 118046 61274 118102
rect 61342 118046 61398 118102
rect 60970 117922 61026 117978
rect 61094 117922 61150 117978
rect 61218 117922 61274 117978
rect 61342 117922 61398 117978
rect 60970 100294 61026 100350
rect 61094 100294 61150 100350
rect 61218 100294 61274 100350
rect 61342 100294 61398 100350
rect 60970 100170 61026 100226
rect 61094 100170 61150 100226
rect 61218 100170 61274 100226
rect 61342 100170 61398 100226
rect 60970 100046 61026 100102
rect 61094 100046 61150 100102
rect 61218 100046 61274 100102
rect 61342 100046 61398 100102
rect 60970 99922 61026 99978
rect 61094 99922 61150 99978
rect 61218 99922 61274 99978
rect 61342 99922 61398 99978
rect 60970 82294 61026 82350
rect 61094 82294 61150 82350
rect 61218 82294 61274 82350
rect 61342 82294 61398 82350
rect 60970 82170 61026 82226
rect 61094 82170 61150 82226
rect 61218 82170 61274 82226
rect 61342 82170 61398 82226
rect 60970 82046 61026 82102
rect 61094 82046 61150 82102
rect 61218 82046 61274 82102
rect 61342 82046 61398 82102
rect 60970 81922 61026 81978
rect 61094 81922 61150 81978
rect 61218 81922 61274 81978
rect 61342 81922 61398 81978
rect 60970 64294 61026 64350
rect 61094 64294 61150 64350
rect 61218 64294 61274 64350
rect 61342 64294 61398 64350
rect 60970 64170 61026 64226
rect 61094 64170 61150 64226
rect 61218 64170 61274 64226
rect 61342 64170 61398 64226
rect 60970 64046 61026 64102
rect 61094 64046 61150 64102
rect 61218 64046 61274 64102
rect 61342 64046 61398 64102
rect 60970 63922 61026 63978
rect 61094 63922 61150 63978
rect 61218 63922 61274 63978
rect 61342 63922 61398 63978
rect 60970 46294 61026 46350
rect 61094 46294 61150 46350
rect 61218 46294 61274 46350
rect 61342 46294 61398 46350
rect 60970 46170 61026 46226
rect 61094 46170 61150 46226
rect 61218 46170 61274 46226
rect 61342 46170 61398 46226
rect 60970 46046 61026 46102
rect 61094 46046 61150 46102
rect 61218 46046 61274 46102
rect 61342 46046 61398 46102
rect 60970 45922 61026 45978
rect 61094 45922 61150 45978
rect 61218 45922 61274 45978
rect 61342 45922 61398 45978
rect 60970 28294 61026 28350
rect 61094 28294 61150 28350
rect 61218 28294 61274 28350
rect 61342 28294 61398 28350
rect 60970 28170 61026 28226
rect 61094 28170 61150 28226
rect 61218 28170 61274 28226
rect 61342 28170 61398 28226
rect 60970 28046 61026 28102
rect 61094 28046 61150 28102
rect 61218 28046 61274 28102
rect 61342 28046 61398 28102
rect 60970 27922 61026 27978
rect 61094 27922 61150 27978
rect 61218 27922 61274 27978
rect 61342 27922 61398 27978
rect 60970 10294 61026 10350
rect 61094 10294 61150 10350
rect 61218 10294 61274 10350
rect 61342 10294 61398 10350
rect 60970 10170 61026 10226
rect 61094 10170 61150 10226
rect 61218 10170 61274 10226
rect 61342 10170 61398 10226
rect 60970 10046 61026 10102
rect 61094 10046 61150 10102
rect 61218 10046 61274 10102
rect 61342 10046 61398 10102
rect 60970 9922 61026 9978
rect 61094 9922 61150 9978
rect 61218 9922 61274 9978
rect 61342 9922 61398 9978
rect 60970 -1176 61026 -1120
rect 61094 -1176 61150 -1120
rect 61218 -1176 61274 -1120
rect 61342 -1176 61398 -1120
rect 60970 -1300 61026 -1244
rect 61094 -1300 61150 -1244
rect 61218 -1300 61274 -1244
rect 61342 -1300 61398 -1244
rect 60970 -1424 61026 -1368
rect 61094 -1424 61150 -1368
rect 61218 -1424 61274 -1368
rect 61342 -1424 61398 -1368
rect 60970 -1548 61026 -1492
rect 61094 -1548 61150 -1492
rect 61218 -1548 61274 -1492
rect 61342 -1548 61398 -1492
rect 75250 597156 75306 597212
rect 75374 597156 75430 597212
rect 75498 597156 75554 597212
rect 75622 597156 75678 597212
rect 75250 597032 75306 597088
rect 75374 597032 75430 597088
rect 75498 597032 75554 597088
rect 75622 597032 75678 597088
rect 75250 596908 75306 596964
rect 75374 596908 75430 596964
rect 75498 596908 75554 596964
rect 75622 596908 75678 596964
rect 75250 596784 75306 596840
rect 75374 596784 75430 596840
rect 75498 596784 75554 596840
rect 75622 596784 75678 596840
rect 75250 580294 75306 580350
rect 75374 580294 75430 580350
rect 75498 580294 75554 580350
rect 75622 580294 75678 580350
rect 75250 580170 75306 580226
rect 75374 580170 75430 580226
rect 75498 580170 75554 580226
rect 75622 580170 75678 580226
rect 75250 580046 75306 580102
rect 75374 580046 75430 580102
rect 75498 580046 75554 580102
rect 75622 580046 75678 580102
rect 75250 579922 75306 579978
rect 75374 579922 75430 579978
rect 75498 579922 75554 579978
rect 75622 579922 75678 579978
rect 75250 562294 75306 562350
rect 75374 562294 75430 562350
rect 75498 562294 75554 562350
rect 75622 562294 75678 562350
rect 75250 562170 75306 562226
rect 75374 562170 75430 562226
rect 75498 562170 75554 562226
rect 75622 562170 75678 562226
rect 75250 562046 75306 562102
rect 75374 562046 75430 562102
rect 75498 562046 75554 562102
rect 75622 562046 75678 562102
rect 75250 561922 75306 561978
rect 75374 561922 75430 561978
rect 75498 561922 75554 561978
rect 75622 561922 75678 561978
rect 75250 544294 75306 544350
rect 75374 544294 75430 544350
rect 75498 544294 75554 544350
rect 75622 544294 75678 544350
rect 75250 544170 75306 544226
rect 75374 544170 75430 544226
rect 75498 544170 75554 544226
rect 75622 544170 75678 544226
rect 75250 544046 75306 544102
rect 75374 544046 75430 544102
rect 75498 544046 75554 544102
rect 75622 544046 75678 544102
rect 75250 543922 75306 543978
rect 75374 543922 75430 543978
rect 75498 543922 75554 543978
rect 75622 543922 75678 543978
rect 75250 526294 75306 526350
rect 75374 526294 75430 526350
rect 75498 526294 75554 526350
rect 75622 526294 75678 526350
rect 75250 526170 75306 526226
rect 75374 526170 75430 526226
rect 75498 526170 75554 526226
rect 75622 526170 75678 526226
rect 75250 526046 75306 526102
rect 75374 526046 75430 526102
rect 75498 526046 75554 526102
rect 75622 526046 75678 526102
rect 75250 525922 75306 525978
rect 75374 525922 75430 525978
rect 75498 525922 75554 525978
rect 75622 525922 75678 525978
rect 75250 508294 75306 508350
rect 75374 508294 75430 508350
rect 75498 508294 75554 508350
rect 75622 508294 75678 508350
rect 75250 508170 75306 508226
rect 75374 508170 75430 508226
rect 75498 508170 75554 508226
rect 75622 508170 75678 508226
rect 75250 508046 75306 508102
rect 75374 508046 75430 508102
rect 75498 508046 75554 508102
rect 75622 508046 75678 508102
rect 75250 507922 75306 507978
rect 75374 507922 75430 507978
rect 75498 507922 75554 507978
rect 75622 507922 75678 507978
rect 75250 490294 75306 490350
rect 75374 490294 75430 490350
rect 75498 490294 75554 490350
rect 75622 490294 75678 490350
rect 75250 490170 75306 490226
rect 75374 490170 75430 490226
rect 75498 490170 75554 490226
rect 75622 490170 75678 490226
rect 75250 490046 75306 490102
rect 75374 490046 75430 490102
rect 75498 490046 75554 490102
rect 75622 490046 75678 490102
rect 75250 489922 75306 489978
rect 75374 489922 75430 489978
rect 75498 489922 75554 489978
rect 75622 489922 75678 489978
rect 75250 472294 75306 472350
rect 75374 472294 75430 472350
rect 75498 472294 75554 472350
rect 75622 472294 75678 472350
rect 75250 472170 75306 472226
rect 75374 472170 75430 472226
rect 75498 472170 75554 472226
rect 75622 472170 75678 472226
rect 75250 472046 75306 472102
rect 75374 472046 75430 472102
rect 75498 472046 75554 472102
rect 75622 472046 75678 472102
rect 75250 471922 75306 471978
rect 75374 471922 75430 471978
rect 75498 471922 75554 471978
rect 75622 471922 75678 471978
rect 75250 454294 75306 454350
rect 75374 454294 75430 454350
rect 75498 454294 75554 454350
rect 75622 454294 75678 454350
rect 75250 454170 75306 454226
rect 75374 454170 75430 454226
rect 75498 454170 75554 454226
rect 75622 454170 75678 454226
rect 75250 454046 75306 454102
rect 75374 454046 75430 454102
rect 75498 454046 75554 454102
rect 75622 454046 75678 454102
rect 75250 453922 75306 453978
rect 75374 453922 75430 453978
rect 75498 453922 75554 453978
rect 75622 453922 75678 453978
rect 75250 436294 75306 436350
rect 75374 436294 75430 436350
rect 75498 436294 75554 436350
rect 75622 436294 75678 436350
rect 75250 436170 75306 436226
rect 75374 436170 75430 436226
rect 75498 436170 75554 436226
rect 75622 436170 75678 436226
rect 75250 436046 75306 436102
rect 75374 436046 75430 436102
rect 75498 436046 75554 436102
rect 75622 436046 75678 436102
rect 75250 435922 75306 435978
rect 75374 435922 75430 435978
rect 75498 435922 75554 435978
rect 75622 435922 75678 435978
rect 75250 418294 75306 418350
rect 75374 418294 75430 418350
rect 75498 418294 75554 418350
rect 75622 418294 75678 418350
rect 75250 418170 75306 418226
rect 75374 418170 75430 418226
rect 75498 418170 75554 418226
rect 75622 418170 75678 418226
rect 75250 418046 75306 418102
rect 75374 418046 75430 418102
rect 75498 418046 75554 418102
rect 75622 418046 75678 418102
rect 75250 417922 75306 417978
rect 75374 417922 75430 417978
rect 75498 417922 75554 417978
rect 75622 417922 75678 417978
rect 75250 400294 75306 400350
rect 75374 400294 75430 400350
rect 75498 400294 75554 400350
rect 75622 400294 75678 400350
rect 75250 400170 75306 400226
rect 75374 400170 75430 400226
rect 75498 400170 75554 400226
rect 75622 400170 75678 400226
rect 75250 400046 75306 400102
rect 75374 400046 75430 400102
rect 75498 400046 75554 400102
rect 75622 400046 75678 400102
rect 75250 399922 75306 399978
rect 75374 399922 75430 399978
rect 75498 399922 75554 399978
rect 75622 399922 75678 399978
rect 75250 382294 75306 382350
rect 75374 382294 75430 382350
rect 75498 382294 75554 382350
rect 75622 382294 75678 382350
rect 75250 382170 75306 382226
rect 75374 382170 75430 382226
rect 75498 382170 75554 382226
rect 75622 382170 75678 382226
rect 75250 382046 75306 382102
rect 75374 382046 75430 382102
rect 75498 382046 75554 382102
rect 75622 382046 75678 382102
rect 75250 381922 75306 381978
rect 75374 381922 75430 381978
rect 75498 381922 75554 381978
rect 75622 381922 75678 381978
rect 75250 364294 75306 364350
rect 75374 364294 75430 364350
rect 75498 364294 75554 364350
rect 75622 364294 75678 364350
rect 75250 364170 75306 364226
rect 75374 364170 75430 364226
rect 75498 364170 75554 364226
rect 75622 364170 75678 364226
rect 75250 364046 75306 364102
rect 75374 364046 75430 364102
rect 75498 364046 75554 364102
rect 75622 364046 75678 364102
rect 75250 363922 75306 363978
rect 75374 363922 75430 363978
rect 75498 363922 75554 363978
rect 75622 363922 75678 363978
rect 75250 346294 75306 346350
rect 75374 346294 75430 346350
rect 75498 346294 75554 346350
rect 75622 346294 75678 346350
rect 75250 346170 75306 346226
rect 75374 346170 75430 346226
rect 75498 346170 75554 346226
rect 75622 346170 75678 346226
rect 75250 346046 75306 346102
rect 75374 346046 75430 346102
rect 75498 346046 75554 346102
rect 75622 346046 75678 346102
rect 75250 345922 75306 345978
rect 75374 345922 75430 345978
rect 75498 345922 75554 345978
rect 75622 345922 75678 345978
rect 75250 328294 75306 328350
rect 75374 328294 75430 328350
rect 75498 328294 75554 328350
rect 75622 328294 75678 328350
rect 75250 328170 75306 328226
rect 75374 328170 75430 328226
rect 75498 328170 75554 328226
rect 75622 328170 75678 328226
rect 75250 328046 75306 328102
rect 75374 328046 75430 328102
rect 75498 328046 75554 328102
rect 75622 328046 75678 328102
rect 75250 327922 75306 327978
rect 75374 327922 75430 327978
rect 75498 327922 75554 327978
rect 75622 327922 75678 327978
rect 75250 310294 75306 310350
rect 75374 310294 75430 310350
rect 75498 310294 75554 310350
rect 75622 310294 75678 310350
rect 75250 310170 75306 310226
rect 75374 310170 75430 310226
rect 75498 310170 75554 310226
rect 75622 310170 75678 310226
rect 75250 310046 75306 310102
rect 75374 310046 75430 310102
rect 75498 310046 75554 310102
rect 75622 310046 75678 310102
rect 75250 309922 75306 309978
rect 75374 309922 75430 309978
rect 75498 309922 75554 309978
rect 75622 309922 75678 309978
rect 75250 292294 75306 292350
rect 75374 292294 75430 292350
rect 75498 292294 75554 292350
rect 75622 292294 75678 292350
rect 75250 292170 75306 292226
rect 75374 292170 75430 292226
rect 75498 292170 75554 292226
rect 75622 292170 75678 292226
rect 75250 292046 75306 292102
rect 75374 292046 75430 292102
rect 75498 292046 75554 292102
rect 75622 292046 75678 292102
rect 75250 291922 75306 291978
rect 75374 291922 75430 291978
rect 75498 291922 75554 291978
rect 75622 291922 75678 291978
rect 75250 274294 75306 274350
rect 75374 274294 75430 274350
rect 75498 274294 75554 274350
rect 75622 274294 75678 274350
rect 75250 274170 75306 274226
rect 75374 274170 75430 274226
rect 75498 274170 75554 274226
rect 75622 274170 75678 274226
rect 75250 274046 75306 274102
rect 75374 274046 75430 274102
rect 75498 274046 75554 274102
rect 75622 274046 75678 274102
rect 75250 273922 75306 273978
rect 75374 273922 75430 273978
rect 75498 273922 75554 273978
rect 75622 273922 75678 273978
rect 75250 256294 75306 256350
rect 75374 256294 75430 256350
rect 75498 256294 75554 256350
rect 75622 256294 75678 256350
rect 75250 256170 75306 256226
rect 75374 256170 75430 256226
rect 75498 256170 75554 256226
rect 75622 256170 75678 256226
rect 75250 256046 75306 256102
rect 75374 256046 75430 256102
rect 75498 256046 75554 256102
rect 75622 256046 75678 256102
rect 75250 255922 75306 255978
rect 75374 255922 75430 255978
rect 75498 255922 75554 255978
rect 75622 255922 75678 255978
rect 75250 238294 75306 238350
rect 75374 238294 75430 238350
rect 75498 238294 75554 238350
rect 75622 238294 75678 238350
rect 75250 238170 75306 238226
rect 75374 238170 75430 238226
rect 75498 238170 75554 238226
rect 75622 238170 75678 238226
rect 75250 238046 75306 238102
rect 75374 238046 75430 238102
rect 75498 238046 75554 238102
rect 75622 238046 75678 238102
rect 75250 237922 75306 237978
rect 75374 237922 75430 237978
rect 75498 237922 75554 237978
rect 75622 237922 75678 237978
rect 75250 220294 75306 220350
rect 75374 220294 75430 220350
rect 75498 220294 75554 220350
rect 75622 220294 75678 220350
rect 75250 220170 75306 220226
rect 75374 220170 75430 220226
rect 75498 220170 75554 220226
rect 75622 220170 75678 220226
rect 75250 220046 75306 220102
rect 75374 220046 75430 220102
rect 75498 220046 75554 220102
rect 75622 220046 75678 220102
rect 75250 219922 75306 219978
rect 75374 219922 75430 219978
rect 75498 219922 75554 219978
rect 75622 219922 75678 219978
rect 75250 202294 75306 202350
rect 75374 202294 75430 202350
rect 75498 202294 75554 202350
rect 75622 202294 75678 202350
rect 75250 202170 75306 202226
rect 75374 202170 75430 202226
rect 75498 202170 75554 202226
rect 75622 202170 75678 202226
rect 75250 202046 75306 202102
rect 75374 202046 75430 202102
rect 75498 202046 75554 202102
rect 75622 202046 75678 202102
rect 75250 201922 75306 201978
rect 75374 201922 75430 201978
rect 75498 201922 75554 201978
rect 75622 201922 75678 201978
rect 75250 184294 75306 184350
rect 75374 184294 75430 184350
rect 75498 184294 75554 184350
rect 75622 184294 75678 184350
rect 75250 184170 75306 184226
rect 75374 184170 75430 184226
rect 75498 184170 75554 184226
rect 75622 184170 75678 184226
rect 75250 184046 75306 184102
rect 75374 184046 75430 184102
rect 75498 184046 75554 184102
rect 75622 184046 75678 184102
rect 75250 183922 75306 183978
rect 75374 183922 75430 183978
rect 75498 183922 75554 183978
rect 75622 183922 75678 183978
rect 75250 166294 75306 166350
rect 75374 166294 75430 166350
rect 75498 166294 75554 166350
rect 75622 166294 75678 166350
rect 75250 166170 75306 166226
rect 75374 166170 75430 166226
rect 75498 166170 75554 166226
rect 75622 166170 75678 166226
rect 75250 166046 75306 166102
rect 75374 166046 75430 166102
rect 75498 166046 75554 166102
rect 75622 166046 75678 166102
rect 75250 165922 75306 165978
rect 75374 165922 75430 165978
rect 75498 165922 75554 165978
rect 75622 165922 75678 165978
rect 75250 148294 75306 148350
rect 75374 148294 75430 148350
rect 75498 148294 75554 148350
rect 75622 148294 75678 148350
rect 75250 148170 75306 148226
rect 75374 148170 75430 148226
rect 75498 148170 75554 148226
rect 75622 148170 75678 148226
rect 75250 148046 75306 148102
rect 75374 148046 75430 148102
rect 75498 148046 75554 148102
rect 75622 148046 75678 148102
rect 75250 147922 75306 147978
rect 75374 147922 75430 147978
rect 75498 147922 75554 147978
rect 75622 147922 75678 147978
rect 75250 130294 75306 130350
rect 75374 130294 75430 130350
rect 75498 130294 75554 130350
rect 75622 130294 75678 130350
rect 75250 130170 75306 130226
rect 75374 130170 75430 130226
rect 75498 130170 75554 130226
rect 75622 130170 75678 130226
rect 75250 130046 75306 130102
rect 75374 130046 75430 130102
rect 75498 130046 75554 130102
rect 75622 130046 75678 130102
rect 75250 129922 75306 129978
rect 75374 129922 75430 129978
rect 75498 129922 75554 129978
rect 75622 129922 75678 129978
rect 75250 112294 75306 112350
rect 75374 112294 75430 112350
rect 75498 112294 75554 112350
rect 75622 112294 75678 112350
rect 75250 112170 75306 112226
rect 75374 112170 75430 112226
rect 75498 112170 75554 112226
rect 75622 112170 75678 112226
rect 75250 112046 75306 112102
rect 75374 112046 75430 112102
rect 75498 112046 75554 112102
rect 75622 112046 75678 112102
rect 75250 111922 75306 111978
rect 75374 111922 75430 111978
rect 75498 111922 75554 111978
rect 75622 111922 75678 111978
rect 75250 94294 75306 94350
rect 75374 94294 75430 94350
rect 75498 94294 75554 94350
rect 75622 94294 75678 94350
rect 75250 94170 75306 94226
rect 75374 94170 75430 94226
rect 75498 94170 75554 94226
rect 75622 94170 75678 94226
rect 75250 94046 75306 94102
rect 75374 94046 75430 94102
rect 75498 94046 75554 94102
rect 75622 94046 75678 94102
rect 75250 93922 75306 93978
rect 75374 93922 75430 93978
rect 75498 93922 75554 93978
rect 75622 93922 75678 93978
rect 75250 76294 75306 76350
rect 75374 76294 75430 76350
rect 75498 76294 75554 76350
rect 75622 76294 75678 76350
rect 75250 76170 75306 76226
rect 75374 76170 75430 76226
rect 75498 76170 75554 76226
rect 75622 76170 75678 76226
rect 75250 76046 75306 76102
rect 75374 76046 75430 76102
rect 75498 76046 75554 76102
rect 75622 76046 75678 76102
rect 75250 75922 75306 75978
rect 75374 75922 75430 75978
rect 75498 75922 75554 75978
rect 75622 75922 75678 75978
rect 75250 58294 75306 58350
rect 75374 58294 75430 58350
rect 75498 58294 75554 58350
rect 75622 58294 75678 58350
rect 75250 58170 75306 58226
rect 75374 58170 75430 58226
rect 75498 58170 75554 58226
rect 75622 58170 75678 58226
rect 75250 58046 75306 58102
rect 75374 58046 75430 58102
rect 75498 58046 75554 58102
rect 75622 58046 75678 58102
rect 75250 57922 75306 57978
rect 75374 57922 75430 57978
rect 75498 57922 75554 57978
rect 75622 57922 75678 57978
rect 75250 40294 75306 40350
rect 75374 40294 75430 40350
rect 75498 40294 75554 40350
rect 75622 40294 75678 40350
rect 75250 40170 75306 40226
rect 75374 40170 75430 40226
rect 75498 40170 75554 40226
rect 75622 40170 75678 40226
rect 75250 40046 75306 40102
rect 75374 40046 75430 40102
rect 75498 40046 75554 40102
rect 75622 40046 75678 40102
rect 75250 39922 75306 39978
rect 75374 39922 75430 39978
rect 75498 39922 75554 39978
rect 75622 39922 75678 39978
rect 75250 22294 75306 22350
rect 75374 22294 75430 22350
rect 75498 22294 75554 22350
rect 75622 22294 75678 22350
rect 75250 22170 75306 22226
rect 75374 22170 75430 22226
rect 75498 22170 75554 22226
rect 75622 22170 75678 22226
rect 75250 22046 75306 22102
rect 75374 22046 75430 22102
rect 75498 22046 75554 22102
rect 75622 22046 75678 22102
rect 75250 21922 75306 21978
rect 75374 21922 75430 21978
rect 75498 21922 75554 21978
rect 75622 21922 75678 21978
rect 75250 4294 75306 4350
rect 75374 4294 75430 4350
rect 75498 4294 75554 4350
rect 75622 4294 75678 4350
rect 75250 4170 75306 4226
rect 75374 4170 75430 4226
rect 75498 4170 75554 4226
rect 75622 4170 75678 4226
rect 75250 4046 75306 4102
rect 75374 4046 75430 4102
rect 75498 4046 75554 4102
rect 75622 4046 75678 4102
rect 75250 3922 75306 3978
rect 75374 3922 75430 3978
rect 75498 3922 75554 3978
rect 75622 3922 75678 3978
rect 75250 -216 75306 -160
rect 75374 -216 75430 -160
rect 75498 -216 75554 -160
rect 75622 -216 75678 -160
rect 75250 -340 75306 -284
rect 75374 -340 75430 -284
rect 75498 -340 75554 -284
rect 75622 -340 75678 -284
rect 75250 -464 75306 -408
rect 75374 -464 75430 -408
rect 75498 -464 75554 -408
rect 75622 -464 75678 -408
rect 75250 -588 75306 -532
rect 75374 -588 75430 -532
rect 75498 -588 75554 -532
rect 75622 -588 75678 -532
rect 78970 598116 79026 598172
rect 79094 598116 79150 598172
rect 79218 598116 79274 598172
rect 79342 598116 79398 598172
rect 78970 597992 79026 598048
rect 79094 597992 79150 598048
rect 79218 597992 79274 598048
rect 79342 597992 79398 598048
rect 78970 597868 79026 597924
rect 79094 597868 79150 597924
rect 79218 597868 79274 597924
rect 79342 597868 79398 597924
rect 78970 597744 79026 597800
rect 79094 597744 79150 597800
rect 79218 597744 79274 597800
rect 79342 597744 79398 597800
rect 78970 586294 79026 586350
rect 79094 586294 79150 586350
rect 79218 586294 79274 586350
rect 79342 586294 79398 586350
rect 78970 586170 79026 586226
rect 79094 586170 79150 586226
rect 79218 586170 79274 586226
rect 79342 586170 79398 586226
rect 78970 586046 79026 586102
rect 79094 586046 79150 586102
rect 79218 586046 79274 586102
rect 79342 586046 79398 586102
rect 78970 585922 79026 585978
rect 79094 585922 79150 585978
rect 79218 585922 79274 585978
rect 79342 585922 79398 585978
rect 78970 568294 79026 568350
rect 79094 568294 79150 568350
rect 79218 568294 79274 568350
rect 79342 568294 79398 568350
rect 78970 568170 79026 568226
rect 79094 568170 79150 568226
rect 79218 568170 79274 568226
rect 79342 568170 79398 568226
rect 78970 568046 79026 568102
rect 79094 568046 79150 568102
rect 79218 568046 79274 568102
rect 79342 568046 79398 568102
rect 78970 567922 79026 567978
rect 79094 567922 79150 567978
rect 79218 567922 79274 567978
rect 79342 567922 79398 567978
rect 78970 550294 79026 550350
rect 79094 550294 79150 550350
rect 79218 550294 79274 550350
rect 79342 550294 79398 550350
rect 78970 550170 79026 550226
rect 79094 550170 79150 550226
rect 79218 550170 79274 550226
rect 79342 550170 79398 550226
rect 78970 550046 79026 550102
rect 79094 550046 79150 550102
rect 79218 550046 79274 550102
rect 79342 550046 79398 550102
rect 78970 549922 79026 549978
rect 79094 549922 79150 549978
rect 79218 549922 79274 549978
rect 79342 549922 79398 549978
rect 78970 532294 79026 532350
rect 79094 532294 79150 532350
rect 79218 532294 79274 532350
rect 79342 532294 79398 532350
rect 78970 532170 79026 532226
rect 79094 532170 79150 532226
rect 79218 532170 79274 532226
rect 79342 532170 79398 532226
rect 78970 532046 79026 532102
rect 79094 532046 79150 532102
rect 79218 532046 79274 532102
rect 79342 532046 79398 532102
rect 78970 531922 79026 531978
rect 79094 531922 79150 531978
rect 79218 531922 79274 531978
rect 79342 531922 79398 531978
rect 78970 514294 79026 514350
rect 79094 514294 79150 514350
rect 79218 514294 79274 514350
rect 79342 514294 79398 514350
rect 78970 514170 79026 514226
rect 79094 514170 79150 514226
rect 79218 514170 79274 514226
rect 79342 514170 79398 514226
rect 78970 514046 79026 514102
rect 79094 514046 79150 514102
rect 79218 514046 79274 514102
rect 79342 514046 79398 514102
rect 78970 513922 79026 513978
rect 79094 513922 79150 513978
rect 79218 513922 79274 513978
rect 79342 513922 79398 513978
rect 78970 496294 79026 496350
rect 79094 496294 79150 496350
rect 79218 496294 79274 496350
rect 79342 496294 79398 496350
rect 78970 496170 79026 496226
rect 79094 496170 79150 496226
rect 79218 496170 79274 496226
rect 79342 496170 79398 496226
rect 78970 496046 79026 496102
rect 79094 496046 79150 496102
rect 79218 496046 79274 496102
rect 79342 496046 79398 496102
rect 78970 495922 79026 495978
rect 79094 495922 79150 495978
rect 79218 495922 79274 495978
rect 79342 495922 79398 495978
rect 78970 478294 79026 478350
rect 79094 478294 79150 478350
rect 79218 478294 79274 478350
rect 79342 478294 79398 478350
rect 78970 478170 79026 478226
rect 79094 478170 79150 478226
rect 79218 478170 79274 478226
rect 79342 478170 79398 478226
rect 78970 478046 79026 478102
rect 79094 478046 79150 478102
rect 79218 478046 79274 478102
rect 79342 478046 79398 478102
rect 78970 477922 79026 477978
rect 79094 477922 79150 477978
rect 79218 477922 79274 477978
rect 79342 477922 79398 477978
rect 78970 460294 79026 460350
rect 79094 460294 79150 460350
rect 79218 460294 79274 460350
rect 79342 460294 79398 460350
rect 78970 460170 79026 460226
rect 79094 460170 79150 460226
rect 79218 460170 79274 460226
rect 79342 460170 79398 460226
rect 78970 460046 79026 460102
rect 79094 460046 79150 460102
rect 79218 460046 79274 460102
rect 79342 460046 79398 460102
rect 78970 459922 79026 459978
rect 79094 459922 79150 459978
rect 79218 459922 79274 459978
rect 79342 459922 79398 459978
rect 78970 442294 79026 442350
rect 79094 442294 79150 442350
rect 79218 442294 79274 442350
rect 79342 442294 79398 442350
rect 78970 442170 79026 442226
rect 79094 442170 79150 442226
rect 79218 442170 79274 442226
rect 79342 442170 79398 442226
rect 78970 442046 79026 442102
rect 79094 442046 79150 442102
rect 79218 442046 79274 442102
rect 79342 442046 79398 442102
rect 78970 441922 79026 441978
rect 79094 441922 79150 441978
rect 79218 441922 79274 441978
rect 79342 441922 79398 441978
rect 78970 424294 79026 424350
rect 79094 424294 79150 424350
rect 79218 424294 79274 424350
rect 79342 424294 79398 424350
rect 78970 424170 79026 424226
rect 79094 424170 79150 424226
rect 79218 424170 79274 424226
rect 79342 424170 79398 424226
rect 78970 424046 79026 424102
rect 79094 424046 79150 424102
rect 79218 424046 79274 424102
rect 79342 424046 79398 424102
rect 78970 423922 79026 423978
rect 79094 423922 79150 423978
rect 79218 423922 79274 423978
rect 79342 423922 79398 423978
rect 78970 406294 79026 406350
rect 79094 406294 79150 406350
rect 79218 406294 79274 406350
rect 79342 406294 79398 406350
rect 78970 406170 79026 406226
rect 79094 406170 79150 406226
rect 79218 406170 79274 406226
rect 79342 406170 79398 406226
rect 78970 406046 79026 406102
rect 79094 406046 79150 406102
rect 79218 406046 79274 406102
rect 79342 406046 79398 406102
rect 78970 405922 79026 405978
rect 79094 405922 79150 405978
rect 79218 405922 79274 405978
rect 79342 405922 79398 405978
rect 78970 388294 79026 388350
rect 79094 388294 79150 388350
rect 79218 388294 79274 388350
rect 79342 388294 79398 388350
rect 78970 388170 79026 388226
rect 79094 388170 79150 388226
rect 79218 388170 79274 388226
rect 79342 388170 79398 388226
rect 78970 388046 79026 388102
rect 79094 388046 79150 388102
rect 79218 388046 79274 388102
rect 79342 388046 79398 388102
rect 78970 387922 79026 387978
rect 79094 387922 79150 387978
rect 79218 387922 79274 387978
rect 79342 387922 79398 387978
rect 78970 370294 79026 370350
rect 79094 370294 79150 370350
rect 79218 370294 79274 370350
rect 79342 370294 79398 370350
rect 78970 370170 79026 370226
rect 79094 370170 79150 370226
rect 79218 370170 79274 370226
rect 79342 370170 79398 370226
rect 78970 370046 79026 370102
rect 79094 370046 79150 370102
rect 79218 370046 79274 370102
rect 79342 370046 79398 370102
rect 78970 369922 79026 369978
rect 79094 369922 79150 369978
rect 79218 369922 79274 369978
rect 79342 369922 79398 369978
rect 78970 352294 79026 352350
rect 79094 352294 79150 352350
rect 79218 352294 79274 352350
rect 79342 352294 79398 352350
rect 78970 352170 79026 352226
rect 79094 352170 79150 352226
rect 79218 352170 79274 352226
rect 79342 352170 79398 352226
rect 78970 352046 79026 352102
rect 79094 352046 79150 352102
rect 79218 352046 79274 352102
rect 79342 352046 79398 352102
rect 78970 351922 79026 351978
rect 79094 351922 79150 351978
rect 79218 351922 79274 351978
rect 79342 351922 79398 351978
rect 78970 334294 79026 334350
rect 79094 334294 79150 334350
rect 79218 334294 79274 334350
rect 79342 334294 79398 334350
rect 78970 334170 79026 334226
rect 79094 334170 79150 334226
rect 79218 334170 79274 334226
rect 79342 334170 79398 334226
rect 78970 334046 79026 334102
rect 79094 334046 79150 334102
rect 79218 334046 79274 334102
rect 79342 334046 79398 334102
rect 78970 333922 79026 333978
rect 79094 333922 79150 333978
rect 79218 333922 79274 333978
rect 79342 333922 79398 333978
rect 78970 316294 79026 316350
rect 79094 316294 79150 316350
rect 79218 316294 79274 316350
rect 79342 316294 79398 316350
rect 78970 316170 79026 316226
rect 79094 316170 79150 316226
rect 79218 316170 79274 316226
rect 79342 316170 79398 316226
rect 78970 316046 79026 316102
rect 79094 316046 79150 316102
rect 79218 316046 79274 316102
rect 79342 316046 79398 316102
rect 78970 315922 79026 315978
rect 79094 315922 79150 315978
rect 79218 315922 79274 315978
rect 79342 315922 79398 315978
rect 78970 298294 79026 298350
rect 79094 298294 79150 298350
rect 79218 298294 79274 298350
rect 79342 298294 79398 298350
rect 78970 298170 79026 298226
rect 79094 298170 79150 298226
rect 79218 298170 79274 298226
rect 79342 298170 79398 298226
rect 78970 298046 79026 298102
rect 79094 298046 79150 298102
rect 79218 298046 79274 298102
rect 79342 298046 79398 298102
rect 78970 297922 79026 297978
rect 79094 297922 79150 297978
rect 79218 297922 79274 297978
rect 79342 297922 79398 297978
rect 78970 280294 79026 280350
rect 79094 280294 79150 280350
rect 79218 280294 79274 280350
rect 79342 280294 79398 280350
rect 78970 280170 79026 280226
rect 79094 280170 79150 280226
rect 79218 280170 79274 280226
rect 79342 280170 79398 280226
rect 78970 280046 79026 280102
rect 79094 280046 79150 280102
rect 79218 280046 79274 280102
rect 79342 280046 79398 280102
rect 78970 279922 79026 279978
rect 79094 279922 79150 279978
rect 79218 279922 79274 279978
rect 79342 279922 79398 279978
rect 78970 262294 79026 262350
rect 79094 262294 79150 262350
rect 79218 262294 79274 262350
rect 79342 262294 79398 262350
rect 78970 262170 79026 262226
rect 79094 262170 79150 262226
rect 79218 262170 79274 262226
rect 79342 262170 79398 262226
rect 78970 262046 79026 262102
rect 79094 262046 79150 262102
rect 79218 262046 79274 262102
rect 79342 262046 79398 262102
rect 78970 261922 79026 261978
rect 79094 261922 79150 261978
rect 79218 261922 79274 261978
rect 79342 261922 79398 261978
rect 78970 244294 79026 244350
rect 79094 244294 79150 244350
rect 79218 244294 79274 244350
rect 79342 244294 79398 244350
rect 78970 244170 79026 244226
rect 79094 244170 79150 244226
rect 79218 244170 79274 244226
rect 79342 244170 79398 244226
rect 78970 244046 79026 244102
rect 79094 244046 79150 244102
rect 79218 244046 79274 244102
rect 79342 244046 79398 244102
rect 78970 243922 79026 243978
rect 79094 243922 79150 243978
rect 79218 243922 79274 243978
rect 79342 243922 79398 243978
rect 78970 226294 79026 226350
rect 79094 226294 79150 226350
rect 79218 226294 79274 226350
rect 79342 226294 79398 226350
rect 78970 226170 79026 226226
rect 79094 226170 79150 226226
rect 79218 226170 79274 226226
rect 79342 226170 79398 226226
rect 78970 226046 79026 226102
rect 79094 226046 79150 226102
rect 79218 226046 79274 226102
rect 79342 226046 79398 226102
rect 78970 225922 79026 225978
rect 79094 225922 79150 225978
rect 79218 225922 79274 225978
rect 79342 225922 79398 225978
rect 78970 208294 79026 208350
rect 79094 208294 79150 208350
rect 79218 208294 79274 208350
rect 79342 208294 79398 208350
rect 78970 208170 79026 208226
rect 79094 208170 79150 208226
rect 79218 208170 79274 208226
rect 79342 208170 79398 208226
rect 78970 208046 79026 208102
rect 79094 208046 79150 208102
rect 79218 208046 79274 208102
rect 79342 208046 79398 208102
rect 78970 207922 79026 207978
rect 79094 207922 79150 207978
rect 79218 207922 79274 207978
rect 79342 207922 79398 207978
rect 78970 190294 79026 190350
rect 79094 190294 79150 190350
rect 79218 190294 79274 190350
rect 79342 190294 79398 190350
rect 78970 190170 79026 190226
rect 79094 190170 79150 190226
rect 79218 190170 79274 190226
rect 79342 190170 79398 190226
rect 78970 190046 79026 190102
rect 79094 190046 79150 190102
rect 79218 190046 79274 190102
rect 79342 190046 79398 190102
rect 78970 189922 79026 189978
rect 79094 189922 79150 189978
rect 79218 189922 79274 189978
rect 79342 189922 79398 189978
rect 78970 172294 79026 172350
rect 79094 172294 79150 172350
rect 79218 172294 79274 172350
rect 79342 172294 79398 172350
rect 78970 172170 79026 172226
rect 79094 172170 79150 172226
rect 79218 172170 79274 172226
rect 79342 172170 79398 172226
rect 78970 172046 79026 172102
rect 79094 172046 79150 172102
rect 79218 172046 79274 172102
rect 79342 172046 79398 172102
rect 78970 171922 79026 171978
rect 79094 171922 79150 171978
rect 79218 171922 79274 171978
rect 79342 171922 79398 171978
rect 78970 154294 79026 154350
rect 79094 154294 79150 154350
rect 79218 154294 79274 154350
rect 79342 154294 79398 154350
rect 78970 154170 79026 154226
rect 79094 154170 79150 154226
rect 79218 154170 79274 154226
rect 79342 154170 79398 154226
rect 78970 154046 79026 154102
rect 79094 154046 79150 154102
rect 79218 154046 79274 154102
rect 79342 154046 79398 154102
rect 78970 153922 79026 153978
rect 79094 153922 79150 153978
rect 79218 153922 79274 153978
rect 79342 153922 79398 153978
rect 78970 136294 79026 136350
rect 79094 136294 79150 136350
rect 79218 136294 79274 136350
rect 79342 136294 79398 136350
rect 78970 136170 79026 136226
rect 79094 136170 79150 136226
rect 79218 136170 79274 136226
rect 79342 136170 79398 136226
rect 78970 136046 79026 136102
rect 79094 136046 79150 136102
rect 79218 136046 79274 136102
rect 79342 136046 79398 136102
rect 78970 135922 79026 135978
rect 79094 135922 79150 135978
rect 79218 135922 79274 135978
rect 79342 135922 79398 135978
rect 78970 118294 79026 118350
rect 79094 118294 79150 118350
rect 79218 118294 79274 118350
rect 79342 118294 79398 118350
rect 78970 118170 79026 118226
rect 79094 118170 79150 118226
rect 79218 118170 79274 118226
rect 79342 118170 79398 118226
rect 78970 118046 79026 118102
rect 79094 118046 79150 118102
rect 79218 118046 79274 118102
rect 79342 118046 79398 118102
rect 78970 117922 79026 117978
rect 79094 117922 79150 117978
rect 79218 117922 79274 117978
rect 79342 117922 79398 117978
rect 78970 100294 79026 100350
rect 79094 100294 79150 100350
rect 79218 100294 79274 100350
rect 79342 100294 79398 100350
rect 78970 100170 79026 100226
rect 79094 100170 79150 100226
rect 79218 100170 79274 100226
rect 79342 100170 79398 100226
rect 78970 100046 79026 100102
rect 79094 100046 79150 100102
rect 79218 100046 79274 100102
rect 79342 100046 79398 100102
rect 78970 99922 79026 99978
rect 79094 99922 79150 99978
rect 79218 99922 79274 99978
rect 79342 99922 79398 99978
rect 78970 82294 79026 82350
rect 79094 82294 79150 82350
rect 79218 82294 79274 82350
rect 79342 82294 79398 82350
rect 78970 82170 79026 82226
rect 79094 82170 79150 82226
rect 79218 82170 79274 82226
rect 79342 82170 79398 82226
rect 78970 82046 79026 82102
rect 79094 82046 79150 82102
rect 79218 82046 79274 82102
rect 79342 82046 79398 82102
rect 78970 81922 79026 81978
rect 79094 81922 79150 81978
rect 79218 81922 79274 81978
rect 79342 81922 79398 81978
rect 78970 64294 79026 64350
rect 79094 64294 79150 64350
rect 79218 64294 79274 64350
rect 79342 64294 79398 64350
rect 78970 64170 79026 64226
rect 79094 64170 79150 64226
rect 79218 64170 79274 64226
rect 79342 64170 79398 64226
rect 78970 64046 79026 64102
rect 79094 64046 79150 64102
rect 79218 64046 79274 64102
rect 79342 64046 79398 64102
rect 78970 63922 79026 63978
rect 79094 63922 79150 63978
rect 79218 63922 79274 63978
rect 79342 63922 79398 63978
rect 78970 46294 79026 46350
rect 79094 46294 79150 46350
rect 79218 46294 79274 46350
rect 79342 46294 79398 46350
rect 78970 46170 79026 46226
rect 79094 46170 79150 46226
rect 79218 46170 79274 46226
rect 79342 46170 79398 46226
rect 78970 46046 79026 46102
rect 79094 46046 79150 46102
rect 79218 46046 79274 46102
rect 79342 46046 79398 46102
rect 78970 45922 79026 45978
rect 79094 45922 79150 45978
rect 79218 45922 79274 45978
rect 79342 45922 79398 45978
rect 78970 28294 79026 28350
rect 79094 28294 79150 28350
rect 79218 28294 79274 28350
rect 79342 28294 79398 28350
rect 78970 28170 79026 28226
rect 79094 28170 79150 28226
rect 79218 28170 79274 28226
rect 79342 28170 79398 28226
rect 78970 28046 79026 28102
rect 79094 28046 79150 28102
rect 79218 28046 79274 28102
rect 79342 28046 79398 28102
rect 78970 27922 79026 27978
rect 79094 27922 79150 27978
rect 79218 27922 79274 27978
rect 79342 27922 79398 27978
rect 78970 10294 79026 10350
rect 79094 10294 79150 10350
rect 79218 10294 79274 10350
rect 79342 10294 79398 10350
rect 78970 10170 79026 10226
rect 79094 10170 79150 10226
rect 79218 10170 79274 10226
rect 79342 10170 79398 10226
rect 78970 10046 79026 10102
rect 79094 10046 79150 10102
rect 79218 10046 79274 10102
rect 79342 10046 79398 10102
rect 78970 9922 79026 9978
rect 79094 9922 79150 9978
rect 79218 9922 79274 9978
rect 79342 9922 79398 9978
rect 78970 -1176 79026 -1120
rect 79094 -1176 79150 -1120
rect 79218 -1176 79274 -1120
rect 79342 -1176 79398 -1120
rect 78970 -1300 79026 -1244
rect 79094 -1300 79150 -1244
rect 79218 -1300 79274 -1244
rect 79342 -1300 79398 -1244
rect 78970 -1424 79026 -1368
rect 79094 -1424 79150 -1368
rect 79218 -1424 79274 -1368
rect 79342 -1424 79398 -1368
rect 78970 -1548 79026 -1492
rect 79094 -1548 79150 -1492
rect 79218 -1548 79274 -1492
rect 79342 -1548 79398 -1492
rect 93250 597156 93306 597212
rect 93374 597156 93430 597212
rect 93498 597156 93554 597212
rect 93622 597156 93678 597212
rect 93250 597032 93306 597088
rect 93374 597032 93430 597088
rect 93498 597032 93554 597088
rect 93622 597032 93678 597088
rect 93250 596908 93306 596964
rect 93374 596908 93430 596964
rect 93498 596908 93554 596964
rect 93622 596908 93678 596964
rect 93250 596784 93306 596840
rect 93374 596784 93430 596840
rect 93498 596784 93554 596840
rect 93622 596784 93678 596840
rect 93250 580294 93306 580350
rect 93374 580294 93430 580350
rect 93498 580294 93554 580350
rect 93622 580294 93678 580350
rect 93250 580170 93306 580226
rect 93374 580170 93430 580226
rect 93498 580170 93554 580226
rect 93622 580170 93678 580226
rect 93250 580046 93306 580102
rect 93374 580046 93430 580102
rect 93498 580046 93554 580102
rect 93622 580046 93678 580102
rect 93250 579922 93306 579978
rect 93374 579922 93430 579978
rect 93498 579922 93554 579978
rect 93622 579922 93678 579978
rect 93250 562294 93306 562350
rect 93374 562294 93430 562350
rect 93498 562294 93554 562350
rect 93622 562294 93678 562350
rect 93250 562170 93306 562226
rect 93374 562170 93430 562226
rect 93498 562170 93554 562226
rect 93622 562170 93678 562226
rect 93250 562046 93306 562102
rect 93374 562046 93430 562102
rect 93498 562046 93554 562102
rect 93622 562046 93678 562102
rect 93250 561922 93306 561978
rect 93374 561922 93430 561978
rect 93498 561922 93554 561978
rect 93622 561922 93678 561978
rect 93250 544294 93306 544350
rect 93374 544294 93430 544350
rect 93498 544294 93554 544350
rect 93622 544294 93678 544350
rect 93250 544170 93306 544226
rect 93374 544170 93430 544226
rect 93498 544170 93554 544226
rect 93622 544170 93678 544226
rect 93250 544046 93306 544102
rect 93374 544046 93430 544102
rect 93498 544046 93554 544102
rect 93622 544046 93678 544102
rect 93250 543922 93306 543978
rect 93374 543922 93430 543978
rect 93498 543922 93554 543978
rect 93622 543922 93678 543978
rect 93250 526294 93306 526350
rect 93374 526294 93430 526350
rect 93498 526294 93554 526350
rect 93622 526294 93678 526350
rect 93250 526170 93306 526226
rect 93374 526170 93430 526226
rect 93498 526170 93554 526226
rect 93622 526170 93678 526226
rect 93250 526046 93306 526102
rect 93374 526046 93430 526102
rect 93498 526046 93554 526102
rect 93622 526046 93678 526102
rect 93250 525922 93306 525978
rect 93374 525922 93430 525978
rect 93498 525922 93554 525978
rect 93622 525922 93678 525978
rect 93250 508294 93306 508350
rect 93374 508294 93430 508350
rect 93498 508294 93554 508350
rect 93622 508294 93678 508350
rect 93250 508170 93306 508226
rect 93374 508170 93430 508226
rect 93498 508170 93554 508226
rect 93622 508170 93678 508226
rect 93250 508046 93306 508102
rect 93374 508046 93430 508102
rect 93498 508046 93554 508102
rect 93622 508046 93678 508102
rect 93250 507922 93306 507978
rect 93374 507922 93430 507978
rect 93498 507922 93554 507978
rect 93622 507922 93678 507978
rect 93250 490294 93306 490350
rect 93374 490294 93430 490350
rect 93498 490294 93554 490350
rect 93622 490294 93678 490350
rect 93250 490170 93306 490226
rect 93374 490170 93430 490226
rect 93498 490170 93554 490226
rect 93622 490170 93678 490226
rect 93250 490046 93306 490102
rect 93374 490046 93430 490102
rect 93498 490046 93554 490102
rect 93622 490046 93678 490102
rect 93250 489922 93306 489978
rect 93374 489922 93430 489978
rect 93498 489922 93554 489978
rect 93622 489922 93678 489978
rect 93250 472294 93306 472350
rect 93374 472294 93430 472350
rect 93498 472294 93554 472350
rect 93622 472294 93678 472350
rect 93250 472170 93306 472226
rect 93374 472170 93430 472226
rect 93498 472170 93554 472226
rect 93622 472170 93678 472226
rect 93250 472046 93306 472102
rect 93374 472046 93430 472102
rect 93498 472046 93554 472102
rect 93622 472046 93678 472102
rect 93250 471922 93306 471978
rect 93374 471922 93430 471978
rect 93498 471922 93554 471978
rect 93622 471922 93678 471978
rect 93250 454294 93306 454350
rect 93374 454294 93430 454350
rect 93498 454294 93554 454350
rect 93622 454294 93678 454350
rect 93250 454170 93306 454226
rect 93374 454170 93430 454226
rect 93498 454170 93554 454226
rect 93622 454170 93678 454226
rect 93250 454046 93306 454102
rect 93374 454046 93430 454102
rect 93498 454046 93554 454102
rect 93622 454046 93678 454102
rect 93250 453922 93306 453978
rect 93374 453922 93430 453978
rect 93498 453922 93554 453978
rect 93622 453922 93678 453978
rect 93250 436294 93306 436350
rect 93374 436294 93430 436350
rect 93498 436294 93554 436350
rect 93622 436294 93678 436350
rect 93250 436170 93306 436226
rect 93374 436170 93430 436226
rect 93498 436170 93554 436226
rect 93622 436170 93678 436226
rect 93250 436046 93306 436102
rect 93374 436046 93430 436102
rect 93498 436046 93554 436102
rect 93622 436046 93678 436102
rect 93250 435922 93306 435978
rect 93374 435922 93430 435978
rect 93498 435922 93554 435978
rect 93622 435922 93678 435978
rect 93250 418294 93306 418350
rect 93374 418294 93430 418350
rect 93498 418294 93554 418350
rect 93622 418294 93678 418350
rect 93250 418170 93306 418226
rect 93374 418170 93430 418226
rect 93498 418170 93554 418226
rect 93622 418170 93678 418226
rect 93250 418046 93306 418102
rect 93374 418046 93430 418102
rect 93498 418046 93554 418102
rect 93622 418046 93678 418102
rect 93250 417922 93306 417978
rect 93374 417922 93430 417978
rect 93498 417922 93554 417978
rect 93622 417922 93678 417978
rect 93250 400294 93306 400350
rect 93374 400294 93430 400350
rect 93498 400294 93554 400350
rect 93622 400294 93678 400350
rect 93250 400170 93306 400226
rect 93374 400170 93430 400226
rect 93498 400170 93554 400226
rect 93622 400170 93678 400226
rect 93250 400046 93306 400102
rect 93374 400046 93430 400102
rect 93498 400046 93554 400102
rect 93622 400046 93678 400102
rect 93250 399922 93306 399978
rect 93374 399922 93430 399978
rect 93498 399922 93554 399978
rect 93622 399922 93678 399978
rect 93250 382294 93306 382350
rect 93374 382294 93430 382350
rect 93498 382294 93554 382350
rect 93622 382294 93678 382350
rect 93250 382170 93306 382226
rect 93374 382170 93430 382226
rect 93498 382170 93554 382226
rect 93622 382170 93678 382226
rect 93250 382046 93306 382102
rect 93374 382046 93430 382102
rect 93498 382046 93554 382102
rect 93622 382046 93678 382102
rect 93250 381922 93306 381978
rect 93374 381922 93430 381978
rect 93498 381922 93554 381978
rect 93622 381922 93678 381978
rect 93250 364294 93306 364350
rect 93374 364294 93430 364350
rect 93498 364294 93554 364350
rect 93622 364294 93678 364350
rect 93250 364170 93306 364226
rect 93374 364170 93430 364226
rect 93498 364170 93554 364226
rect 93622 364170 93678 364226
rect 93250 364046 93306 364102
rect 93374 364046 93430 364102
rect 93498 364046 93554 364102
rect 93622 364046 93678 364102
rect 93250 363922 93306 363978
rect 93374 363922 93430 363978
rect 93498 363922 93554 363978
rect 93622 363922 93678 363978
rect 93250 346294 93306 346350
rect 93374 346294 93430 346350
rect 93498 346294 93554 346350
rect 93622 346294 93678 346350
rect 93250 346170 93306 346226
rect 93374 346170 93430 346226
rect 93498 346170 93554 346226
rect 93622 346170 93678 346226
rect 93250 346046 93306 346102
rect 93374 346046 93430 346102
rect 93498 346046 93554 346102
rect 93622 346046 93678 346102
rect 93250 345922 93306 345978
rect 93374 345922 93430 345978
rect 93498 345922 93554 345978
rect 93622 345922 93678 345978
rect 93250 328294 93306 328350
rect 93374 328294 93430 328350
rect 93498 328294 93554 328350
rect 93622 328294 93678 328350
rect 93250 328170 93306 328226
rect 93374 328170 93430 328226
rect 93498 328170 93554 328226
rect 93622 328170 93678 328226
rect 93250 328046 93306 328102
rect 93374 328046 93430 328102
rect 93498 328046 93554 328102
rect 93622 328046 93678 328102
rect 93250 327922 93306 327978
rect 93374 327922 93430 327978
rect 93498 327922 93554 327978
rect 93622 327922 93678 327978
rect 93250 310294 93306 310350
rect 93374 310294 93430 310350
rect 93498 310294 93554 310350
rect 93622 310294 93678 310350
rect 93250 310170 93306 310226
rect 93374 310170 93430 310226
rect 93498 310170 93554 310226
rect 93622 310170 93678 310226
rect 93250 310046 93306 310102
rect 93374 310046 93430 310102
rect 93498 310046 93554 310102
rect 93622 310046 93678 310102
rect 93250 309922 93306 309978
rect 93374 309922 93430 309978
rect 93498 309922 93554 309978
rect 93622 309922 93678 309978
rect 93250 292294 93306 292350
rect 93374 292294 93430 292350
rect 93498 292294 93554 292350
rect 93622 292294 93678 292350
rect 93250 292170 93306 292226
rect 93374 292170 93430 292226
rect 93498 292170 93554 292226
rect 93622 292170 93678 292226
rect 93250 292046 93306 292102
rect 93374 292046 93430 292102
rect 93498 292046 93554 292102
rect 93622 292046 93678 292102
rect 93250 291922 93306 291978
rect 93374 291922 93430 291978
rect 93498 291922 93554 291978
rect 93622 291922 93678 291978
rect 93250 274294 93306 274350
rect 93374 274294 93430 274350
rect 93498 274294 93554 274350
rect 93622 274294 93678 274350
rect 93250 274170 93306 274226
rect 93374 274170 93430 274226
rect 93498 274170 93554 274226
rect 93622 274170 93678 274226
rect 93250 274046 93306 274102
rect 93374 274046 93430 274102
rect 93498 274046 93554 274102
rect 93622 274046 93678 274102
rect 93250 273922 93306 273978
rect 93374 273922 93430 273978
rect 93498 273922 93554 273978
rect 93622 273922 93678 273978
rect 93250 256294 93306 256350
rect 93374 256294 93430 256350
rect 93498 256294 93554 256350
rect 93622 256294 93678 256350
rect 93250 256170 93306 256226
rect 93374 256170 93430 256226
rect 93498 256170 93554 256226
rect 93622 256170 93678 256226
rect 93250 256046 93306 256102
rect 93374 256046 93430 256102
rect 93498 256046 93554 256102
rect 93622 256046 93678 256102
rect 93250 255922 93306 255978
rect 93374 255922 93430 255978
rect 93498 255922 93554 255978
rect 93622 255922 93678 255978
rect 93250 238294 93306 238350
rect 93374 238294 93430 238350
rect 93498 238294 93554 238350
rect 93622 238294 93678 238350
rect 93250 238170 93306 238226
rect 93374 238170 93430 238226
rect 93498 238170 93554 238226
rect 93622 238170 93678 238226
rect 93250 238046 93306 238102
rect 93374 238046 93430 238102
rect 93498 238046 93554 238102
rect 93622 238046 93678 238102
rect 93250 237922 93306 237978
rect 93374 237922 93430 237978
rect 93498 237922 93554 237978
rect 93622 237922 93678 237978
rect 93250 220294 93306 220350
rect 93374 220294 93430 220350
rect 93498 220294 93554 220350
rect 93622 220294 93678 220350
rect 93250 220170 93306 220226
rect 93374 220170 93430 220226
rect 93498 220170 93554 220226
rect 93622 220170 93678 220226
rect 93250 220046 93306 220102
rect 93374 220046 93430 220102
rect 93498 220046 93554 220102
rect 93622 220046 93678 220102
rect 93250 219922 93306 219978
rect 93374 219922 93430 219978
rect 93498 219922 93554 219978
rect 93622 219922 93678 219978
rect 93250 202294 93306 202350
rect 93374 202294 93430 202350
rect 93498 202294 93554 202350
rect 93622 202294 93678 202350
rect 93250 202170 93306 202226
rect 93374 202170 93430 202226
rect 93498 202170 93554 202226
rect 93622 202170 93678 202226
rect 93250 202046 93306 202102
rect 93374 202046 93430 202102
rect 93498 202046 93554 202102
rect 93622 202046 93678 202102
rect 93250 201922 93306 201978
rect 93374 201922 93430 201978
rect 93498 201922 93554 201978
rect 93622 201922 93678 201978
rect 93250 184294 93306 184350
rect 93374 184294 93430 184350
rect 93498 184294 93554 184350
rect 93622 184294 93678 184350
rect 93250 184170 93306 184226
rect 93374 184170 93430 184226
rect 93498 184170 93554 184226
rect 93622 184170 93678 184226
rect 93250 184046 93306 184102
rect 93374 184046 93430 184102
rect 93498 184046 93554 184102
rect 93622 184046 93678 184102
rect 93250 183922 93306 183978
rect 93374 183922 93430 183978
rect 93498 183922 93554 183978
rect 93622 183922 93678 183978
rect 93250 166294 93306 166350
rect 93374 166294 93430 166350
rect 93498 166294 93554 166350
rect 93622 166294 93678 166350
rect 93250 166170 93306 166226
rect 93374 166170 93430 166226
rect 93498 166170 93554 166226
rect 93622 166170 93678 166226
rect 93250 166046 93306 166102
rect 93374 166046 93430 166102
rect 93498 166046 93554 166102
rect 93622 166046 93678 166102
rect 93250 165922 93306 165978
rect 93374 165922 93430 165978
rect 93498 165922 93554 165978
rect 93622 165922 93678 165978
rect 93250 148294 93306 148350
rect 93374 148294 93430 148350
rect 93498 148294 93554 148350
rect 93622 148294 93678 148350
rect 93250 148170 93306 148226
rect 93374 148170 93430 148226
rect 93498 148170 93554 148226
rect 93622 148170 93678 148226
rect 93250 148046 93306 148102
rect 93374 148046 93430 148102
rect 93498 148046 93554 148102
rect 93622 148046 93678 148102
rect 93250 147922 93306 147978
rect 93374 147922 93430 147978
rect 93498 147922 93554 147978
rect 93622 147922 93678 147978
rect 93250 130294 93306 130350
rect 93374 130294 93430 130350
rect 93498 130294 93554 130350
rect 93622 130294 93678 130350
rect 93250 130170 93306 130226
rect 93374 130170 93430 130226
rect 93498 130170 93554 130226
rect 93622 130170 93678 130226
rect 93250 130046 93306 130102
rect 93374 130046 93430 130102
rect 93498 130046 93554 130102
rect 93622 130046 93678 130102
rect 93250 129922 93306 129978
rect 93374 129922 93430 129978
rect 93498 129922 93554 129978
rect 93622 129922 93678 129978
rect 93250 112294 93306 112350
rect 93374 112294 93430 112350
rect 93498 112294 93554 112350
rect 93622 112294 93678 112350
rect 93250 112170 93306 112226
rect 93374 112170 93430 112226
rect 93498 112170 93554 112226
rect 93622 112170 93678 112226
rect 93250 112046 93306 112102
rect 93374 112046 93430 112102
rect 93498 112046 93554 112102
rect 93622 112046 93678 112102
rect 93250 111922 93306 111978
rect 93374 111922 93430 111978
rect 93498 111922 93554 111978
rect 93622 111922 93678 111978
rect 93250 94294 93306 94350
rect 93374 94294 93430 94350
rect 93498 94294 93554 94350
rect 93622 94294 93678 94350
rect 93250 94170 93306 94226
rect 93374 94170 93430 94226
rect 93498 94170 93554 94226
rect 93622 94170 93678 94226
rect 93250 94046 93306 94102
rect 93374 94046 93430 94102
rect 93498 94046 93554 94102
rect 93622 94046 93678 94102
rect 93250 93922 93306 93978
rect 93374 93922 93430 93978
rect 93498 93922 93554 93978
rect 93622 93922 93678 93978
rect 93250 76294 93306 76350
rect 93374 76294 93430 76350
rect 93498 76294 93554 76350
rect 93622 76294 93678 76350
rect 93250 76170 93306 76226
rect 93374 76170 93430 76226
rect 93498 76170 93554 76226
rect 93622 76170 93678 76226
rect 93250 76046 93306 76102
rect 93374 76046 93430 76102
rect 93498 76046 93554 76102
rect 93622 76046 93678 76102
rect 93250 75922 93306 75978
rect 93374 75922 93430 75978
rect 93498 75922 93554 75978
rect 93622 75922 93678 75978
rect 93250 58294 93306 58350
rect 93374 58294 93430 58350
rect 93498 58294 93554 58350
rect 93622 58294 93678 58350
rect 93250 58170 93306 58226
rect 93374 58170 93430 58226
rect 93498 58170 93554 58226
rect 93622 58170 93678 58226
rect 93250 58046 93306 58102
rect 93374 58046 93430 58102
rect 93498 58046 93554 58102
rect 93622 58046 93678 58102
rect 93250 57922 93306 57978
rect 93374 57922 93430 57978
rect 93498 57922 93554 57978
rect 93622 57922 93678 57978
rect 93250 40294 93306 40350
rect 93374 40294 93430 40350
rect 93498 40294 93554 40350
rect 93622 40294 93678 40350
rect 93250 40170 93306 40226
rect 93374 40170 93430 40226
rect 93498 40170 93554 40226
rect 93622 40170 93678 40226
rect 93250 40046 93306 40102
rect 93374 40046 93430 40102
rect 93498 40046 93554 40102
rect 93622 40046 93678 40102
rect 93250 39922 93306 39978
rect 93374 39922 93430 39978
rect 93498 39922 93554 39978
rect 93622 39922 93678 39978
rect 93250 22294 93306 22350
rect 93374 22294 93430 22350
rect 93498 22294 93554 22350
rect 93622 22294 93678 22350
rect 93250 22170 93306 22226
rect 93374 22170 93430 22226
rect 93498 22170 93554 22226
rect 93622 22170 93678 22226
rect 93250 22046 93306 22102
rect 93374 22046 93430 22102
rect 93498 22046 93554 22102
rect 93622 22046 93678 22102
rect 93250 21922 93306 21978
rect 93374 21922 93430 21978
rect 93498 21922 93554 21978
rect 93622 21922 93678 21978
rect 93250 4294 93306 4350
rect 93374 4294 93430 4350
rect 93498 4294 93554 4350
rect 93622 4294 93678 4350
rect 93250 4170 93306 4226
rect 93374 4170 93430 4226
rect 93498 4170 93554 4226
rect 93622 4170 93678 4226
rect 93250 4046 93306 4102
rect 93374 4046 93430 4102
rect 93498 4046 93554 4102
rect 93622 4046 93678 4102
rect 93250 3922 93306 3978
rect 93374 3922 93430 3978
rect 93498 3922 93554 3978
rect 93622 3922 93678 3978
rect 93250 -216 93306 -160
rect 93374 -216 93430 -160
rect 93498 -216 93554 -160
rect 93622 -216 93678 -160
rect 93250 -340 93306 -284
rect 93374 -340 93430 -284
rect 93498 -340 93554 -284
rect 93622 -340 93678 -284
rect 93250 -464 93306 -408
rect 93374 -464 93430 -408
rect 93498 -464 93554 -408
rect 93622 -464 93678 -408
rect 93250 -588 93306 -532
rect 93374 -588 93430 -532
rect 93498 -588 93554 -532
rect 93622 -588 93678 -532
rect 96970 598116 97026 598172
rect 97094 598116 97150 598172
rect 97218 598116 97274 598172
rect 97342 598116 97398 598172
rect 96970 597992 97026 598048
rect 97094 597992 97150 598048
rect 97218 597992 97274 598048
rect 97342 597992 97398 598048
rect 96970 597868 97026 597924
rect 97094 597868 97150 597924
rect 97218 597868 97274 597924
rect 97342 597868 97398 597924
rect 96970 597744 97026 597800
rect 97094 597744 97150 597800
rect 97218 597744 97274 597800
rect 97342 597744 97398 597800
rect 96970 586294 97026 586350
rect 97094 586294 97150 586350
rect 97218 586294 97274 586350
rect 97342 586294 97398 586350
rect 96970 586170 97026 586226
rect 97094 586170 97150 586226
rect 97218 586170 97274 586226
rect 97342 586170 97398 586226
rect 96970 586046 97026 586102
rect 97094 586046 97150 586102
rect 97218 586046 97274 586102
rect 97342 586046 97398 586102
rect 96970 585922 97026 585978
rect 97094 585922 97150 585978
rect 97218 585922 97274 585978
rect 97342 585922 97398 585978
rect 96970 568294 97026 568350
rect 97094 568294 97150 568350
rect 97218 568294 97274 568350
rect 97342 568294 97398 568350
rect 96970 568170 97026 568226
rect 97094 568170 97150 568226
rect 97218 568170 97274 568226
rect 97342 568170 97398 568226
rect 96970 568046 97026 568102
rect 97094 568046 97150 568102
rect 97218 568046 97274 568102
rect 97342 568046 97398 568102
rect 96970 567922 97026 567978
rect 97094 567922 97150 567978
rect 97218 567922 97274 567978
rect 97342 567922 97398 567978
rect 96970 550294 97026 550350
rect 97094 550294 97150 550350
rect 97218 550294 97274 550350
rect 97342 550294 97398 550350
rect 96970 550170 97026 550226
rect 97094 550170 97150 550226
rect 97218 550170 97274 550226
rect 97342 550170 97398 550226
rect 96970 550046 97026 550102
rect 97094 550046 97150 550102
rect 97218 550046 97274 550102
rect 97342 550046 97398 550102
rect 96970 549922 97026 549978
rect 97094 549922 97150 549978
rect 97218 549922 97274 549978
rect 97342 549922 97398 549978
rect 96970 532294 97026 532350
rect 97094 532294 97150 532350
rect 97218 532294 97274 532350
rect 97342 532294 97398 532350
rect 96970 532170 97026 532226
rect 97094 532170 97150 532226
rect 97218 532170 97274 532226
rect 97342 532170 97398 532226
rect 96970 532046 97026 532102
rect 97094 532046 97150 532102
rect 97218 532046 97274 532102
rect 97342 532046 97398 532102
rect 96970 531922 97026 531978
rect 97094 531922 97150 531978
rect 97218 531922 97274 531978
rect 97342 531922 97398 531978
rect 96970 514294 97026 514350
rect 97094 514294 97150 514350
rect 97218 514294 97274 514350
rect 97342 514294 97398 514350
rect 96970 514170 97026 514226
rect 97094 514170 97150 514226
rect 97218 514170 97274 514226
rect 97342 514170 97398 514226
rect 96970 514046 97026 514102
rect 97094 514046 97150 514102
rect 97218 514046 97274 514102
rect 97342 514046 97398 514102
rect 96970 513922 97026 513978
rect 97094 513922 97150 513978
rect 97218 513922 97274 513978
rect 97342 513922 97398 513978
rect 96970 496294 97026 496350
rect 97094 496294 97150 496350
rect 97218 496294 97274 496350
rect 97342 496294 97398 496350
rect 96970 496170 97026 496226
rect 97094 496170 97150 496226
rect 97218 496170 97274 496226
rect 97342 496170 97398 496226
rect 96970 496046 97026 496102
rect 97094 496046 97150 496102
rect 97218 496046 97274 496102
rect 97342 496046 97398 496102
rect 96970 495922 97026 495978
rect 97094 495922 97150 495978
rect 97218 495922 97274 495978
rect 97342 495922 97398 495978
rect 96970 478294 97026 478350
rect 97094 478294 97150 478350
rect 97218 478294 97274 478350
rect 97342 478294 97398 478350
rect 96970 478170 97026 478226
rect 97094 478170 97150 478226
rect 97218 478170 97274 478226
rect 97342 478170 97398 478226
rect 96970 478046 97026 478102
rect 97094 478046 97150 478102
rect 97218 478046 97274 478102
rect 97342 478046 97398 478102
rect 96970 477922 97026 477978
rect 97094 477922 97150 477978
rect 97218 477922 97274 477978
rect 97342 477922 97398 477978
rect 96970 460294 97026 460350
rect 97094 460294 97150 460350
rect 97218 460294 97274 460350
rect 97342 460294 97398 460350
rect 96970 460170 97026 460226
rect 97094 460170 97150 460226
rect 97218 460170 97274 460226
rect 97342 460170 97398 460226
rect 96970 460046 97026 460102
rect 97094 460046 97150 460102
rect 97218 460046 97274 460102
rect 97342 460046 97398 460102
rect 96970 459922 97026 459978
rect 97094 459922 97150 459978
rect 97218 459922 97274 459978
rect 97342 459922 97398 459978
rect 96970 442294 97026 442350
rect 97094 442294 97150 442350
rect 97218 442294 97274 442350
rect 97342 442294 97398 442350
rect 96970 442170 97026 442226
rect 97094 442170 97150 442226
rect 97218 442170 97274 442226
rect 97342 442170 97398 442226
rect 96970 442046 97026 442102
rect 97094 442046 97150 442102
rect 97218 442046 97274 442102
rect 97342 442046 97398 442102
rect 96970 441922 97026 441978
rect 97094 441922 97150 441978
rect 97218 441922 97274 441978
rect 97342 441922 97398 441978
rect 96970 424294 97026 424350
rect 97094 424294 97150 424350
rect 97218 424294 97274 424350
rect 97342 424294 97398 424350
rect 96970 424170 97026 424226
rect 97094 424170 97150 424226
rect 97218 424170 97274 424226
rect 97342 424170 97398 424226
rect 96970 424046 97026 424102
rect 97094 424046 97150 424102
rect 97218 424046 97274 424102
rect 97342 424046 97398 424102
rect 96970 423922 97026 423978
rect 97094 423922 97150 423978
rect 97218 423922 97274 423978
rect 97342 423922 97398 423978
rect 96970 406294 97026 406350
rect 97094 406294 97150 406350
rect 97218 406294 97274 406350
rect 97342 406294 97398 406350
rect 96970 406170 97026 406226
rect 97094 406170 97150 406226
rect 97218 406170 97274 406226
rect 97342 406170 97398 406226
rect 96970 406046 97026 406102
rect 97094 406046 97150 406102
rect 97218 406046 97274 406102
rect 97342 406046 97398 406102
rect 96970 405922 97026 405978
rect 97094 405922 97150 405978
rect 97218 405922 97274 405978
rect 97342 405922 97398 405978
rect 96970 388294 97026 388350
rect 97094 388294 97150 388350
rect 97218 388294 97274 388350
rect 97342 388294 97398 388350
rect 96970 388170 97026 388226
rect 97094 388170 97150 388226
rect 97218 388170 97274 388226
rect 97342 388170 97398 388226
rect 96970 388046 97026 388102
rect 97094 388046 97150 388102
rect 97218 388046 97274 388102
rect 97342 388046 97398 388102
rect 96970 387922 97026 387978
rect 97094 387922 97150 387978
rect 97218 387922 97274 387978
rect 97342 387922 97398 387978
rect 96970 370294 97026 370350
rect 97094 370294 97150 370350
rect 97218 370294 97274 370350
rect 97342 370294 97398 370350
rect 96970 370170 97026 370226
rect 97094 370170 97150 370226
rect 97218 370170 97274 370226
rect 97342 370170 97398 370226
rect 96970 370046 97026 370102
rect 97094 370046 97150 370102
rect 97218 370046 97274 370102
rect 97342 370046 97398 370102
rect 96970 369922 97026 369978
rect 97094 369922 97150 369978
rect 97218 369922 97274 369978
rect 97342 369922 97398 369978
rect 96970 352294 97026 352350
rect 97094 352294 97150 352350
rect 97218 352294 97274 352350
rect 97342 352294 97398 352350
rect 96970 352170 97026 352226
rect 97094 352170 97150 352226
rect 97218 352170 97274 352226
rect 97342 352170 97398 352226
rect 96970 352046 97026 352102
rect 97094 352046 97150 352102
rect 97218 352046 97274 352102
rect 97342 352046 97398 352102
rect 96970 351922 97026 351978
rect 97094 351922 97150 351978
rect 97218 351922 97274 351978
rect 97342 351922 97398 351978
rect 96970 334294 97026 334350
rect 97094 334294 97150 334350
rect 97218 334294 97274 334350
rect 97342 334294 97398 334350
rect 96970 334170 97026 334226
rect 97094 334170 97150 334226
rect 97218 334170 97274 334226
rect 97342 334170 97398 334226
rect 96970 334046 97026 334102
rect 97094 334046 97150 334102
rect 97218 334046 97274 334102
rect 97342 334046 97398 334102
rect 96970 333922 97026 333978
rect 97094 333922 97150 333978
rect 97218 333922 97274 333978
rect 97342 333922 97398 333978
rect 96970 316294 97026 316350
rect 97094 316294 97150 316350
rect 97218 316294 97274 316350
rect 97342 316294 97398 316350
rect 96970 316170 97026 316226
rect 97094 316170 97150 316226
rect 97218 316170 97274 316226
rect 97342 316170 97398 316226
rect 96970 316046 97026 316102
rect 97094 316046 97150 316102
rect 97218 316046 97274 316102
rect 97342 316046 97398 316102
rect 96970 315922 97026 315978
rect 97094 315922 97150 315978
rect 97218 315922 97274 315978
rect 97342 315922 97398 315978
rect 96970 298294 97026 298350
rect 97094 298294 97150 298350
rect 97218 298294 97274 298350
rect 97342 298294 97398 298350
rect 96970 298170 97026 298226
rect 97094 298170 97150 298226
rect 97218 298170 97274 298226
rect 97342 298170 97398 298226
rect 96970 298046 97026 298102
rect 97094 298046 97150 298102
rect 97218 298046 97274 298102
rect 97342 298046 97398 298102
rect 96970 297922 97026 297978
rect 97094 297922 97150 297978
rect 97218 297922 97274 297978
rect 97342 297922 97398 297978
rect 96970 280294 97026 280350
rect 97094 280294 97150 280350
rect 97218 280294 97274 280350
rect 97342 280294 97398 280350
rect 96970 280170 97026 280226
rect 97094 280170 97150 280226
rect 97218 280170 97274 280226
rect 97342 280170 97398 280226
rect 96970 280046 97026 280102
rect 97094 280046 97150 280102
rect 97218 280046 97274 280102
rect 97342 280046 97398 280102
rect 96970 279922 97026 279978
rect 97094 279922 97150 279978
rect 97218 279922 97274 279978
rect 97342 279922 97398 279978
rect 96970 262294 97026 262350
rect 97094 262294 97150 262350
rect 97218 262294 97274 262350
rect 97342 262294 97398 262350
rect 96970 262170 97026 262226
rect 97094 262170 97150 262226
rect 97218 262170 97274 262226
rect 97342 262170 97398 262226
rect 96970 262046 97026 262102
rect 97094 262046 97150 262102
rect 97218 262046 97274 262102
rect 97342 262046 97398 262102
rect 96970 261922 97026 261978
rect 97094 261922 97150 261978
rect 97218 261922 97274 261978
rect 97342 261922 97398 261978
rect 96970 244294 97026 244350
rect 97094 244294 97150 244350
rect 97218 244294 97274 244350
rect 97342 244294 97398 244350
rect 96970 244170 97026 244226
rect 97094 244170 97150 244226
rect 97218 244170 97274 244226
rect 97342 244170 97398 244226
rect 96970 244046 97026 244102
rect 97094 244046 97150 244102
rect 97218 244046 97274 244102
rect 97342 244046 97398 244102
rect 96970 243922 97026 243978
rect 97094 243922 97150 243978
rect 97218 243922 97274 243978
rect 97342 243922 97398 243978
rect 96970 226294 97026 226350
rect 97094 226294 97150 226350
rect 97218 226294 97274 226350
rect 97342 226294 97398 226350
rect 96970 226170 97026 226226
rect 97094 226170 97150 226226
rect 97218 226170 97274 226226
rect 97342 226170 97398 226226
rect 96970 226046 97026 226102
rect 97094 226046 97150 226102
rect 97218 226046 97274 226102
rect 97342 226046 97398 226102
rect 96970 225922 97026 225978
rect 97094 225922 97150 225978
rect 97218 225922 97274 225978
rect 97342 225922 97398 225978
rect 96970 208294 97026 208350
rect 97094 208294 97150 208350
rect 97218 208294 97274 208350
rect 97342 208294 97398 208350
rect 96970 208170 97026 208226
rect 97094 208170 97150 208226
rect 97218 208170 97274 208226
rect 97342 208170 97398 208226
rect 96970 208046 97026 208102
rect 97094 208046 97150 208102
rect 97218 208046 97274 208102
rect 97342 208046 97398 208102
rect 96970 207922 97026 207978
rect 97094 207922 97150 207978
rect 97218 207922 97274 207978
rect 97342 207922 97398 207978
rect 96970 190294 97026 190350
rect 97094 190294 97150 190350
rect 97218 190294 97274 190350
rect 97342 190294 97398 190350
rect 96970 190170 97026 190226
rect 97094 190170 97150 190226
rect 97218 190170 97274 190226
rect 97342 190170 97398 190226
rect 96970 190046 97026 190102
rect 97094 190046 97150 190102
rect 97218 190046 97274 190102
rect 97342 190046 97398 190102
rect 96970 189922 97026 189978
rect 97094 189922 97150 189978
rect 97218 189922 97274 189978
rect 97342 189922 97398 189978
rect 96970 172294 97026 172350
rect 97094 172294 97150 172350
rect 97218 172294 97274 172350
rect 97342 172294 97398 172350
rect 96970 172170 97026 172226
rect 97094 172170 97150 172226
rect 97218 172170 97274 172226
rect 97342 172170 97398 172226
rect 96970 172046 97026 172102
rect 97094 172046 97150 172102
rect 97218 172046 97274 172102
rect 97342 172046 97398 172102
rect 96970 171922 97026 171978
rect 97094 171922 97150 171978
rect 97218 171922 97274 171978
rect 97342 171922 97398 171978
rect 96970 154294 97026 154350
rect 97094 154294 97150 154350
rect 97218 154294 97274 154350
rect 97342 154294 97398 154350
rect 96970 154170 97026 154226
rect 97094 154170 97150 154226
rect 97218 154170 97274 154226
rect 97342 154170 97398 154226
rect 96970 154046 97026 154102
rect 97094 154046 97150 154102
rect 97218 154046 97274 154102
rect 97342 154046 97398 154102
rect 96970 153922 97026 153978
rect 97094 153922 97150 153978
rect 97218 153922 97274 153978
rect 97342 153922 97398 153978
rect 96970 136294 97026 136350
rect 97094 136294 97150 136350
rect 97218 136294 97274 136350
rect 97342 136294 97398 136350
rect 96970 136170 97026 136226
rect 97094 136170 97150 136226
rect 97218 136170 97274 136226
rect 97342 136170 97398 136226
rect 96970 136046 97026 136102
rect 97094 136046 97150 136102
rect 97218 136046 97274 136102
rect 97342 136046 97398 136102
rect 96970 135922 97026 135978
rect 97094 135922 97150 135978
rect 97218 135922 97274 135978
rect 97342 135922 97398 135978
rect 96970 118294 97026 118350
rect 97094 118294 97150 118350
rect 97218 118294 97274 118350
rect 97342 118294 97398 118350
rect 96970 118170 97026 118226
rect 97094 118170 97150 118226
rect 97218 118170 97274 118226
rect 97342 118170 97398 118226
rect 96970 118046 97026 118102
rect 97094 118046 97150 118102
rect 97218 118046 97274 118102
rect 97342 118046 97398 118102
rect 96970 117922 97026 117978
rect 97094 117922 97150 117978
rect 97218 117922 97274 117978
rect 97342 117922 97398 117978
rect 96970 100294 97026 100350
rect 97094 100294 97150 100350
rect 97218 100294 97274 100350
rect 97342 100294 97398 100350
rect 96970 100170 97026 100226
rect 97094 100170 97150 100226
rect 97218 100170 97274 100226
rect 97342 100170 97398 100226
rect 96970 100046 97026 100102
rect 97094 100046 97150 100102
rect 97218 100046 97274 100102
rect 97342 100046 97398 100102
rect 96970 99922 97026 99978
rect 97094 99922 97150 99978
rect 97218 99922 97274 99978
rect 97342 99922 97398 99978
rect 96970 82294 97026 82350
rect 97094 82294 97150 82350
rect 97218 82294 97274 82350
rect 97342 82294 97398 82350
rect 96970 82170 97026 82226
rect 97094 82170 97150 82226
rect 97218 82170 97274 82226
rect 97342 82170 97398 82226
rect 96970 82046 97026 82102
rect 97094 82046 97150 82102
rect 97218 82046 97274 82102
rect 97342 82046 97398 82102
rect 96970 81922 97026 81978
rect 97094 81922 97150 81978
rect 97218 81922 97274 81978
rect 97342 81922 97398 81978
rect 96970 64294 97026 64350
rect 97094 64294 97150 64350
rect 97218 64294 97274 64350
rect 97342 64294 97398 64350
rect 96970 64170 97026 64226
rect 97094 64170 97150 64226
rect 97218 64170 97274 64226
rect 97342 64170 97398 64226
rect 96970 64046 97026 64102
rect 97094 64046 97150 64102
rect 97218 64046 97274 64102
rect 97342 64046 97398 64102
rect 96970 63922 97026 63978
rect 97094 63922 97150 63978
rect 97218 63922 97274 63978
rect 97342 63922 97398 63978
rect 96970 46294 97026 46350
rect 97094 46294 97150 46350
rect 97218 46294 97274 46350
rect 97342 46294 97398 46350
rect 96970 46170 97026 46226
rect 97094 46170 97150 46226
rect 97218 46170 97274 46226
rect 97342 46170 97398 46226
rect 96970 46046 97026 46102
rect 97094 46046 97150 46102
rect 97218 46046 97274 46102
rect 97342 46046 97398 46102
rect 96970 45922 97026 45978
rect 97094 45922 97150 45978
rect 97218 45922 97274 45978
rect 97342 45922 97398 45978
rect 96970 28294 97026 28350
rect 97094 28294 97150 28350
rect 97218 28294 97274 28350
rect 97342 28294 97398 28350
rect 96970 28170 97026 28226
rect 97094 28170 97150 28226
rect 97218 28170 97274 28226
rect 97342 28170 97398 28226
rect 96970 28046 97026 28102
rect 97094 28046 97150 28102
rect 97218 28046 97274 28102
rect 97342 28046 97398 28102
rect 96970 27922 97026 27978
rect 97094 27922 97150 27978
rect 97218 27922 97274 27978
rect 97342 27922 97398 27978
rect 96970 10294 97026 10350
rect 97094 10294 97150 10350
rect 97218 10294 97274 10350
rect 97342 10294 97398 10350
rect 96970 10170 97026 10226
rect 97094 10170 97150 10226
rect 97218 10170 97274 10226
rect 97342 10170 97398 10226
rect 96970 10046 97026 10102
rect 97094 10046 97150 10102
rect 97218 10046 97274 10102
rect 97342 10046 97398 10102
rect 96970 9922 97026 9978
rect 97094 9922 97150 9978
rect 97218 9922 97274 9978
rect 97342 9922 97398 9978
rect 96970 -1176 97026 -1120
rect 97094 -1176 97150 -1120
rect 97218 -1176 97274 -1120
rect 97342 -1176 97398 -1120
rect 96970 -1300 97026 -1244
rect 97094 -1300 97150 -1244
rect 97218 -1300 97274 -1244
rect 97342 -1300 97398 -1244
rect 96970 -1424 97026 -1368
rect 97094 -1424 97150 -1368
rect 97218 -1424 97274 -1368
rect 97342 -1424 97398 -1368
rect 96970 -1548 97026 -1492
rect 97094 -1548 97150 -1492
rect 97218 -1548 97274 -1492
rect 97342 -1548 97398 -1492
rect 111250 597156 111306 597212
rect 111374 597156 111430 597212
rect 111498 597156 111554 597212
rect 111622 597156 111678 597212
rect 111250 597032 111306 597088
rect 111374 597032 111430 597088
rect 111498 597032 111554 597088
rect 111622 597032 111678 597088
rect 111250 596908 111306 596964
rect 111374 596908 111430 596964
rect 111498 596908 111554 596964
rect 111622 596908 111678 596964
rect 111250 596784 111306 596840
rect 111374 596784 111430 596840
rect 111498 596784 111554 596840
rect 111622 596784 111678 596840
rect 111250 580294 111306 580350
rect 111374 580294 111430 580350
rect 111498 580294 111554 580350
rect 111622 580294 111678 580350
rect 111250 580170 111306 580226
rect 111374 580170 111430 580226
rect 111498 580170 111554 580226
rect 111622 580170 111678 580226
rect 111250 580046 111306 580102
rect 111374 580046 111430 580102
rect 111498 580046 111554 580102
rect 111622 580046 111678 580102
rect 111250 579922 111306 579978
rect 111374 579922 111430 579978
rect 111498 579922 111554 579978
rect 111622 579922 111678 579978
rect 111250 562294 111306 562350
rect 111374 562294 111430 562350
rect 111498 562294 111554 562350
rect 111622 562294 111678 562350
rect 111250 562170 111306 562226
rect 111374 562170 111430 562226
rect 111498 562170 111554 562226
rect 111622 562170 111678 562226
rect 111250 562046 111306 562102
rect 111374 562046 111430 562102
rect 111498 562046 111554 562102
rect 111622 562046 111678 562102
rect 111250 561922 111306 561978
rect 111374 561922 111430 561978
rect 111498 561922 111554 561978
rect 111622 561922 111678 561978
rect 111250 544294 111306 544350
rect 111374 544294 111430 544350
rect 111498 544294 111554 544350
rect 111622 544294 111678 544350
rect 111250 544170 111306 544226
rect 111374 544170 111430 544226
rect 111498 544170 111554 544226
rect 111622 544170 111678 544226
rect 111250 544046 111306 544102
rect 111374 544046 111430 544102
rect 111498 544046 111554 544102
rect 111622 544046 111678 544102
rect 111250 543922 111306 543978
rect 111374 543922 111430 543978
rect 111498 543922 111554 543978
rect 111622 543922 111678 543978
rect 111250 526294 111306 526350
rect 111374 526294 111430 526350
rect 111498 526294 111554 526350
rect 111622 526294 111678 526350
rect 111250 526170 111306 526226
rect 111374 526170 111430 526226
rect 111498 526170 111554 526226
rect 111622 526170 111678 526226
rect 111250 526046 111306 526102
rect 111374 526046 111430 526102
rect 111498 526046 111554 526102
rect 111622 526046 111678 526102
rect 111250 525922 111306 525978
rect 111374 525922 111430 525978
rect 111498 525922 111554 525978
rect 111622 525922 111678 525978
rect 111250 508294 111306 508350
rect 111374 508294 111430 508350
rect 111498 508294 111554 508350
rect 111622 508294 111678 508350
rect 111250 508170 111306 508226
rect 111374 508170 111430 508226
rect 111498 508170 111554 508226
rect 111622 508170 111678 508226
rect 111250 508046 111306 508102
rect 111374 508046 111430 508102
rect 111498 508046 111554 508102
rect 111622 508046 111678 508102
rect 111250 507922 111306 507978
rect 111374 507922 111430 507978
rect 111498 507922 111554 507978
rect 111622 507922 111678 507978
rect 111250 490294 111306 490350
rect 111374 490294 111430 490350
rect 111498 490294 111554 490350
rect 111622 490294 111678 490350
rect 111250 490170 111306 490226
rect 111374 490170 111430 490226
rect 111498 490170 111554 490226
rect 111622 490170 111678 490226
rect 111250 490046 111306 490102
rect 111374 490046 111430 490102
rect 111498 490046 111554 490102
rect 111622 490046 111678 490102
rect 111250 489922 111306 489978
rect 111374 489922 111430 489978
rect 111498 489922 111554 489978
rect 111622 489922 111678 489978
rect 111250 472294 111306 472350
rect 111374 472294 111430 472350
rect 111498 472294 111554 472350
rect 111622 472294 111678 472350
rect 111250 472170 111306 472226
rect 111374 472170 111430 472226
rect 111498 472170 111554 472226
rect 111622 472170 111678 472226
rect 111250 472046 111306 472102
rect 111374 472046 111430 472102
rect 111498 472046 111554 472102
rect 111622 472046 111678 472102
rect 111250 471922 111306 471978
rect 111374 471922 111430 471978
rect 111498 471922 111554 471978
rect 111622 471922 111678 471978
rect 111250 454294 111306 454350
rect 111374 454294 111430 454350
rect 111498 454294 111554 454350
rect 111622 454294 111678 454350
rect 111250 454170 111306 454226
rect 111374 454170 111430 454226
rect 111498 454170 111554 454226
rect 111622 454170 111678 454226
rect 111250 454046 111306 454102
rect 111374 454046 111430 454102
rect 111498 454046 111554 454102
rect 111622 454046 111678 454102
rect 111250 453922 111306 453978
rect 111374 453922 111430 453978
rect 111498 453922 111554 453978
rect 111622 453922 111678 453978
rect 111250 436294 111306 436350
rect 111374 436294 111430 436350
rect 111498 436294 111554 436350
rect 111622 436294 111678 436350
rect 111250 436170 111306 436226
rect 111374 436170 111430 436226
rect 111498 436170 111554 436226
rect 111622 436170 111678 436226
rect 111250 436046 111306 436102
rect 111374 436046 111430 436102
rect 111498 436046 111554 436102
rect 111622 436046 111678 436102
rect 111250 435922 111306 435978
rect 111374 435922 111430 435978
rect 111498 435922 111554 435978
rect 111622 435922 111678 435978
rect 111250 418294 111306 418350
rect 111374 418294 111430 418350
rect 111498 418294 111554 418350
rect 111622 418294 111678 418350
rect 111250 418170 111306 418226
rect 111374 418170 111430 418226
rect 111498 418170 111554 418226
rect 111622 418170 111678 418226
rect 111250 418046 111306 418102
rect 111374 418046 111430 418102
rect 111498 418046 111554 418102
rect 111622 418046 111678 418102
rect 111250 417922 111306 417978
rect 111374 417922 111430 417978
rect 111498 417922 111554 417978
rect 111622 417922 111678 417978
rect 111250 400294 111306 400350
rect 111374 400294 111430 400350
rect 111498 400294 111554 400350
rect 111622 400294 111678 400350
rect 111250 400170 111306 400226
rect 111374 400170 111430 400226
rect 111498 400170 111554 400226
rect 111622 400170 111678 400226
rect 111250 400046 111306 400102
rect 111374 400046 111430 400102
rect 111498 400046 111554 400102
rect 111622 400046 111678 400102
rect 111250 399922 111306 399978
rect 111374 399922 111430 399978
rect 111498 399922 111554 399978
rect 111622 399922 111678 399978
rect 111250 382294 111306 382350
rect 111374 382294 111430 382350
rect 111498 382294 111554 382350
rect 111622 382294 111678 382350
rect 111250 382170 111306 382226
rect 111374 382170 111430 382226
rect 111498 382170 111554 382226
rect 111622 382170 111678 382226
rect 111250 382046 111306 382102
rect 111374 382046 111430 382102
rect 111498 382046 111554 382102
rect 111622 382046 111678 382102
rect 111250 381922 111306 381978
rect 111374 381922 111430 381978
rect 111498 381922 111554 381978
rect 111622 381922 111678 381978
rect 111250 364294 111306 364350
rect 111374 364294 111430 364350
rect 111498 364294 111554 364350
rect 111622 364294 111678 364350
rect 111250 364170 111306 364226
rect 111374 364170 111430 364226
rect 111498 364170 111554 364226
rect 111622 364170 111678 364226
rect 111250 364046 111306 364102
rect 111374 364046 111430 364102
rect 111498 364046 111554 364102
rect 111622 364046 111678 364102
rect 111250 363922 111306 363978
rect 111374 363922 111430 363978
rect 111498 363922 111554 363978
rect 111622 363922 111678 363978
rect 111250 346294 111306 346350
rect 111374 346294 111430 346350
rect 111498 346294 111554 346350
rect 111622 346294 111678 346350
rect 111250 346170 111306 346226
rect 111374 346170 111430 346226
rect 111498 346170 111554 346226
rect 111622 346170 111678 346226
rect 111250 346046 111306 346102
rect 111374 346046 111430 346102
rect 111498 346046 111554 346102
rect 111622 346046 111678 346102
rect 111250 345922 111306 345978
rect 111374 345922 111430 345978
rect 111498 345922 111554 345978
rect 111622 345922 111678 345978
rect 111250 328294 111306 328350
rect 111374 328294 111430 328350
rect 111498 328294 111554 328350
rect 111622 328294 111678 328350
rect 111250 328170 111306 328226
rect 111374 328170 111430 328226
rect 111498 328170 111554 328226
rect 111622 328170 111678 328226
rect 111250 328046 111306 328102
rect 111374 328046 111430 328102
rect 111498 328046 111554 328102
rect 111622 328046 111678 328102
rect 111250 327922 111306 327978
rect 111374 327922 111430 327978
rect 111498 327922 111554 327978
rect 111622 327922 111678 327978
rect 111250 310294 111306 310350
rect 111374 310294 111430 310350
rect 111498 310294 111554 310350
rect 111622 310294 111678 310350
rect 111250 310170 111306 310226
rect 111374 310170 111430 310226
rect 111498 310170 111554 310226
rect 111622 310170 111678 310226
rect 111250 310046 111306 310102
rect 111374 310046 111430 310102
rect 111498 310046 111554 310102
rect 111622 310046 111678 310102
rect 111250 309922 111306 309978
rect 111374 309922 111430 309978
rect 111498 309922 111554 309978
rect 111622 309922 111678 309978
rect 111250 292294 111306 292350
rect 111374 292294 111430 292350
rect 111498 292294 111554 292350
rect 111622 292294 111678 292350
rect 111250 292170 111306 292226
rect 111374 292170 111430 292226
rect 111498 292170 111554 292226
rect 111622 292170 111678 292226
rect 111250 292046 111306 292102
rect 111374 292046 111430 292102
rect 111498 292046 111554 292102
rect 111622 292046 111678 292102
rect 111250 291922 111306 291978
rect 111374 291922 111430 291978
rect 111498 291922 111554 291978
rect 111622 291922 111678 291978
rect 111250 274294 111306 274350
rect 111374 274294 111430 274350
rect 111498 274294 111554 274350
rect 111622 274294 111678 274350
rect 111250 274170 111306 274226
rect 111374 274170 111430 274226
rect 111498 274170 111554 274226
rect 111622 274170 111678 274226
rect 111250 274046 111306 274102
rect 111374 274046 111430 274102
rect 111498 274046 111554 274102
rect 111622 274046 111678 274102
rect 111250 273922 111306 273978
rect 111374 273922 111430 273978
rect 111498 273922 111554 273978
rect 111622 273922 111678 273978
rect 111250 256294 111306 256350
rect 111374 256294 111430 256350
rect 111498 256294 111554 256350
rect 111622 256294 111678 256350
rect 111250 256170 111306 256226
rect 111374 256170 111430 256226
rect 111498 256170 111554 256226
rect 111622 256170 111678 256226
rect 111250 256046 111306 256102
rect 111374 256046 111430 256102
rect 111498 256046 111554 256102
rect 111622 256046 111678 256102
rect 111250 255922 111306 255978
rect 111374 255922 111430 255978
rect 111498 255922 111554 255978
rect 111622 255922 111678 255978
rect 111250 238294 111306 238350
rect 111374 238294 111430 238350
rect 111498 238294 111554 238350
rect 111622 238294 111678 238350
rect 111250 238170 111306 238226
rect 111374 238170 111430 238226
rect 111498 238170 111554 238226
rect 111622 238170 111678 238226
rect 111250 238046 111306 238102
rect 111374 238046 111430 238102
rect 111498 238046 111554 238102
rect 111622 238046 111678 238102
rect 111250 237922 111306 237978
rect 111374 237922 111430 237978
rect 111498 237922 111554 237978
rect 111622 237922 111678 237978
rect 111250 220294 111306 220350
rect 111374 220294 111430 220350
rect 111498 220294 111554 220350
rect 111622 220294 111678 220350
rect 111250 220170 111306 220226
rect 111374 220170 111430 220226
rect 111498 220170 111554 220226
rect 111622 220170 111678 220226
rect 111250 220046 111306 220102
rect 111374 220046 111430 220102
rect 111498 220046 111554 220102
rect 111622 220046 111678 220102
rect 111250 219922 111306 219978
rect 111374 219922 111430 219978
rect 111498 219922 111554 219978
rect 111622 219922 111678 219978
rect 111250 202294 111306 202350
rect 111374 202294 111430 202350
rect 111498 202294 111554 202350
rect 111622 202294 111678 202350
rect 111250 202170 111306 202226
rect 111374 202170 111430 202226
rect 111498 202170 111554 202226
rect 111622 202170 111678 202226
rect 111250 202046 111306 202102
rect 111374 202046 111430 202102
rect 111498 202046 111554 202102
rect 111622 202046 111678 202102
rect 111250 201922 111306 201978
rect 111374 201922 111430 201978
rect 111498 201922 111554 201978
rect 111622 201922 111678 201978
rect 111250 184294 111306 184350
rect 111374 184294 111430 184350
rect 111498 184294 111554 184350
rect 111622 184294 111678 184350
rect 111250 184170 111306 184226
rect 111374 184170 111430 184226
rect 111498 184170 111554 184226
rect 111622 184170 111678 184226
rect 111250 184046 111306 184102
rect 111374 184046 111430 184102
rect 111498 184046 111554 184102
rect 111622 184046 111678 184102
rect 111250 183922 111306 183978
rect 111374 183922 111430 183978
rect 111498 183922 111554 183978
rect 111622 183922 111678 183978
rect 111250 166294 111306 166350
rect 111374 166294 111430 166350
rect 111498 166294 111554 166350
rect 111622 166294 111678 166350
rect 111250 166170 111306 166226
rect 111374 166170 111430 166226
rect 111498 166170 111554 166226
rect 111622 166170 111678 166226
rect 111250 166046 111306 166102
rect 111374 166046 111430 166102
rect 111498 166046 111554 166102
rect 111622 166046 111678 166102
rect 111250 165922 111306 165978
rect 111374 165922 111430 165978
rect 111498 165922 111554 165978
rect 111622 165922 111678 165978
rect 111250 148294 111306 148350
rect 111374 148294 111430 148350
rect 111498 148294 111554 148350
rect 111622 148294 111678 148350
rect 111250 148170 111306 148226
rect 111374 148170 111430 148226
rect 111498 148170 111554 148226
rect 111622 148170 111678 148226
rect 111250 148046 111306 148102
rect 111374 148046 111430 148102
rect 111498 148046 111554 148102
rect 111622 148046 111678 148102
rect 111250 147922 111306 147978
rect 111374 147922 111430 147978
rect 111498 147922 111554 147978
rect 111622 147922 111678 147978
rect 111250 130294 111306 130350
rect 111374 130294 111430 130350
rect 111498 130294 111554 130350
rect 111622 130294 111678 130350
rect 111250 130170 111306 130226
rect 111374 130170 111430 130226
rect 111498 130170 111554 130226
rect 111622 130170 111678 130226
rect 111250 130046 111306 130102
rect 111374 130046 111430 130102
rect 111498 130046 111554 130102
rect 111622 130046 111678 130102
rect 111250 129922 111306 129978
rect 111374 129922 111430 129978
rect 111498 129922 111554 129978
rect 111622 129922 111678 129978
rect 111250 112294 111306 112350
rect 111374 112294 111430 112350
rect 111498 112294 111554 112350
rect 111622 112294 111678 112350
rect 111250 112170 111306 112226
rect 111374 112170 111430 112226
rect 111498 112170 111554 112226
rect 111622 112170 111678 112226
rect 111250 112046 111306 112102
rect 111374 112046 111430 112102
rect 111498 112046 111554 112102
rect 111622 112046 111678 112102
rect 111250 111922 111306 111978
rect 111374 111922 111430 111978
rect 111498 111922 111554 111978
rect 111622 111922 111678 111978
rect 111250 94294 111306 94350
rect 111374 94294 111430 94350
rect 111498 94294 111554 94350
rect 111622 94294 111678 94350
rect 111250 94170 111306 94226
rect 111374 94170 111430 94226
rect 111498 94170 111554 94226
rect 111622 94170 111678 94226
rect 111250 94046 111306 94102
rect 111374 94046 111430 94102
rect 111498 94046 111554 94102
rect 111622 94046 111678 94102
rect 111250 93922 111306 93978
rect 111374 93922 111430 93978
rect 111498 93922 111554 93978
rect 111622 93922 111678 93978
rect 111250 76294 111306 76350
rect 111374 76294 111430 76350
rect 111498 76294 111554 76350
rect 111622 76294 111678 76350
rect 111250 76170 111306 76226
rect 111374 76170 111430 76226
rect 111498 76170 111554 76226
rect 111622 76170 111678 76226
rect 111250 76046 111306 76102
rect 111374 76046 111430 76102
rect 111498 76046 111554 76102
rect 111622 76046 111678 76102
rect 111250 75922 111306 75978
rect 111374 75922 111430 75978
rect 111498 75922 111554 75978
rect 111622 75922 111678 75978
rect 111250 58294 111306 58350
rect 111374 58294 111430 58350
rect 111498 58294 111554 58350
rect 111622 58294 111678 58350
rect 111250 58170 111306 58226
rect 111374 58170 111430 58226
rect 111498 58170 111554 58226
rect 111622 58170 111678 58226
rect 111250 58046 111306 58102
rect 111374 58046 111430 58102
rect 111498 58046 111554 58102
rect 111622 58046 111678 58102
rect 111250 57922 111306 57978
rect 111374 57922 111430 57978
rect 111498 57922 111554 57978
rect 111622 57922 111678 57978
rect 111250 40294 111306 40350
rect 111374 40294 111430 40350
rect 111498 40294 111554 40350
rect 111622 40294 111678 40350
rect 111250 40170 111306 40226
rect 111374 40170 111430 40226
rect 111498 40170 111554 40226
rect 111622 40170 111678 40226
rect 111250 40046 111306 40102
rect 111374 40046 111430 40102
rect 111498 40046 111554 40102
rect 111622 40046 111678 40102
rect 111250 39922 111306 39978
rect 111374 39922 111430 39978
rect 111498 39922 111554 39978
rect 111622 39922 111678 39978
rect 111250 22294 111306 22350
rect 111374 22294 111430 22350
rect 111498 22294 111554 22350
rect 111622 22294 111678 22350
rect 111250 22170 111306 22226
rect 111374 22170 111430 22226
rect 111498 22170 111554 22226
rect 111622 22170 111678 22226
rect 111250 22046 111306 22102
rect 111374 22046 111430 22102
rect 111498 22046 111554 22102
rect 111622 22046 111678 22102
rect 111250 21922 111306 21978
rect 111374 21922 111430 21978
rect 111498 21922 111554 21978
rect 111622 21922 111678 21978
rect 111250 4294 111306 4350
rect 111374 4294 111430 4350
rect 111498 4294 111554 4350
rect 111622 4294 111678 4350
rect 111250 4170 111306 4226
rect 111374 4170 111430 4226
rect 111498 4170 111554 4226
rect 111622 4170 111678 4226
rect 111250 4046 111306 4102
rect 111374 4046 111430 4102
rect 111498 4046 111554 4102
rect 111622 4046 111678 4102
rect 111250 3922 111306 3978
rect 111374 3922 111430 3978
rect 111498 3922 111554 3978
rect 111622 3922 111678 3978
rect 111250 -216 111306 -160
rect 111374 -216 111430 -160
rect 111498 -216 111554 -160
rect 111622 -216 111678 -160
rect 111250 -340 111306 -284
rect 111374 -340 111430 -284
rect 111498 -340 111554 -284
rect 111622 -340 111678 -284
rect 111250 -464 111306 -408
rect 111374 -464 111430 -408
rect 111498 -464 111554 -408
rect 111622 -464 111678 -408
rect 111250 -588 111306 -532
rect 111374 -588 111430 -532
rect 111498 -588 111554 -532
rect 111622 -588 111678 -532
rect 114970 598116 115026 598172
rect 115094 598116 115150 598172
rect 115218 598116 115274 598172
rect 115342 598116 115398 598172
rect 114970 597992 115026 598048
rect 115094 597992 115150 598048
rect 115218 597992 115274 598048
rect 115342 597992 115398 598048
rect 114970 597868 115026 597924
rect 115094 597868 115150 597924
rect 115218 597868 115274 597924
rect 115342 597868 115398 597924
rect 114970 597744 115026 597800
rect 115094 597744 115150 597800
rect 115218 597744 115274 597800
rect 115342 597744 115398 597800
rect 114970 586294 115026 586350
rect 115094 586294 115150 586350
rect 115218 586294 115274 586350
rect 115342 586294 115398 586350
rect 114970 586170 115026 586226
rect 115094 586170 115150 586226
rect 115218 586170 115274 586226
rect 115342 586170 115398 586226
rect 114970 586046 115026 586102
rect 115094 586046 115150 586102
rect 115218 586046 115274 586102
rect 115342 586046 115398 586102
rect 114970 585922 115026 585978
rect 115094 585922 115150 585978
rect 115218 585922 115274 585978
rect 115342 585922 115398 585978
rect 114970 568294 115026 568350
rect 115094 568294 115150 568350
rect 115218 568294 115274 568350
rect 115342 568294 115398 568350
rect 114970 568170 115026 568226
rect 115094 568170 115150 568226
rect 115218 568170 115274 568226
rect 115342 568170 115398 568226
rect 114970 568046 115026 568102
rect 115094 568046 115150 568102
rect 115218 568046 115274 568102
rect 115342 568046 115398 568102
rect 114970 567922 115026 567978
rect 115094 567922 115150 567978
rect 115218 567922 115274 567978
rect 115342 567922 115398 567978
rect 114970 550294 115026 550350
rect 115094 550294 115150 550350
rect 115218 550294 115274 550350
rect 115342 550294 115398 550350
rect 114970 550170 115026 550226
rect 115094 550170 115150 550226
rect 115218 550170 115274 550226
rect 115342 550170 115398 550226
rect 114970 550046 115026 550102
rect 115094 550046 115150 550102
rect 115218 550046 115274 550102
rect 115342 550046 115398 550102
rect 114970 549922 115026 549978
rect 115094 549922 115150 549978
rect 115218 549922 115274 549978
rect 115342 549922 115398 549978
rect 114970 532294 115026 532350
rect 115094 532294 115150 532350
rect 115218 532294 115274 532350
rect 115342 532294 115398 532350
rect 114970 532170 115026 532226
rect 115094 532170 115150 532226
rect 115218 532170 115274 532226
rect 115342 532170 115398 532226
rect 114970 532046 115026 532102
rect 115094 532046 115150 532102
rect 115218 532046 115274 532102
rect 115342 532046 115398 532102
rect 114970 531922 115026 531978
rect 115094 531922 115150 531978
rect 115218 531922 115274 531978
rect 115342 531922 115398 531978
rect 114970 514294 115026 514350
rect 115094 514294 115150 514350
rect 115218 514294 115274 514350
rect 115342 514294 115398 514350
rect 114970 514170 115026 514226
rect 115094 514170 115150 514226
rect 115218 514170 115274 514226
rect 115342 514170 115398 514226
rect 114970 514046 115026 514102
rect 115094 514046 115150 514102
rect 115218 514046 115274 514102
rect 115342 514046 115398 514102
rect 114970 513922 115026 513978
rect 115094 513922 115150 513978
rect 115218 513922 115274 513978
rect 115342 513922 115398 513978
rect 114970 496294 115026 496350
rect 115094 496294 115150 496350
rect 115218 496294 115274 496350
rect 115342 496294 115398 496350
rect 114970 496170 115026 496226
rect 115094 496170 115150 496226
rect 115218 496170 115274 496226
rect 115342 496170 115398 496226
rect 114970 496046 115026 496102
rect 115094 496046 115150 496102
rect 115218 496046 115274 496102
rect 115342 496046 115398 496102
rect 114970 495922 115026 495978
rect 115094 495922 115150 495978
rect 115218 495922 115274 495978
rect 115342 495922 115398 495978
rect 114970 478294 115026 478350
rect 115094 478294 115150 478350
rect 115218 478294 115274 478350
rect 115342 478294 115398 478350
rect 114970 478170 115026 478226
rect 115094 478170 115150 478226
rect 115218 478170 115274 478226
rect 115342 478170 115398 478226
rect 114970 478046 115026 478102
rect 115094 478046 115150 478102
rect 115218 478046 115274 478102
rect 115342 478046 115398 478102
rect 114970 477922 115026 477978
rect 115094 477922 115150 477978
rect 115218 477922 115274 477978
rect 115342 477922 115398 477978
rect 114970 460294 115026 460350
rect 115094 460294 115150 460350
rect 115218 460294 115274 460350
rect 115342 460294 115398 460350
rect 114970 460170 115026 460226
rect 115094 460170 115150 460226
rect 115218 460170 115274 460226
rect 115342 460170 115398 460226
rect 114970 460046 115026 460102
rect 115094 460046 115150 460102
rect 115218 460046 115274 460102
rect 115342 460046 115398 460102
rect 114970 459922 115026 459978
rect 115094 459922 115150 459978
rect 115218 459922 115274 459978
rect 115342 459922 115398 459978
rect 114970 442294 115026 442350
rect 115094 442294 115150 442350
rect 115218 442294 115274 442350
rect 115342 442294 115398 442350
rect 114970 442170 115026 442226
rect 115094 442170 115150 442226
rect 115218 442170 115274 442226
rect 115342 442170 115398 442226
rect 114970 442046 115026 442102
rect 115094 442046 115150 442102
rect 115218 442046 115274 442102
rect 115342 442046 115398 442102
rect 114970 441922 115026 441978
rect 115094 441922 115150 441978
rect 115218 441922 115274 441978
rect 115342 441922 115398 441978
rect 114970 424294 115026 424350
rect 115094 424294 115150 424350
rect 115218 424294 115274 424350
rect 115342 424294 115398 424350
rect 114970 424170 115026 424226
rect 115094 424170 115150 424226
rect 115218 424170 115274 424226
rect 115342 424170 115398 424226
rect 114970 424046 115026 424102
rect 115094 424046 115150 424102
rect 115218 424046 115274 424102
rect 115342 424046 115398 424102
rect 114970 423922 115026 423978
rect 115094 423922 115150 423978
rect 115218 423922 115274 423978
rect 115342 423922 115398 423978
rect 114970 406294 115026 406350
rect 115094 406294 115150 406350
rect 115218 406294 115274 406350
rect 115342 406294 115398 406350
rect 114970 406170 115026 406226
rect 115094 406170 115150 406226
rect 115218 406170 115274 406226
rect 115342 406170 115398 406226
rect 114970 406046 115026 406102
rect 115094 406046 115150 406102
rect 115218 406046 115274 406102
rect 115342 406046 115398 406102
rect 114970 405922 115026 405978
rect 115094 405922 115150 405978
rect 115218 405922 115274 405978
rect 115342 405922 115398 405978
rect 114970 388294 115026 388350
rect 115094 388294 115150 388350
rect 115218 388294 115274 388350
rect 115342 388294 115398 388350
rect 114970 388170 115026 388226
rect 115094 388170 115150 388226
rect 115218 388170 115274 388226
rect 115342 388170 115398 388226
rect 114970 388046 115026 388102
rect 115094 388046 115150 388102
rect 115218 388046 115274 388102
rect 115342 388046 115398 388102
rect 114970 387922 115026 387978
rect 115094 387922 115150 387978
rect 115218 387922 115274 387978
rect 115342 387922 115398 387978
rect 114970 370294 115026 370350
rect 115094 370294 115150 370350
rect 115218 370294 115274 370350
rect 115342 370294 115398 370350
rect 114970 370170 115026 370226
rect 115094 370170 115150 370226
rect 115218 370170 115274 370226
rect 115342 370170 115398 370226
rect 114970 370046 115026 370102
rect 115094 370046 115150 370102
rect 115218 370046 115274 370102
rect 115342 370046 115398 370102
rect 114970 369922 115026 369978
rect 115094 369922 115150 369978
rect 115218 369922 115274 369978
rect 115342 369922 115398 369978
rect 114970 352294 115026 352350
rect 115094 352294 115150 352350
rect 115218 352294 115274 352350
rect 115342 352294 115398 352350
rect 114970 352170 115026 352226
rect 115094 352170 115150 352226
rect 115218 352170 115274 352226
rect 115342 352170 115398 352226
rect 114970 352046 115026 352102
rect 115094 352046 115150 352102
rect 115218 352046 115274 352102
rect 115342 352046 115398 352102
rect 114970 351922 115026 351978
rect 115094 351922 115150 351978
rect 115218 351922 115274 351978
rect 115342 351922 115398 351978
rect 114970 334294 115026 334350
rect 115094 334294 115150 334350
rect 115218 334294 115274 334350
rect 115342 334294 115398 334350
rect 114970 334170 115026 334226
rect 115094 334170 115150 334226
rect 115218 334170 115274 334226
rect 115342 334170 115398 334226
rect 114970 334046 115026 334102
rect 115094 334046 115150 334102
rect 115218 334046 115274 334102
rect 115342 334046 115398 334102
rect 114970 333922 115026 333978
rect 115094 333922 115150 333978
rect 115218 333922 115274 333978
rect 115342 333922 115398 333978
rect 114970 316294 115026 316350
rect 115094 316294 115150 316350
rect 115218 316294 115274 316350
rect 115342 316294 115398 316350
rect 114970 316170 115026 316226
rect 115094 316170 115150 316226
rect 115218 316170 115274 316226
rect 115342 316170 115398 316226
rect 114970 316046 115026 316102
rect 115094 316046 115150 316102
rect 115218 316046 115274 316102
rect 115342 316046 115398 316102
rect 114970 315922 115026 315978
rect 115094 315922 115150 315978
rect 115218 315922 115274 315978
rect 115342 315922 115398 315978
rect 114970 298294 115026 298350
rect 115094 298294 115150 298350
rect 115218 298294 115274 298350
rect 115342 298294 115398 298350
rect 114970 298170 115026 298226
rect 115094 298170 115150 298226
rect 115218 298170 115274 298226
rect 115342 298170 115398 298226
rect 114970 298046 115026 298102
rect 115094 298046 115150 298102
rect 115218 298046 115274 298102
rect 115342 298046 115398 298102
rect 114970 297922 115026 297978
rect 115094 297922 115150 297978
rect 115218 297922 115274 297978
rect 115342 297922 115398 297978
rect 114970 280294 115026 280350
rect 115094 280294 115150 280350
rect 115218 280294 115274 280350
rect 115342 280294 115398 280350
rect 114970 280170 115026 280226
rect 115094 280170 115150 280226
rect 115218 280170 115274 280226
rect 115342 280170 115398 280226
rect 114970 280046 115026 280102
rect 115094 280046 115150 280102
rect 115218 280046 115274 280102
rect 115342 280046 115398 280102
rect 114970 279922 115026 279978
rect 115094 279922 115150 279978
rect 115218 279922 115274 279978
rect 115342 279922 115398 279978
rect 114970 262294 115026 262350
rect 115094 262294 115150 262350
rect 115218 262294 115274 262350
rect 115342 262294 115398 262350
rect 114970 262170 115026 262226
rect 115094 262170 115150 262226
rect 115218 262170 115274 262226
rect 115342 262170 115398 262226
rect 114970 262046 115026 262102
rect 115094 262046 115150 262102
rect 115218 262046 115274 262102
rect 115342 262046 115398 262102
rect 114970 261922 115026 261978
rect 115094 261922 115150 261978
rect 115218 261922 115274 261978
rect 115342 261922 115398 261978
rect 114970 244294 115026 244350
rect 115094 244294 115150 244350
rect 115218 244294 115274 244350
rect 115342 244294 115398 244350
rect 114970 244170 115026 244226
rect 115094 244170 115150 244226
rect 115218 244170 115274 244226
rect 115342 244170 115398 244226
rect 114970 244046 115026 244102
rect 115094 244046 115150 244102
rect 115218 244046 115274 244102
rect 115342 244046 115398 244102
rect 114970 243922 115026 243978
rect 115094 243922 115150 243978
rect 115218 243922 115274 243978
rect 115342 243922 115398 243978
rect 114970 226294 115026 226350
rect 115094 226294 115150 226350
rect 115218 226294 115274 226350
rect 115342 226294 115398 226350
rect 114970 226170 115026 226226
rect 115094 226170 115150 226226
rect 115218 226170 115274 226226
rect 115342 226170 115398 226226
rect 114970 226046 115026 226102
rect 115094 226046 115150 226102
rect 115218 226046 115274 226102
rect 115342 226046 115398 226102
rect 114970 225922 115026 225978
rect 115094 225922 115150 225978
rect 115218 225922 115274 225978
rect 115342 225922 115398 225978
rect 114970 208294 115026 208350
rect 115094 208294 115150 208350
rect 115218 208294 115274 208350
rect 115342 208294 115398 208350
rect 114970 208170 115026 208226
rect 115094 208170 115150 208226
rect 115218 208170 115274 208226
rect 115342 208170 115398 208226
rect 114970 208046 115026 208102
rect 115094 208046 115150 208102
rect 115218 208046 115274 208102
rect 115342 208046 115398 208102
rect 114970 207922 115026 207978
rect 115094 207922 115150 207978
rect 115218 207922 115274 207978
rect 115342 207922 115398 207978
rect 114970 190294 115026 190350
rect 115094 190294 115150 190350
rect 115218 190294 115274 190350
rect 115342 190294 115398 190350
rect 114970 190170 115026 190226
rect 115094 190170 115150 190226
rect 115218 190170 115274 190226
rect 115342 190170 115398 190226
rect 114970 190046 115026 190102
rect 115094 190046 115150 190102
rect 115218 190046 115274 190102
rect 115342 190046 115398 190102
rect 114970 189922 115026 189978
rect 115094 189922 115150 189978
rect 115218 189922 115274 189978
rect 115342 189922 115398 189978
rect 114970 172294 115026 172350
rect 115094 172294 115150 172350
rect 115218 172294 115274 172350
rect 115342 172294 115398 172350
rect 114970 172170 115026 172226
rect 115094 172170 115150 172226
rect 115218 172170 115274 172226
rect 115342 172170 115398 172226
rect 114970 172046 115026 172102
rect 115094 172046 115150 172102
rect 115218 172046 115274 172102
rect 115342 172046 115398 172102
rect 114970 171922 115026 171978
rect 115094 171922 115150 171978
rect 115218 171922 115274 171978
rect 115342 171922 115398 171978
rect 114970 154294 115026 154350
rect 115094 154294 115150 154350
rect 115218 154294 115274 154350
rect 115342 154294 115398 154350
rect 114970 154170 115026 154226
rect 115094 154170 115150 154226
rect 115218 154170 115274 154226
rect 115342 154170 115398 154226
rect 114970 154046 115026 154102
rect 115094 154046 115150 154102
rect 115218 154046 115274 154102
rect 115342 154046 115398 154102
rect 114970 153922 115026 153978
rect 115094 153922 115150 153978
rect 115218 153922 115274 153978
rect 115342 153922 115398 153978
rect 114970 136294 115026 136350
rect 115094 136294 115150 136350
rect 115218 136294 115274 136350
rect 115342 136294 115398 136350
rect 114970 136170 115026 136226
rect 115094 136170 115150 136226
rect 115218 136170 115274 136226
rect 115342 136170 115398 136226
rect 114970 136046 115026 136102
rect 115094 136046 115150 136102
rect 115218 136046 115274 136102
rect 115342 136046 115398 136102
rect 114970 135922 115026 135978
rect 115094 135922 115150 135978
rect 115218 135922 115274 135978
rect 115342 135922 115398 135978
rect 114970 118294 115026 118350
rect 115094 118294 115150 118350
rect 115218 118294 115274 118350
rect 115342 118294 115398 118350
rect 114970 118170 115026 118226
rect 115094 118170 115150 118226
rect 115218 118170 115274 118226
rect 115342 118170 115398 118226
rect 114970 118046 115026 118102
rect 115094 118046 115150 118102
rect 115218 118046 115274 118102
rect 115342 118046 115398 118102
rect 114970 117922 115026 117978
rect 115094 117922 115150 117978
rect 115218 117922 115274 117978
rect 115342 117922 115398 117978
rect 114970 100294 115026 100350
rect 115094 100294 115150 100350
rect 115218 100294 115274 100350
rect 115342 100294 115398 100350
rect 114970 100170 115026 100226
rect 115094 100170 115150 100226
rect 115218 100170 115274 100226
rect 115342 100170 115398 100226
rect 114970 100046 115026 100102
rect 115094 100046 115150 100102
rect 115218 100046 115274 100102
rect 115342 100046 115398 100102
rect 114970 99922 115026 99978
rect 115094 99922 115150 99978
rect 115218 99922 115274 99978
rect 115342 99922 115398 99978
rect 114970 82294 115026 82350
rect 115094 82294 115150 82350
rect 115218 82294 115274 82350
rect 115342 82294 115398 82350
rect 114970 82170 115026 82226
rect 115094 82170 115150 82226
rect 115218 82170 115274 82226
rect 115342 82170 115398 82226
rect 114970 82046 115026 82102
rect 115094 82046 115150 82102
rect 115218 82046 115274 82102
rect 115342 82046 115398 82102
rect 114970 81922 115026 81978
rect 115094 81922 115150 81978
rect 115218 81922 115274 81978
rect 115342 81922 115398 81978
rect 114970 64294 115026 64350
rect 115094 64294 115150 64350
rect 115218 64294 115274 64350
rect 115342 64294 115398 64350
rect 114970 64170 115026 64226
rect 115094 64170 115150 64226
rect 115218 64170 115274 64226
rect 115342 64170 115398 64226
rect 114970 64046 115026 64102
rect 115094 64046 115150 64102
rect 115218 64046 115274 64102
rect 115342 64046 115398 64102
rect 114970 63922 115026 63978
rect 115094 63922 115150 63978
rect 115218 63922 115274 63978
rect 115342 63922 115398 63978
rect 114970 46294 115026 46350
rect 115094 46294 115150 46350
rect 115218 46294 115274 46350
rect 115342 46294 115398 46350
rect 114970 46170 115026 46226
rect 115094 46170 115150 46226
rect 115218 46170 115274 46226
rect 115342 46170 115398 46226
rect 114970 46046 115026 46102
rect 115094 46046 115150 46102
rect 115218 46046 115274 46102
rect 115342 46046 115398 46102
rect 114970 45922 115026 45978
rect 115094 45922 115150 45978
rect 115218 45922 115274 45978
rect 115342 45922 115398 45978
rect 114970 28294 115026 28350
rect 115094 28294 115150 28350
rect 115218 28294 115274 28350
rect 115342 28294 115398 28350
rect 114970 28170 115026 28226
rect 115094 28170 115150 28226
rect 115218 28170 115274 28226
rect 115342 28170 115398 28226
rect 114970 28046 115026 28102
rect 115094 28046 115150 28102
rect 115218 28046 115274 28102
rect 115342 28046 115398 28102
rect 114970 27922 115026 27978
rect 115094 27922 115150 27978
rect 115218 27922 115274 27978
rect 115342 27922 115398 27978
rect 114970 10294 115026 10350
rect 115094 10294 115150 10350
rect 115218 10294 115274 10350
rect 115342 10294 115398 10350
rect 114970 10170 115026 10226
rect 115094 10170 115150 10226
rect 115218 10170 115274 10226
rect 115342 10170 115398 10226
rect 114970 10046 115026 10102
rect 115094 10046 115150 10102
rect 115218 10046 115274 10102
rect 115342 10046 115398 10102
rect 114970 9922 115026 9978
rect 115094 9922 115150 9978
rect 115218 9922 115274 9978
rect 115342 9922 115398 9978
rect 114970 -1176 115026 -1120
rect 115094 -1176 115150 -1120
rect 115218 -1176 115274 -1120
rect 115342 -1176 115398 -1120
rect 114970 -1300 115026 -1244
rect 115094 -1300 115150 -1244
rect 115218 -1300 115274 -1244
rect 115342 -1300 115398 -1244
rect 114970 -1424 115026 -1368
rect 115094 -1424 115150 -1368
rect 115218 -1424 115274 -1368
rect 115342 -1424 115398 -1368
rect 114970 -1548 115026 -1492
rect 115094 -1548 115150 -1492
rect 115218 -1548 115274 -1492
rect 115342 -1548 115398 -1492
rect 129250 597156 129306 597212
rect 129374 597156 129430 597212
rect 129498 597156 129554 597212
rect 129622 597156 129678 597212
rect 129250 597032 129306 597088
rect 129374 597032 129430 597088
rect 129498 597032 129554 597088
rect 129622 597032 129678 597088
rect 129250 596908 129306 596964
rect 129374 596908 129430 596964
rect 129498 596908 129554 596964
rect 129622 596908 129678 596964
rect 129250 596784 129306 596840
rect 129374 596784 129430 596840
rect 129498 596784 129554 596840
rect 129622 596784 129678 596840
rect 129250 580294 129306 580350
rect 129374 580294 129430 580350
rect 129498 580294 129554 580350
rect 129622 580294 129678 580350
rect 129250 580170 129306 580226
rect 129374 580170 129430 580226
rect 129498 580170 129554 580226
rect 129622 580170 129678 580226
rect 129250 580046 129306 580102
rect 129374 580046 129430 580102
rect 129498 580046 129554 580102
rect 129622 580046 129678 580102
rect 129250 579922 129306 579978
rect 129374 579922 129430 579978
rect 129498 579922 129554 579978
rect 129622 579922 129678 579978
rect 129250 562294 129306 562350
rect 129374 562294 129430 562350
rect 129498 562294 129554 562350
rect 129622 562294 129678 562350
rect 129250 562170 129306 562226
rect 129374 562170 129430 562226
rect 129498 562170 129554 562226
rect 129622 562170 129678 562226
rect 129250 562046 129306 562102
rect 129374 562046 129430 562102
rect 129498 562046 129554 562102
rect 129622 562046 129678 562102
rect 129250 561922 129306 561978
rect 129374 561922 129430 561978
rect 129498 561922 129554 561978
rect 129622 561922 129678 561978
rect 129250 544294 129306 544350
rect 129374 544294 129430 544350
rect 129498 544294 129554 544350
rect 129622 544294 129678 544350
rect 129250 544170 129306 544226
rect 129374 544170 129430 544226
rect 129498 544170 129554 544226
rect 129622 544170 129678 544226
rect 129250 544046 129306 544102
rect 129374 544046 129430 544102
rect 129498 544046 129554 544102
rect 129622 544046 129678 544102
rect 129250 543922 129306 543978
rect 129374 543922 129430 543978
rect 129498 543922 129554 543978
rect 129622 543922 129678 543978
rect 129250 526294 129306 526350
rect 129374 526294 129430 526350
rect 129498 526294 129554 526350
rect 129622 526294 129678 526350
rect 129250 526170 129306 526226
rect 129374 526170 129430 526226
rect 129498 526170 129554 526226
rect 129622 526170 129678 526226
rect 129250 526046 129306 526102
rect 129374 526046 129430 526102
rect 129498 526046 129554 526102
rect 129622 526046 129678 526102
rect 129250 525922 129306 525978
rect 129374 525922 129430 525978
rect 129498 525922 129554 525978
rect 129622 525922 129678 525978
rect 129250 508294 129306 508350
rect 129374 508294 129430 508350
rect 129498 508294 129554 508350
rect 129622 508294 129678 508350
rect 129250 508170 129306 508226
rect 129374 508170 129430 508226
rect 129498 508170 129554 508226
rect 129622 508170 129678 508226
rect 129250 508046 129306 508102
rect 129374 508046 129430 508102
rect 129498 508046 129554 508102
rect 129622 508046 129678 508102
rect 129250 507922 129306 507978
rect 129374 507922 129430 507978
rect 129498 507922 129554 507978
rect 129622 507922 129678 507978
rect 129250 490294 129306 490350
rect 129374 490294 129430 490350
rect 129498 490294 129554 490350
rect 129622 490294 129678 490350
rect 129250 490170 129306 490226
rect 129374 490170 129430 490226
rect 129498 490170 129554 490226
rect 129622 490170 129678 490226
rect 129250 490046 129306 490102
rect 129374 490046 129430 490102
rect 129498 490046 129554 490102
rect 129622 490046 129678 490102
rect 129250 489922 129306 489978
rect 129374 489922 129430 489978
rect 129498 489922 129554 489978
rect 129622 489922 129678 489978
rect 129250 472294 129306 472350
rect 129374 472294 129430 472350
rect 129498 472294 129554 472350
rect 129622 472294 129678 472350
rect 129250 472170 129306 472226
rect 129374 472170 129430 472226
rect 129498 472170 129554 472226
rect 129622 472170 129678 472226
rect 129250 472046 129306 472102
rect 129374 472046 129430 472102
rect 129498 472046 129554 472102
rect 129622 472046 129678 472102
rect 129250 471922 129306 471978
rect 129374 471922 129430 471978
rect 129498 471922 129554 471978
rect 129622 471922 129678 471978
rect 129250 454294 129306 454350
rect 129374 454294 129430 454350
rect 129498 454294 129554 454350
rect 129622 454294 129678 454350
rect 129250 454170 129306 454226
rect 129374 454170 129430 454226
rect 129498 454170 129554 454226
rect 129622 454170 129678 454226
rect 129250 454046 129306 454102
rect 129374 454046 129430 454102
rect 129498 454046 129554 454102
rect 129622 454046 129678 454102
rect 129250 453922 129306 453978
rect 129374 453922 129430 453978
rect 129498 453922 129554 453978
rect 129622 453922 129678 453978
rect 129250 436294 129306 436350
rect 129374 436294 129430 436350
rect 129498 436294 129554 436350
rect 129622 436294 129678 436350
rect 129250 436170 129306 436226
rect 129374 436170 129430 436226
rect 129498 436170 129554 436226
rect 129622 436170 129678 436226
rect 129250 436046 129306 436102
rect 129374 436046 129430 436102
rect 129498 436046 129554 436102
rect 129622 436046 129678 436102
rect 129250 435922 129306 435978
rect 129374 435922 129430 435978
rect 129498 435922 129554 435978
rect 129622 435922 129678 435978
rect 129250 418294 129306 418350
rect 129374 418294 129430 418350
rect 129498 418294 129554 418350
rect 129622 418294 129678 418350
rect 129250 418170 129306 418226
rect 129374 418170 129430 418226
rect 129498 418170 129554 418226
rect 129622 418170 129678 418226
rect 129250 418046 129306 418102
rect 129374 418046 129430 418102
rect 129498 418046 129554 418102
rect 129622 418046 129678 418102
rect 129250 417922 129306 417978
rect 129374 417922 129430 417978
rect 129498 417922 129554 417978
rect 129622 417922 129678 417978
rect 129250 400294 129306 400350
rect 129374 400294 129430 400350
rect 129498 400294 129554 400350
rect 129622 400294 129678 400350
rect 129250 400170 129306 400226
rect 129374 400170 129430 400226
rect 129498 400170 129554 400226
rect 129622 400170 129678 400226
rect 129250 400046 129306 400102
rect 129374 400046 129430 400102
rect 129498 400046 129554 400102
rect 129622 400046 129678 400102
rect 129250 399922 129306 399978
rect 129374 399922 129430 399978
rect 129498 399922 129554 399978
rect 129622 399922 129678 399978
rect 129250 382294 129306 382350
rect 129374 382294 129430 382350
rect 129498 382294 129554 382350
rect 129622 382294 129678 382350
rect 129250 382170 129306 382226
rect 129374 382170 129430 382226
rect 129498 382170 129554 382226
rect 129622 382170 129678 382226
rect 129250 382046 129306 382102
rect 129374 382046 129430 382102
rect 129498 382046 129554 382102
rect 129622 382046 129678 382102
rect 129250 381922 129306 381978
rect 129374 381922 129430 381978
rect 129498 381922 129554 381978
rect 129622 381922 129678 381978
rect 129250 364294 129306 364350
rect 129374 364294 129430 364350
rect 129498 364294 129554 364350
rect 129622 364294 129678 364350
rect 129250 364170 129306 364226
rect 129374 364170 129430 364226
rect 129498 364170 129554 364226
rect 129622 364170 129678 364226
rect 129250 364046 129306 364102
rect 129374 364046 129430 364102
rect 129498 364046 129554 364102
rect 129622 364046 129678 364102
rect 129250 363922 129306 363978
rect 129374 363922 129430 363978
rect 129498 363922 129554 363978
rect 129622 363922 129678 363978
rect 129250 346294 129306 346350
rect 129374 346294 129430 346350
rect 129498 346294 129554 346350
rect 129622 346294 129678 346350
rect 129250 346170 129306 346226
rect 129374 346170 129430 346226
rect 129498 346170 129554 346226
rect 129622 346170 129678 346226
rect 129250 346046 129306 346102
rect 129374 346046 129430 346102
rect 129498 346046 129554 346102
rect 129622 346046 129678 346102
rect 129250 345922 129306 345978
rect 129374 345922 129430 345978
rect 129498 345922 129554 345978
rect 129622 345922 129678 345978
rect 129250 328294 129306 328350
rect 129374 328294 129430 328350
rect 129498 328294 129554 328350
rect 129622 328294 129678 328350
rect 129250 328170 129306 328226
rect 129374 328170 129430 328226
rect 129498 328170 129554 328226
rect 129622 328170 129678 328226
rect 129250 328046 129306 328102
rect 129374 328046 129430 328102
rect 129498 328046 129554 328102
rect 129622 328046 129678 328102
rect 129250 327922 129306 327978
rect 129374 327922 129430 327978
rect 129498 327922 129554 327978
rect 129622 327922 129678 327978
rect 129250 310294 129306 310350
rect 129374 310294 129430 310350
rect 129498 310294 129554 310350
rect 129622 310294 129678 310350
rect 129250 310170 129306 310226
rect 129374 310170 129430 310226
rect 129498 310170 129554 310226
rect 129622 310170 129678 310226
rect 129250 310046 129306 310102
rect 129374 310046 129430 310102
rect 129498 310046 129554 310102
rect 129622 310046 129678 310102
rect 129250 309922 129306 309978
rect 129374 309922 129430 309978
rect 129498 309922 129554 309978
rect 129622 309922 129678 309978
rect 129250 292294 129306 292350
rect 129374 292294 129430 292350
rect 129498 292294 129554 292350
rect 129622 292294 129678 292350
rect 129250 292170 129306 292226
rect 129374 292170 129430 292226
rect 129498 292170 129554 292226
rect 129622 292170 129678 292226
rect 129250 292046 129306 292102
rect 129374 292046 129430 292102
rect 129498 292046 129554 292102
rect 129622 292046 129678 292102
rect 129250 291922 129306 291978
rect 129374 291922 129430 291978
rect 129498 291922 129554 291978
rect 129622 291922 129678 291978
rect 129250 274294 129306 274350
rect 129374 274294 129430 274350
rect 129498 274294 129554 274350
rect 129622 274294 129678 274350
rect 129250 274170 129306 274226
rect 129374 274170 129430 274226
rect 129498 274170 129554 274226
rect 129622 274170 129678 274226
rect 129250 274046 129306 274102
rect 129374 274046 129430 274102
rect 129498 274046 129554 274102
rect 129622 274046 129678 274102
rect 129250 273922 129306 273978
rect 129374 273922 129430 273978
rect 129498 273922 129554 273978
rect 129622 273922 129678 273978
rect 129250 256294 129306 256350
rect 129374 256294 129430 256350
rect 129498 256294 129554 256350
rect 129622 256294 129678 256350
rect 129250 256170 129306 256226
rect 129374 256170 129430 256226
rect 129498 256170 129554 256226
rect 129622 256170 129678 256226
rect 129250 256046 129306 256102
rect 129374 256046 129430 256102
rect 129498 256046 129554 256102
rect 129622 256046 129678 256102
rect 129250 255922 129306 255978
rect 129374 255922 129430 255978
rect 129498 255922 129554 255978
rect 129622 255922 129678 255978
rect 129250 238294 129306 238350
rect 129374 238294 129430 238350
rect 129498 238294 129554 238350
rect 129622 238294 129678 238350
rect 129250 238170 129306 238226
rect 129374 238170 129430 238226
rect 129498 238170 129554 238226
rect 129622 238170 129678 238226
rect 129250 238046 129306 238102
rect 129374 238046 129430 238102
rect 129498 238046 129554 238102
rect 129622 238046 129678 238102
rect 129250 237922 129306 237978
rect 129374 237922 129430 237978
rect 129498 237922 129554 237978
rect 129622 237922 129678 237978
rect 129250 220294 129306 220350
rect 129374 220294 129430 220350
rect 129498 220294 129554 220350
rect 129622 220294 129678 220350
rect 129250 220170 129306 220226
rect 129374 220170 129430 220226
rect 129498 220170 129554 220226
rect 129622 220170 129678 220226
rect 129250 220046 129306 220102
rect 129374 220046 129430 220102
rect 129498 220046 129554 220102
rect 129622 220046 129678 220102
rect 129250 219922 129306 219978
rect 129374 219922 129430 219978
rect 129498 219922 129554 219978
rect 129622 219922 129678 219978
rect 129250 202294 129306 202350
rect 129374 202294 129430 202350
rect 129498 202294 129554 202350
rect 129622 202294 129678 202350
rect 129250 202170 129306 202226
rect 129374 202170 129430 202226
rect 129498 202170 129554 202226
rect 129622 202170 129678 202226
rect 129250 202046 129306 202102
rect 129374 202046 129430 202102
rect 129498 202046 129554 202102
rect 129622 202046 129678 202102
rect 129250 201922 129306 201978
rect 129374 201922 129430 201978
rect 129498 201922 129554 201978
rect 129622 201922 129678 201978
rect 129250 184294 129306 184350
rect 129374 184294 129430 184350
rect 129498 184294 129554 184350
rect 129622 184294 129678 184350
rect 129250 184170 129306 184226
rect 129374 184170 129430 184226
rect 129498 184170 129554 184226
rect 129622 184170 129678 184226
rect 129250 184046 129306 184102
rect 129374 184046 129430 184102
rect 129498 184046 129554 184102
rect 129622 184046 129678 184102
rect 129250 183922 129306 183978
rect 129374 183922 129430 183978
rect 129498 183922 129554 183978
rect 129622 183922 129678 183978
rect 129250 166294 129306 166350
rect 129374 166294 129430 166350
rect 129498 166294 129554 166350
rect 129622 166294 129678 166350
rect 129250 166170 129306 166226
rect 129374 166170 129430 166226
rect 129498 166170 129554 166226
rect 129622 166170 129678 166226
rect 129250 166046 129306 166102
rect 129374 166046 129430 166102
rect 129498 166046 129554 166102
rect 129622 166046 129678 166102
rect 129250 165922 129306 165978
rect 129374 165922 129430 165978
rect 129498 165922 129554 165978
rect 129622 165922 129678 165978
rect 129250 148294 129306 148350
rect 129374 148294 129430 148350
rect 129498 148294 129554 148350
rect 129622 148294 129678 148350
rect 129250 148170 129306 148226
rect 129374 148170 129430 148226
rect 129498 148170 129554 148226
rect 129622 148170 129678 148226
rect 129250 148046 129306 148102
rect 129374 148046 129430 148102
rect 129498 148046 129554 148102
rect 129622 148046 129678 148102
rect 129250 147922 129306 147978
rect 129374 147922 129430 147978
rect 129498 147922 129554 147978
rect 129622 147922 129678 147978
rect 129250 130294 129306 130350
rect 129374 130294 129430 130350
rect 129498 130294 129554 130350
rect 129622 130294 129678 130350
rect 129250 130170 129306 130226
rect 129374 130170 129430 130226
rect 129498 130170 129554 130226
rect 129622 130170 129678 130226
rect 129250 130046 129306 130102
rect 129374 130046 129430 130102
rect 129498 130046 129554 130102
rect 129622 130046 129678 130102
rect 129250 129922 129306 129978
rect 129374 129922 129430 129978
rect 129498 129922 129554 129978
rect 129622 129922 129678 129978
rect 129250 112294 129306 112350
rect 129374 112294 129430 112350
rect 129498 112294 129554 112350
rect 129622 112294 129678 112350
rect 129250 112170 129306 112226
rect 129374 112170 129430 112226
rect 129498 112170 129554 112226
rect 129622 112170 129678 112226
rect 129250 112046 129306 112102
rect 129374 112046 129430 112102
rect 129498 112046 129554 112102
rect 129622 112046 129678 112102
rect 129250 111922 129306 111978
rect 129374 111922 129430 111978
rect 129498 111922 129554 111978
rect 129622 111922 129678 111978
rect 129250 94294 129306 94350
rect 129374 94294 129430 94350
rect 129498 94294 129554 94350
rect 129622 94294 129678 94350
rect 129250 94170 129306 94226
rect 129374 94170 129430 94226
rect 129498 94170 129554 94226
rect 129622 94170 129678 94226
rect 129250 94046 129306 94102
rect 129374 94046 129430 94102
rect 129498 94046 129554 94102
rect 129622 94046 129678 94102
rect 129250 93922 129306 93978
rect 129374 93922 129430 93978
rect 129498 93922 129554 93978
rect 129622 93922 129678 93978
rect 129250 76294 129306 76350
rect 129374 76294 129430 76350
rect 129498 76294 129554 76350
rect 129622 76294 129678 76350
rect 129250 76170 129306 76226
rect 129374 76170 129430 76226
rect 129498 76170 129554 76226
rect 129622 76170 129678 76226
rect 129250 76046 129306 76102
rect 129374 76046 129430 76102
rect 129498 76046 129554 76102
rect 129622 76046 129678 76102
rect 129250 75922 129306 75978
rect 129374 75922 129430 75978
rect 129498 75922 129554 75978
rect 129622 75922 129678 75978
rect 129250 58294 129306 58350
rect 129374 58294 129430 58350
rect 129498 58294 129554 58350
rect 129622 58294 129678 58350
rect 129250 58170 129306 58226
rect 129374 58170 129430 58226
rect 129498 58170 129554 58226
rect 129622 58170 129678 58226
rect 129250 58046 129306 58102
rect 129374 58046 129430 58102
rect 129498 58046 129554 58102
rect 129622 58046 129678 58102
rect 129250 57922 129306 57978
rect 129374 57922 129430 57978
rect 129498 57922 129554 57978
rect 129622 57922 129678 57978
rect 129250 40294 129306 40350
rect 129374 40294 129430 40350
rect 129498 40294 129554 40350
rect 129622 40294 129678 40350
rect 129250 40170 129306 40226
rect 129374 40170 129430 40226
rect 129498 40170 129554 40226
rect 129622 40170 129678 40226
rect 129250 40046 129306 40102
rect 129374 40046 129430 40102
rect 129498 40046 129554 40102
rect 129622 40046 129678 40102
rect 129250 39922 129306 39978
rect 129374 39922 129430 39978
rect 129498 39922 129554 39978
rect 129622 39922 129678 39978
rect 129250 22294 129306 22350
rect 129374 22294 129430 22350
rect 129498 22294 129554 22350
rect 129622 22294 129678 22350
rect 129250 22170 129306 22226
rect 129374 22170 129430 22226
rect 129498 22170 129554 22226
rect 129622 22170 129678 22226
rect 129250 22046 129306 22102
rect 129374 22046 129430 22102
rect 129498 22046 129554 22102
rect 129622 22046 129678 22102
rect 129250 21922 129306 21978
rect 129374 21922 129430 21978
rect 129498 21922 129554 21978
rect 129622 21922 129678 21978
rect 129250 4294 129306 4350
rect 129374 4294 129430 4350
rect 129498 4294 129554 4350
rect 129622 4294 129678 4350
rect 129250 4170 129306 4226
rect 129374 4170 129430 4226
rect 129498 4170 129554 4226
rect 129622 4170 129678 4226
rect 129250 4046 129306 4102
rect 129374 4046 129430 4102
rect 129498 4046 129554 4102
rect 129622 4046 129678 4102
rect 129250 3922 129306 3978
rect 129374 3922 129430 3978
rect 129498 3922 129554 3978
rect 129622 3922 129678 3978
rect 129250 -216 129306 -160
rect 129374 -216 129430 -160
rect 129498 -216 129554 -160
rect 129622 -216 129678 -160
rect 129250 -340 129306 -284
rect 129374 -340 129430 -284
rect 129498 -340 129554 -284
rect 129622 -340 129678 -284
rect 129250 -464 129306 -408
rect 129374 -464 129430 -408
rect 129498 -464 129554 -408
rect 129622 -464 129678 -408
rect 129250 -588 129306 -532
rect 129374 -588 129430 -532
rect 129498 -588 129554 -532
rect 129622 -588 129678 -532
rect 132970 598116 133026 598172
rect 133094 598116 133150 598172
rect 133218 598116 133274 598172
rect 133342 598116 133398 598172
rect 132970 597992 133026 598048
rect 133094 597992 133150 598048
rect 133218 597992 133274 598048
rect 133342 597992 133398 598048
rect 132970 597868 133026 597924
rect 133094 597868 133150 597924
rect 133218 597868 133274 597924
rect 133342 597868 133398 597924
rect 132970 597744 133026 597800
rect 133094 597744 133150 597800
rect 133218 597744 133274 597800
rect 133342 597744 133398 597800
rect 132970 586294 133026 586350
rect 133094 586294 133150 586350
rect 133218 586294 133274 586350
rect 133342 586294 133398 586350
rect 132970 586170 133026 586226
rect 133094 586170 133150 586226
rect 133218 586170 133274 586226
rect 133342 586170 133398 586226
rect 132970 586046 133026 586102
rect 133094 586046 133150 586102
rect 133218 586046 133274 586102
rect 133342 586046 133398 586102
rect 132970 585922 133026 585978
rect 133094 585922 133150 585978
rect 133218 585922 133274 585978
rect 133342 585922 133398 585978
rect 132970 568294 133026 568350
rect 133094 568294 133150 568350
rect 133218 568294 133274 568350
rect 133342 568294 133398 568350
rect 132970 568170 133026 568226
rect 133094 568170 133150 568226
rect 133218 568170 133274 568226
rect 133342 568170 133398 568226
rect 132970 568046 133026 568102
rect 133094 568046 133150 568102
rect 133218 568046 133274 568102
rect 133342 568046 133398 568102
rect 132970 567922 133026 567978
rect 133094 567922 133150 567978
rect 133218 567922 133274 567978
rect 133342 567922 133398 567978
rect 132970 550294 133026 550350
rect 133094 550294 133150 550350
rect 133218 550294 133274 550350
rect 133342 550294 133398 550350
rect 132970 550170 133026 550226
rect 133094 550170 133150 550226
rect 133218 550170 133274 550226
rect 133342 550170 133398 550226
rect 132970 550046 133026 550102
rect 133094 550046 133150 550102
rect 133218 550046 133274 550102
rect 133342 550046 133398 550102
rect 132970 549922 133026 549978
rect 133094 549922 133150 549978
rect 133218 549922 133274 549978
rect 133342 549922 133398 549978
rect 132970 532294 133026 532350
rect 133094 532294 133150 532350
rect 133218 532294 133274 532350
rect 133342 532294 133398 532350
rect 132970 532170 133026 532226
rect 133094 532170 133150 532226
rect 133218 532170 133274 532226
rect 133342 532170 133398 532226
rect 132970 532046 133026 532102
rect 133094 532046 133150 532102
rect 133218 532046 133274 532102
rect 133342 532046 133398 532102
rect 132970 531922 133026 531978
rect 133094 531922 133150 531978
rect 133218 531922 133274 531978
rect 133342 531922 133398 531978
rect 132970 514294 133026 514350
rect 133094 514294 133150 514350
rect 133218 514294 133274 514350
rect 133342 514294 133398 514350
rect 132970 514170 133026 514226
rect 133094 514170 133150 514226
rect 133218 514170 133274 514226
rect 133342 514170 133398 514226
rect 132970 514046 133026 514102
rect 133094 514046 133150 514102
rect 133218 514046 133274 514102
rect 133342 514046 133398 514102
rect 132970 513922 133026 513978
rect 133094 513922 133150 513978
rect 133218 513922 133274 513978
rect 133342 513922 133398 513978
rect 132970 496294 133026 496350
rect 133094 496294 133150 496350
rect 133218 496294 133274 496350
rect 133342 496294 133398 496350
rect 132970 496170 133026 496226
rect 133094 496170 133150 496226
rect 133218 496170 133274 496226
rect 133342 496170 133398 496226
rect 132970 496046 133026 496102
rect 133094 496046 133150 496102
rect 133218 496046 133274 496102
rect 133342 496046 133398 496102
rect 132970 495922 133026 495978
rect 133094 495922 133150 495978
rect 133218 495922 133274 495978
rect 133342 495922 133398 495978
rect 132970 478294 133026 478350
rect 133094 478294 133150 478350
rect 133218 478294 133274 478350
rect 133342 478294 133398 478350
rect 132970 478170 133026 478226
rect 133094 478170 133150 478226
rect 133218 478170 133274 478226
rect 133342 478170 133398 478226
rect 132970 478046 133026 478102
rect 133094 478046 133150 478102
rect 133218 478046 133274 478102
rect 133342 478046 133398 478102
rect 132970 477922 133026 477978
rect 133094 477922 133150 477978
rect 133218 477922 133274 477978
rect 133342 477922 133398 477978
rect 132970 460294 133026 460350
rect 133094 460294 133150 460350
rect 133218 460294 133274 460350
rect 133342 460294 133398 460350
rect 132970 460170 133026 460226
rect 133094 460170 133150 460226
rect 133218 460170 133274 460226
rect 133342 460170 133398 460226
rect 132970 460046 133026 460102
rect 133094 460046 133150 460102
rect 133218 460046 133274 460102
rect 133342 460046 133398 460102
rect 132970 459922 133026 459978
rect 133094 459922 133150 459978
rect 133218 459922 133274 459978
rect 133342 459922 133398 459978
rect 132970 442294 133026 442350
rect 133094 442294 133150 442350
rect 133218 442294 133274 442350
rect 133342 442294 133398 442350
rect 132970 442170 133026 442226
rect 133094 442170 133150 442226
rect 133218 442170 133274 442226
rect 133342 442170 133398 442226
rect 132970 442046 133026 442102
rect 133094 442046 133150 442102
rect 133218 442046 133274 442102
rect 133342 442046 133398 442102
rect 132970 441922 133026 441978
rect 133094 441922 133150 441978
rect 133218 441922 133274 441978
rect 133342 441922 133398 441978
rect 132970 424294 133026 424350
rect 133094 424294 133150 424350
rect 133218 424294 133274 424350
rect 133342 424294 133398 424350
rect 132970 424170 133026 424226
rect 133094 424170 133150 424226
rect 133218 424170 133274 424226
rect 133342 424170 133398 424226
rect 132970 424046 133026 424102
rect 133094 424046 133150 424102
rect 133218 424046 133274 424102
rect 133342 424046 133398 424102
rect 132970 423922 133026 423978
rect 133094 423922 133150 423978
rect 133218 423922 133274 423978
rect 133342 423922 133398 423978
rect 132970 406294 133026 406350
rect 133094 406294 133150 406350
rect 133218 406294 133274 406350
rect 133342 406294 133398 406350
rect 132970 406170 133026 406226
rect 133094 406170 133150 406226
rect 133218 406170 133274 406226
rect 133342 406170 133398 406226
rect 132970 406046 133026 406102
rect 133094 406046 133150 406102
rect 133218 406046 133274 406102
rect 133342 406046 133398 406102
rect 132970 405922 133026 405978
rect 133094 405922 133150 405978
rect 133218 405922 133274 405978
rect 133342 405922 133398 405978
rect 132970 388294 133026 388350
rect 133094 388294 133150 388350
rect 133218 388294 133274 388350
rect 133342 388294 133398 388350
rect 132970 388170 133026 388226
rect 133094 388170 133150 388226
rect 133218 388170 133274 388226
rect 133342 388170 133398 388226
rect 132970 388046 133026 388102
rect 133094 388046 133150 388102
rect 133218 388046 133274 388102
rect 133342 388046 133398 388102
rect 132970 387922 133026 387978
rect 133094 387922 133150 387978
rect 133218 387922 133274 387978
rect 133342 387922 133398 387978
rect 132970 370294 133026 370350
rect 133094 370294 133150 370350
rect 133218 370294 133274 370350
rect 133342 370294 133398 370350
rect 132970 370170 133026 370226
rect 133094 370170 133150 370226
rect 133218 370170 133274 370226
rect 133342 370170 133398 370226
rect 132970 370046 133026 370102
rect 133094 370046 133150 370102
rect 133218 370046 133274 370102
rect 133342 370046 133398 370102
rect 132970 369922 133026 369978
rect 133094 369922 133150 369978
rect 133218 369922 133274 369978
rect 133342 369922 133398 369978
rect 132970 352294 133026 352350
rect 133094 352294 133150 352350
rect 133218 352294 133274 352350
rect 133342 352294 133398 352350
rect 132970 352170 133026 352226
rect 133094 352170 133150 352226
rect 133218 352170 133274 352226
rect 133342 352170 133398 352226
rect 132970 352046 133026 352102
rect 133094 352046 133150 352102
rect 133218 352046 133274 352102
rect 133342 352046 133398 352102
rect 132970 351922 133026 351978
rect 133094 351922 133150 351978
rect 133218 351922 133274 351978
rect 133342 351922 133398 351978
rect 132970 334294 133026 334350
rect 133094 334294 133150 334350
rect 133218 334294 133274 334350
rect 133342 334294 133398 334350
rect 132970 334170 133026 334226
rect 133094 334170 133150 334226
rect 133218 334170 133274 334226
rect 133342 334170 133398 334226
rect 132970 334046 133026 334102
rect 133094 334046 133150 334102
rect 133218 334046 133274 334102
rect 133342 334046 133398 334102
rect 132970 333922 133026 333978
rect 133094 333922 133150 333978
rect 133218 333922 133274 333978
rect 133342 333922 133398 333978
rect 132970 316294 133026 316350
rect 133094 316294 133150 316350
rect 133218 316294 133274 316350
rect 133342 316294 133398 316350
rect 132970 316170 133026 316226
rect 133094 316170 133150 316226
rect 133218 316170 133274 316226
rect 133342 316170 133398 316226
rect 132970 316046 133026 316102
rect 133094 316046 133150 316102
rect 133218 316046 133274 316102
rect 133342 316046 133398 316102
rect 132970 315922 133026 315978
rect 133094 315922 133150 315978
rect 133218 315922 133274 315978
rect 133342 315922 133398 315978
rect 132970 298294 133026 298350
rect 133094 298294 133150 298350
rect 133218 298294 133274 298350
rect 133342 298294 133398 298350
rect 132970 298170 133026 298226
rect 133094 298170 133150 298226
rect 133218 298170 133274 298226
rect 133342 298170 133398 298226
rect 132970 298046 133026 298102
rect 133094 298046 133150 298102
rect 133218 298046 133274 298102
rect 133342 298046 133398 298102
rect 132970 297922 133026 297978
rect 133094 297922 133150 297978
rect 133218 297922 133274 297978
rect 133342 297922 133398 297978
rect 132970 280294 133026 280350
rect 133094 280294 133150 280350
rect 133218 280294 133274 280350
rect 133342 280294 133398 280350
rect 132970 280170 133026 280226
rect 133094 280170 133150 280226
rect 133218 280170 133274 280226
rect 133342 280170 133398 280226
rect 132970 280046 133026 280102
rect 133094 280046 133150 280102
rect 133218 280046 133274 280102
rect 133342 280046 133398 280102
rect 132970 279922 133026 279978
rect 133094 279922 133150 279978
rect 133218 279922 133274 279978
rect 133342 279922 133398 279978
rect 132970 262294 133026 262350
rect 133094 262294 133150 262350
rect 133218 262294 133274 262350
rect 133342 262294 133398 262350
rect 132970 262170 133026 262226
rect 133094 262170 133150 262226
rect 133218 262170 133274 262226
rect 133342 262170 133398 262226
rect 132970 262046 133026 262102
rect 133094 262046 133150 262102
rect 133218 262046 133274 262102
rect 133342 262046 133398 262102
rect 132970 261922 133026 261978
rect 133094 261922 133150 261978
rect 133218 261922 133274 261978
rect 133342 261922 133398 261978
rect 132970 244294 133026 244350
rect 133094 244294 133150 244350
rect 133218 244294 133274 244350
rect 133342 244294 133398 244350
rect 132970 244170 133026 244226
rect 133094 244170 133150 244226
rect 133218 244170 133274 244226
rect 133342 244170 133398 244226
rect 132970 244046 133026 244102
rect 133094 244046 133150 244102
rect 133218 244046 133274 244102
rect 133342 244046 133398 244102
rect 132970 243922 133026 243978
rect 133094 243922 133150 243978
rect 133218 243922 133274 243978
rect 133342 243922 133398 243978
rect 132970 226294 133026 226350
rect 133094 226294 133150 226350
rect 133218 226294 133274 226350
rect 133342 226294 133398 226350
rect 132970 226170 133026 226226
rect 133094 226170 133150 226226
rect 133218 226170 133274 226226
rect 133342 226170 133398 226226
rect 132970 226046 133026 226102
rect 133094 226046 133150 226102
rect 133218 226046 133274 226102
rect 133342 226046 133398 226102
rect 132970 225922 133026 225978
rect 133094 225922 133150 225978
rect 133218 225922 133274 225978
rect 133342 225922 133398 225978
rect 132970 208294 133026 208350
rect 133094 208294 133150 208350
rect 133218 208294 133274 208350
rect 133342 208294 133398 208350
rect 132970 208170 133026 208226
rect 133094 208170 133150 208226
rect 133218 208170 133274 208226
rect 133342 208170 133398 208226
rect 132970 208046 133026 208102
rect 133094 208046 133150 208102
rect 133218 208046 133274 208102
rect 133342 208046 133398 208102
rect 132970 207922 133026 207978
rect 133094 207922 133150 207978
rect 133218 207922 133274 207978
rect 133342 207922 133398 207978
rect 132970 190294 133026 190350
rect 133094 190294 133150 190350
rect 133218 190294 133274 190350
rect 133342 190294 133398 190350
rect 132970 190170 133026 190226
rect 133094 190170 133150 190226
rect 133218 190170 133274 190226
rect 133342 190170 133398 190226
rect 132970 190046 133026 190102
rect 133094 190046 133150 190102
rect 133218 190046 133274 190102
rect 133342 190046 133398 190102
rect 132970 189922 133026 189978
rect 133094 189922 133150 189978
rect 133218 189922 133274 189978
rect 133342 189922 133398 189978
rect 132970 172294 133026 172350
rect 133094 172294 133150 172350
rect 133218 172294 133274 172350
rect 133342 172294 133398 172350
rect 132970 172170 133026 172226
rect 133094 172170 133150 172226
rect 133218 172170 133274 172226
rect 133342 172170 133398 172226
rect 132970 172046 133026 172102
rect 133094 172046 133150 172102
rect 133218 172046 133274 172102
rect 133342 172046 133398 172102
rect 132970 171922 133026 171978
rect 133094 171922 133150 171978
rect 133218 171922 133274 171978
rect 133342 171922 133398 171978
rect 132970 154294 133026 154350
rect 133094 154294 133150 154350
rect 133218 154294 133274 154350
rect 133342 154294 133398 154350
rect 132970 154170 133026 154226
rect 133094 154170 133150 154226
rect 133218 154170 133274 154226
rect 133342 154170 133398 154226
rect 132970 154046 133026 154102
rect 133094 154046 133150 154102
rect 133218 154046 133274 154102
rect 133342 154046 133398 154102
rect 132970 153922 133026 153978
rect 133094 153922 133150 153978
rect 133218 153922 133274 153978
rect 133342 153922 133398 153978
rect 132970 136294 133026 136350
rect 133094 136294 133150 136350
rect 133218 136294 133274 136350
rect 133342 136294 133398 136350
rect 132970 136170 133026 136226
rect 133094 136170 133150 136226
rect 133218 136170 133274 136226
rect 133342 136170 133398 136226
rect 132970 136046 133026 136102
rect 133094 136046 133150 136102
rect 133218 136046 133274 136102
rect 133342 136046 133398 136102
rect 132970 135922 133026 135978
rect 133094 135922 133150 135978
rect 133218 135922 133274 135978
rect 133342 135922 133398 135978
rect 132970 118294 133026 118350
rect 133094 118294 133150 118350
rect 133218 118294 133274 118350
rect 133342 118294 133398 118350
rect 132970 118170 133026 118226
rect 133094 118170 133150 118226
rect 133218 118170 133274 118226
rect 133342 118170 133398 118226
rect 132970 118046 133026 118102
rect 133094 118046 133150 118102
rect 133218 118046 133274 118102
rect 133342 118046 133398 118102
rect 132970 117922 133026 117978
rect 133094 117922 133150 117978
rect 133218 117922 133274 117978
rect 133342 117922 133398 117978
rect 132970 100294 133026 100350
rect 133094 100294 133150 100350
rect 133218 100294 133274 100350
rect 133342 100294 133398 100350
rect 132970 100170 133026 100226
rect 133094 100170 133150 100226
rect 133218 100170 133274 100226
rect 133342 100170 133398 100226
rect 132970 100046 133026 100102
rect 133094 100046 133150 100102
rect 133218 100046 133274 100102
rect 133342 100046 133398 100102
rect 132970 99922 133026 99978
rect 133094 99922 133150 99978
rect 133218 99922 133274 99978
rect 133342 99922 133398 99978
rect 132970 82294 133026 82350
rect 133094 82294 133150 82350
rect 133218 82294 133274 82350
rect 133342 82294 133398 82350
rect 132970 82170 133026 82226
rect 133094 82170 133150 82226
rect 133218 82170 133274 82226
rect 133342 82170 133398 82226
rect 132970 82046 133026 82102
rect 133094 82046 133150 82102
rect 133218 82046 133274 82102
rect 133342 82046 133398 82102
rect 132970 81922 133026 81978
rect 133094 81922 133150 81978
rect 133218 81922 133274 81978
rect 133342 81922 133398 81978
rect 132970 64294 133026 64350
rect 133094 64294 133150 64350
rect 133218 64294 133274 64350
rect 133342 64294 133398 64350
rect 132970 64170 133026 64226
rect 133094 64170 133150 64226
rect 133218 64170 133274 64226
rect 133342 64170 133398 64226
rect 132970 64046 133026 64102
rect 133094 64046 133150 64102
rect 133218 64046 133274 64102
rect 133342 64046 133398 64102
rect 132970 63922 133026 63978
rect 133094 63922 133150 63978
rect 133218 63922 133274 63978
rect 133342 63922 133398 63978
rect 132970 46294 133026 46350
rect 133094 46294 133150 46350
rect 133218 46294 133274 46350
rect 133342 46294 133398 46350
rect 132970 46170 133026 46226
rect 133094 46170 133150 46226
rect 133218 46170 133274 46226
rect 133342 46170 133398 46226
rect 132970 46046 133026 46102
rect 133094 46046 133150 46102
rect 133218 46046 133274 46102
rect 133342 46046 133398 46102
rect 132970 45922 133026 45978
rect 133094 45922 133150 45978
rect 133218 45922 133274 45978
rect 133342 45922 133398 45978
rect 132970 28294 133026 28350
rect 133094 28294 133150 28350
rect 133218 28294 133274 28350
rect 133342 28294 133398 28350
rect 132970 28170 133026 28226
rect 133094 28170 133150 28226
rect 133218 28170 133274 28226
rect 133342 28170 133398 28226
rect 132970 28046 133026 28102
rect 133094 28046 133150 28102
rect 133218 28046 133274 28102
rect 133342 28046 133398 28102
rect 132970 27922 133026 27978
rect 133094 27922 133150 27978
rect 133218 27922 133274 27978
rect 133342 27922 133398 27978
rect 132970 10294 133026 10350
rect 133094 10294 133150 10350
rect 133218 10294 133274 10350
rect 133342 10294 133398 10350
rect 132970 10170 133026 10226
rect 133094 10170 133150 10226
rect 133218 10170 133274 10226
rect 133342 10170 133398 10226
rect 132970 10046 133026 10102
rect 133094 10046 133150 10102
rect 133218 10046 133274 10102
rect 133342 10046 133398 10102
rect 132970 9922 133026 9978
rect 133094 9922 133150 9978
rect 133218 9922 133274 9978
rect 133342 9922 133398 9978
rect 132970 -1176 133026 -1120
rect 133094 -1176 133150 -1120
rect 133218 -1176 133274 -1120
rect 133342 -1176 133398 -1120
rect 132970 -1300 133026 -1244
rect 133094 -1300 133150 -1244
rect 133218 -1300 133274 -1244
rect 133342 -1300 133398 -1244
rect 132970 -1424 133026 -1368
rect 133094 -1424 133150 -1368
rect 133218 -1424 133274 -1368
rect 133342 -1424 133398 -1368
rect 132970 -1548 133026 -1492
rect 133094 -1548 133150 -1492
rect 133218 -1548 133274 -1492
rect 133342 -1548 133398 -1492
rect 147250 597156 147306 597212
rect 147374 597156 147430 597212
rect 147498 597156 147554 597212
rect 147622 597156 147678 597212
rect 147250 597032 147306 597088
rect 147374 597032 147430 597088
rect 147498 597032 147554 597088
rect 147622 597032 147678 597088
rect 147250 596908 147306 596964
rect 147374 596908 147430 596964
rect 147498 596908 147554 596964
rect 147622 596908 147678 596964
rect 147250 596784 147306 596840
rect 147374 596784 147430 596840
rect 147498 596784 147554 596840
rect 147622 596784 147678 596840
rect 147250 580294 147306 580350
rect 147374 580294 147430 580350
rect 147498 580294 147554 580350
rect 147622 580294 147678 580350
rect 147250 580170 147306 580226
rect 147374 580170 147430 580226
rect 147498 580170 147554 580226
rect 147622 580170 147678 580226
rect 147250 580046 147306 580102
rect 147374 580046 147430 580102
rect 147498 580046 147554 580102
rect 147622 580046 147678 580102
rect 147250 579922 147306 579978
rect 147374 579922 147430 579978
rect 147498 579922 147554 579978
rect 147622 579922 147678 579978
rect 147250 562294 147306 562350
rect 147374 562294 147430 562350
rect 147498 562294 147554 562350
rect 147622 562294 147678 562350
rect 147250 562170 147306 562226
rect 147374 562170 147430 562226
rect 147498 562170 147554 562226
rect 147622 562170 147678 562226
rect 147250 562046 147306 562102
rect 147374 562046 147430 562102
rect 147498 562046 147554 562102
rect 147622 562046 147678 562102
rect 147250 561922 147306 561978
rect 147374 561922 147430 561978
rect 147498 561922 147554 561978
rect 147622 561922 147678 561978
rect 147250 544294 147306 544350
rect 147374 544294 147430 544350
rect 147498 544294 147554 544350
rect 147622 544294 147678 544350
rect 147250 544170 147306 544226
rect 147374 544170 147430 544226
rect 147498 544170 147554 544226
rect 147622 544170 147678 544226
rect 147250 544046 147306 544102
rect 147374 544046 147430 544102
rect 147498 544046 147554 544102
rect 147622 544046 147678 544102
rect 147250 543922 147306 543978
rect 147374 543922 147430 543978
rect 147498 543922 147554 543978
rect 147622 543922 147678 543978
rect 147250 526294 147306 526350
rect 147374 526294 147430 526350
rect 147498 526294 147554 526350
rect 147622 526294 147678 526350
rect 147250 526170 147306 526226
rect 147374 526170 147430 526226
rect 147498 526170 147554 526226
rect 147622 526170 147678 526226
rect 147250 526046 147306 526102
rect 147374 526046 147430 526102
rect 147498 526046 147554 526102
rect 147622 526046 147678 526102
rect 147250 525922 147306 525978
rect 147374 525922 147430 525978
rect 147498 525922 147554 525978
rect 147622 525922 147678 525978
rect 147250 508294 147306 508350
rect 147374 508294 147430 508350
rect 147498 508294 147554 508350
rect 147622 508294 147678 508350
rect 147250 508170 147306 508226
rect 147374 508170 147430 508226
rect 147498 508170 147554 508226
rect 147622 508170 147678 508226
rect 147250 508046 147306 508102
rect 147374 508046 147430 508102
rect 147498 508046 147554 508102
rect 147622 508046 147678 508102
rect 147250 507922 147306 507978
rect 147374 507922 147430 507978
rect 147498 507922 147554 507978
rect 147622 507922 147678 507978
rect 147250 490294 147306 490350
rect 147374 490294 147430 490350
rect 147498 490294 147554 490350
rect 147622 490294 147678 490350
rect 147250 490170 147306 490226
rect 147374 490170 147430 490226
rect 147498 490170 147554 490226
rect 147622 490170 147678 490226
rect 147250 490046 147306 490102
rect 147374 490046 147430 490102
rect 147498 490046 147554 490102
rect 147622 490046 147678 490102
rect 147250 489922 147306 489978
rect 147374 489922 147430 489978
rect 147498 489922 147554 489978
rect 147622 489922 147678 489978
rect 147250 472294 147306 472350
rect 147374 472294 147430 472350
rect 147498 472294 147554 472350
rect 147622 472294 147678 472350
rect 147250 472170 147306 472226
rect 147374 472170 147430 472226
rect 147498 472170 147554 472226
rect 147622 472170 147678 472226
rect 147250 472046 147306 472102
rect 147374 472046 147430 472102
rect 147498 472046 147554 472102
rect 147622 472046 147678 472102
rect 147250 471922 147306 471978
rect 147374 471922 147430 471978
rect 147498 471922 147554 471978
rect 147622 471922 147678 471978
rect 147250 454294 147306 454350
rect 147374 454294 147430 454350
rect 147498 454294 147554 454350
rect 147622 454294 147678 454350
rect 147250 454170 147306 454226
rect 147374 454170 147430 454226
rect 147498 454170 147554 454226
rect 147622 454170 147678 454226
rect 147250 454046 147306 454102
rect 147374 454046 147430 454102
rect 147498 454046 147554 454102
rect 147622 454046 147678 454102
rect 147250 453922 147306 453978
rect 147374 453922 147430 453978
rect 147498 453922 147554 453978
rect 147622 453922 147678 453978
rect 147250 436294 147306 436350
rect 147374 436294 147430 436350
rect 147498 436294 147554 436350
rect 147622 436294 147678 436350
rect 147250 436170 147306 436226
rect 147374 436170 147430 436226
rect 147498 436170 147554 436226
rect 147622 436170 147678 436226
rect 147250 436046 147306 436102
rect 147374 436046 147430 436102
rect 147498 436046 147554 436102
rect 147622 436046 147678 436102
rect 147250 435922 147306 435978
rect 147374 435922 147430 435978
rect 147498 435922 147554 435978
rect 147622 435922 147678 435978
rect 147250 418294 147306 418350
rect 147374 418294 147430 418350
rect 147498 418294 147554 418350
rect 147622 418294 147678 418350
rect 147250 418170 147306 418226
rect 147374 418170 147430 418226
rect 147498 418170 147554 418226
rect 147622 418170 147678 418226
rect 147250 418046 147306 418102
rect 147374 418046 147430 418102
rect 147498 418046 147554 418102
rect 147622 418046 147678 418102
rect 147250 417922 147306 417978
rect 147374 417922 147430 417978
rect 147498 417922 147554 417978
rect 147622 417922 147678 417978
rect 147250 400294 147306 400350
rect 147374 400294 147430 400350
rect 147498 400294 147554 400350
rect 147622 400294 147678 400350
rect 147250 400170 147306 400226
rect 147374 400170 147430 400226
rect 147498 400170 147554 400226
rect 147622 400170 147678 400226
rect 147250 400046 147306 400102
rect 147374 400046 147430 400102
rect 147498 400046 147554 400102
rect 147622 400046 147678 400102
rect 147250 399922 147306 399978
rect 147374 399922 147430 399978
rect 147498 399922 147554 399978
rect 147622 399922 147678 399978
rect 147250 382294 147306 382350
rect 147374 382294 147430 382350
rect 147498 382294 147554 382350
rect 147622 382294 147678 382350
rect 147250 382170 147306 382226
rect 147374 382170 147430 382226
rect 147498 382170 147554 382226
rect 147622 382170 147678 382226
rect 147250 382046 147306 382102
rect 147374 382046 147430 382102
rect 147498 382046 147554 382102
rect 147622 382046 147678 382102
rect 147250 381922 147306 381978
rect 147374 381922 147430 381978
rect 147498 381922 147554 381978
rect 147622 381922 147678 381978
rect 147250 364294 147306 364350
rect 147374 364294 147430 364350
rect 147498 364294 147554 364350
rect 147622 364294 147678 364350
rect 147250 364170 147306 364226
rect 147374 364170 147430 364226
rect 147498 364170 147554 364226
rect 147622 364170 147678 364226
rect 147250 364046 147306 364102
rect 147374 364046 147430 364102
rect 147498 364046 147554 364102
rect 147622 364046 147678 364102
rect 147250 363922 147306 363978
rect 147374 363922 147430 363978
rect 147498 363922 147554 363978
rect 147622 363922 147678 363978
rect 147250 346294 147306 346350
rect 147374 346294 147430 346350
rect 147498 346294 147554 346350
rect 147622 346294 147678 346350
rect 147250 346170 147306 346226
rect 147374 346170 147430 346226
rect 147498 346170 147554 346226
rect 147622 346170 147678 346226
rect 147250 346046 147306 346102
rect 147374 346046 147430 346102
rect 147498 346046 147554 346102
rect 147622 346046 147678 346102
rect 147250 345922 147306 345978
rect 147374 345922 147430 345978
rect 147498 345922 147554 345978
rect 147622 345922 147678 345978
rect 147250 328294 147306 328350
rect 147374 328294 147430 328350
rect 147498 328294 147554 328350
rect 147622 328294 147678 328350
rect 147250 328170 147306 328226
rect 147374 328170 147430 328226
rect 147498 328170 147554 328226
rect 147622 328170 147678 328226
rect 147250 328046 147306 328102
rect 147374 328046 147430 328102
rect 147498 328046 147554 328102
rect 147622 328046 147678 328102
rect 147250 327922 147306 327978
rect 147374 327922 147430 327978
rect 147498 327922 147554 327978
rect 147622 327922 147678 327978
rect 147250 310294 147306 310350
rect 147374 310294 147430 310350
rect 147498 310294 147554 310350
rect 147622 310294 147678 310350
rect 147250 310170 147306 310226
rect 147374 310170 147430 310226
rect 147498 310170 147554 310226
rect 147622 310170 147678 310226
rect 147250 310046 147306 310102
rect 147374 310046 147430 310102
rect 147498 310046 147554 310102
rect 147622 310046 147678 310102
rect 147250 309922 147306 309978
rect 147374 309922 147430 309978
rect 147498 309922 147554 309978
rect 147622 309922 147678 309978
rect 147250 292294 147306 292350
rect 147374 292294 147430 292350
rect 147498 292294 147554 292350
rect 147622 292294 147678 292350
rect 147250 292170 147306 292226
rect 147374 292170 147430 292226
rect 147498 292170 147554 292226
rect 147622 292170 147678 292226
rect 147250 292046 147306 292102
rect 147374 292046 147430 292102
rect 147498 292046 147554 292102
rect 147622 292046 147678 292102
rect 147250 291922 147306 291978
rect 147374 291922 147430 291978
rect 147498 291922 147554 291978
rect 147622 291922 147678 291978
rect 147250 274294 147306 274350
rect 147374 274294 147430 274350
rect 147498 274294 147554 274350
rect 147622 274294 147678 274350
rect 147250 274170 147306 274226
rect 147374 274170 147430 274226
rect 147498 274170 147554 274226
rect 147622 274170 147678 274226
rect 147250 274046 147306 274102
rect 147374 274046 147430 274102
rect 147498 274046 147554 274102
rect 147622 274046 147678 274102
rect 147250 273922 147306 273978
rect 147374 273922 147430 273978
rect 147498 273922 147554 273978
rect 147622 273922 147678 273978
rect 147250 256294 147306 256350
rect 147374 256294 147430 256350
rect 147498 256294 147554 256350
rect 147622 256294 147678 256350
rect 147250 256170 147306 256226
rect 147374 256170 147430 256226
rect 147498 256170 147554 256226
rect 147622 256170 147678 256226
rect 147250 256046 147306 256102
rect 147374 256046 147430 256102
rect 147498 256046 147554 256102
rect 147622 256046 147678 256102
rect 147250 255922 147306 255978
rect 147374 255922 147430 255978
rect 147498 255922 147554 255978
rect 147622 255922 147678 255978
rect 147250 238294 147306 238350
rect 147374 238294 147430 238350
rect 147498 238294 147554 238350
rect 147622 238294 147678 238350
rect 147250 238170 147306 238226
rect 147374 238170 147430 238226
rect 147498 238170 147554 238226
rect 147622 238170 147678 238226
rect 147250 238046 147306 238102
rect 147374 238046 147430 238102
rect 147498 238046 147554 238102
rect 147622 238046 147678 238102
rect 147250 237922 147306 237978
rect 147374 237922 147430 237978
rect 147498 237922 147554 237978
rect 147622 237922 147678 237978
rect 147250 220294 147306 220350
rect 147374 220294 147430 220350
rect 147498 220294 147554 220350
rect 147622 220294 147678 220350
rect 147250 220170 147306 220226
rect 147374 220170 147430 220226
rect 147498 220170 147554 220226
rect 147622 220170 147678 220226
rect 147250 220046 147306 220102
rect 147374 220046 147430 220102
rect 147498 220046 147554 220102
rect 147622 220046 147678 220102
rect 147250 219922 147306 219978
rect 147374 219922 147430 219978
rect 147498 219922 147554 219978
rect 147622 219922 147678 219978
rect 147250 202294 147306 202350
rect 147374 202294 147430 202350
rect 147498 202294 147554 202350
rect 147622 202294 147678 202350
rect 147250 202170 147306 202226
rect 147374 202170 147430 202226
rect 147498 202170 147554 202226
rect 147622 202170 147678 202226
rect 147250 202046 147306 202102
rect 147374 202046 147430 202102
rect 147498 202046 147554 202102
rect 147622 202046 147678 202102
rect 147250 201922 147306 201978
rect 147374 201922 147430 201978
rect 147498 201922 147554 201978
rect 147622 201922 147678 201978
rect 147250 184294 147306 184350
rect 147374 184294 147430 184350
rect 147498 184294 147554 184350
rect 147622 184294 147678 184350
rect 147250 184170 147306 184226
rect 147374 184170 147430 184226
rect 147498 184170 147554 184226
rect 147622 184170 147678 184226
rect 147250 184046 147306 184102
rect 147374 184046 147430 184102
rect 147498 184046 147554 184102
rect 147622 184046 147678 184102
rect 147250 183922 147306 183978
rect 147374 183922 147430 183978
rect 147498 183922 147554 183978
rect 147622 183922 147678 183978
rect 147250 166294 147306 166350
rect 147374 166294 147430 166350
rect 147498 166294 147554 166350
rect 147622 166294 147678 166350
rect 147250 166170 147306 166226
rect 147374 166170 147430 166226
rect 147498 166170 147554 166226
rect 147622 166170 147678 166226
rect 147250 166046 147306 166102
rect 147374 166046 147430 166102
rect 147498 166046 147554 166102
rect 147622 166046 147678 166102
rect 147250 165922 147306 165978
rect 147374 165922 147430 165978
rect 147498 165922 147554 165978
rect 147622 165922 147678 165978
rect 147250 148294 147306 148350
rect 147374 148294 147430 148350
rect 147498 148294 147554 148350
rect 147622 148294 147678 148350
rect 147250 148170 147306 148226
rect 147374 148170 147430 148226
rect 147498 148170 147554 148226
rect 147622 148170 147678 148226
rect 147250 148046 147306 148102
rect 147374 148046 147430 148102
rect 147498 148046 147554 148102
rect 147622 148046 147678 148102
rect 147250 147922 147306 147978
rect 147374 147922 147430 147978
rect 147498 147922 147554 147978
rect 147622 147922 147678 147978
rect 147250 130294 147306 130350
rect 147374 130294 147430 130350
rect 147498 130294 147554 130350
rect 147622 130294 147678 130350
rect 147250 130170 147306 130226
rect 147374 130170 147430 130226
rect 147498 130170 147554 130226
rect 147622 130170 147678 130226
rect 147250 130046 147306 130102
rect 147374 130046 147430 130102
rect 147498 130046 147554 130102
rect 147622 130046 147678 130102
rect 147250 129922 147306 129978
rect 147374 129922 147430 129978
rect 147498 129922 147554 129978
rect 147622 129922 147678 129978
rect 147250 112294 147306 112350
rect 147374 112294 147430 112350
rect 147498 112294 147554 112350
rect 147622 112294 147678 112350
rect 147250 112170 147306 112226
rect 147374 112170 147430 112226
rect 147498 112170 147554 112226
rect 147622 112170 147678 112226
rect 147250 112046 147306 112102
rect 147374 112046 147430 112102
rect 147498 112046 147554 112102
rect 147622 112046 147678 112102
rect 147250 111922 147306 111978
rect 147374 111922 147430 111978
rect 147498 111922 147554 111978
rect 147622 111922 147678 111978
rect 147250 94294 147306 94350
rect 147374 94294 147430 94350
rect 147498 94294 147554 94350
rect 147622 94294 147678 94350
rect 147250 94170 147306 94226
rect 147374 94170 147430 94226
rect 147498 94170 147554 94226
rect 147622 94170 147678 94226
rect 147250 94046 147306 94102
rect 147374 94046 147430 94102
rect 147498 94046 147554 94102
rect 147622 94046 147678 94102
rect 147250 93922 147306 93978
rect 147374 93922 147430 93978
rect 147498 93922 147554 93978
rect 147622 93922 147678 93978
rect 147250 76294 147306 76350
rect 147374 76294 147430 76350
rect 147498 76294 147554 76350
rect 147622 76294 147678 76350
rect 147250 76170 147306 76226
rect 147374 76170 147430 76226
rect 147498 76170 147554 76226
rect 147622 76170 147678 76226
rect 147250 76046 147306 76102
rect 147374 76046 147430 76102
rect 147498 76046 147554 76102
rect 147622 76046 147678 76102
rect 147250 75922 147306 75978
rect 147374 75922 147430 75978
rect 147498 75922 147554 75978
rect 147622 75922 147678 75978
rect 147250 58294 147306 58350
rect 147374 58294 147430 58350
rect 147498 58294 147554 58350
rect 147622 58294 147678 58350
rect 147250 58170 147306 58226
rect 147374 58170 147430 58226
rect 147498 58170 147554 58226
rect 147622 58170 147678 58226
rect 147250 58046 147306 58102
rect 147374 58046 147430 58102
rect 147498 58046 147554 58102
rect 147622 58046 147678 58102
rect 147250 57922 147306 57978
rect 147374 57922 147430 57978
rect 147498 57922 147554 57978
rect 147622 57922 147678 57978
rect 147250 40294 147306 40350
rect 147374 40294 147430 40350
rect 147498 40294 147554 40350
rect 147622 40294 147678 40350
rect 147250 40170 147306 40226
rect 147374 40170 147430 40226
rect 147498 40170 147554 40226
rect 147622 40170 147678 40226
rect 147250 40046 147306 40102
rect 147374 40046 147430 40102
rect 147498 40046 147554 40102
rect 147622 40046 147678 40102
rect 147250 39922 147306 39978
rect 147374 39922 147430 39978
rect 147498 39922 147554 39978
rect 147622 39922 147678 39978
rect 147250 22294 147306 22350
rect 147374 22294 147430 22350
rect 147498 22294 147554 22350
rect 147622 22294 147678 22350
rect 147250 22170 147306 22226
rect 147374 22170 147430 22226
rect 147498 22170 147554 22226
rect 147622 22170 147678 22226
rect 147250 22046 147306 22102
rect 147374 22046 147430 22102
rect 147498 22046 147554 22102
rect 147622 22046 147678 22102
rect 147250 21922 147306 21978
rect 147374 21922 147430 21978
rect 147498 21922 147554 21978
rect 147622 21922 147678 21978
rect 147250 4294 147306 4350
rect 147374 4294 147430 4350
rect 147498 4294 147554 4350
rect 147622 4294 147678 4350
rect 147250 4170 147306 4226
rect 147374 4170 147430 4226
rect 147498 4170 147554 4226
rect 147622 4170 147678 4226
rect 147250 4046 147306 4102
rect 147374 4046 147430 4102
rect 147498 4046 147554 4102
rect 147622 4046 147678 4102
rect 147250 3922 147306 3978
rect 147374 3922 147430 3978
rect 147498 3922 147554 3978
rect 147622 3922 147678 3978
rect 147250 -216 147306 -160
rect 147374 -216 147430 -160
rect 147498 -216 147554 -160
rect 147622 -216 147678 -160
rect 147250 -340 147306 -284
rect 147374 -340 147430 -284
rect 147498 -340 147554 -284
rect 147622 -340 147678 -284
rect 147250 -464 147306 -408
rect 147374 -464 147430 -408
rect 147498 -464 147554 -408
rect 147622 -464 147678 -408
rect 147250 -588 147306 -532
rect 147374 -588 147430 -532
rect 147498 -588 147554 -532
rect 147622 -588 147678 -532
rect 150970 598116 151026 598172
rect 151094 598116 151150 598172
rect 151218 598116 151274 598172
rect 151342 598116 151398 598172
rect 150970 597992 151026 598048
rect 151094 597992 151150 598048
rect 151218 597992 151274 598048
rect 151342 597992 151398 598048
rect 150970 597868 151026 597924
rect 151094 597868 151150 597924
rect 151218 597868 151274 597924
rect 151342 597868 151398 597924
rect 150970 597744 151026 597800
rect 151094 597744 151150 597800
rect 151218 597744 151274 597800
rect 151342 597744 151398 597800
rect 150970 586294 151026 586350
rect 151094 586294 151150 586350
rect 151218 586294 151274 586350
rect 151342 586294 151398 586350
rect 150970 586170 151026 586226
rect 151094 586170 151150 586226
rect 151218 586170 151274 586226
rect 151342 586170 151398 586226
rect 150970 586046 151026 586102
rect 151094 586046 151150 586102
rect 151218 586046 151274 586102
rect 151342 586046 151398 586102
rect 150970 585922 151026 585978
rect 151094 585922 151150 585978
rect 151218 585922 151274 585978
rect 151342 585922 151398 585978
rect 150970 568294 151026 568350
rect 151094 568294 151150 568350
rect 151218 568294 151274 568350
rect 151342 568294 151398 568350
rect 150970 568170 151026 568226
rect 151094 568170 151150 568226
rect 151218 568170 151274 568226
rect 151342 568170 151398 568226
rect 150970 568046 151026 568102
rect 151094 568046 151150 568102
rect 151218 568046 151274 568102
rect 151342 568046 151398 568102
rect 150970 567922 151026 567978
rect 151094 567922 151150 567978
rect 151218 567922 151274 567978
rect 151342 567922 151398 567978
rect 150970 550294 151026 550350
rect 151094 550294 151150 550350
rect 151218 550294 151274 550350
rect 151342 550294 151398 550350
rect 150970 550170 151026 550226
rect 151094 550170 151150 550226
rect 151218 550170 151274 550226
rect 151342 550170 151398 550226
rect 150970 550046 151026 550102
rect 151094 550046 151150 550102
rect 151218 550046 151274 550102
rect 151342 550046 151398 550102
rect 150970 549922 151026 549978
rect 151094 549922 151150 549978
rect 151218 549922 151274 549978
rect 151342 549922 151398 549978
rect 150970 532294 151026 532350
rect 151094 532294 151150 532350
rect 151218 532294 151274 532350
rect 151342 532294 151398 532350
rect 150970 532170 151026 532226
rect 151094 532170 151150 532226
rect 151218 532170 151274 532226
rect 151342 532170 151398 532226
rect 150970 532046 151026 532102
rect 151094 532046 151150 532102
rect 151218 532046 151274 532102
rect 151342 532046 151398 532102
rect 150970 531922 151026 531978
rect 151094 531922 151150 531978
rect 151218 531922 151274 531978
rect 151342 531922 151398 531978
rect 150970 514294 151026 514350
rect 151094 514294 151150 514350
rect 151218 514294 151274 514350
rect 151342 514294 151398 514350
rect 150970 514170 151026 514226
rect 151094 514170 151150 514226
rect 151218 514170 151274 514226
rect 151342 514170 151398 514226
rect 150970 514046 151026 514102
rect 151094 514046 151150 514102
rect 151218 514046 151274 514102
rect 151342 514046 151398 514102
rect 150970 513922 151026 513978
rect 151094 513922 151150 513978
rect 151218 513922 151274 513978
rect 151342 513922 151398 513978
rect 150970 496294 151026 496350
rect 151094 496294 151150 496350
rect 151218 496294 151274 496350
rect 151342 496294 151398 496350
rect 150970 496170 151026 496226
rect 151094 496170 151150 496226
rect 151218 496170 151274 496226
rect 151342 496170 151398 496226
rect 150970 496046 151026 496102
rect 151094 496046 151150 496102
rect 151218 496046 151274 496102
rect 151342 496046 151398 496102
rect 150970 495922 151026 495978
rect 151094 495922 151150 495978
rect 151218 495922 151274 495978
rect 151342 495922 151398 495978
rect 150970 478294 151026 478350
rect 151094 478294 151150 478350
rect 151218 478294 151274 478350
rect 151342 478294 151398 478350
rect 150970 478170 151026 478226
rect 151094 478170 151150 478226
rect 151218 478170 151274 478226
rect 151342 478170 151398 478226
rect 150970 478046 151026 478102
rect 151094 478046 151150 478102
rect 151218 478046 151274 478102
rect 151342 478046 151398 478102
rect 150970 477922 151026 477978
rect 151094 477922 151150 477978
rect 151218 477922 151274 477978
rect 151342 477922 151398 477978
rect 150970 460294 151026 460350
rect 151094 460294 151150 460350
rect 151218 460294 151274 460350
rect 151342 460294 151398 460350
rect 150970 460170 151026 460226
rect 151094 460170 151150 460226
rect 151218 460170 151274 460226
rect 151342 460170 151398 460226
rect 150970 460046 151026 460102
rect 151094 460046 151150 460102
rect 151218 460046 151274 460102
rect 151342 460046 151398 460102
rect 150970 459922 151026 459978
rect 151094 459922 151150 459978
rect 151218 459922 151274 459978
rect 151342 459922 151398 459978
rect 150970 442294 151026 442350
rect 151094 442294 151150 442350
rect 151218 442294 151274 442350
rect 151342 442294 151398 442350
rect 150970 442170 151026 442226
rect 151094 442170 151150 442226
rect 151218 442170 151274 442226
rect 151342 442170 151398 442226
rect 150970 442046 151026 442102
rect 151094 442046 151150 442102
rect 151218 442046 151274 442102
rect 151342 442046 151398 442102
rect 150970 441922 151026 441978
rect 151094 441922 151150 441978
rect 151218 441922 151274 441978
rect 151342 441922 151398 441978
rect 150970 424294 151026 424350
rect 151094 424294 151150 424350
rect 151218 424294 151274 424350
rect 151342 424294 151398 424350
rect 150970 424170 151026 424226
rect 151094 424170 151150 424226
rect 151218 424170 151274 424226
rect 151342 424170 151398 424226
rect 150970 424046 151026 424102
rect 151094 424046 151150 424102
rect 151218 424046 151274 424102
rect 151342 424046 151398 424102
rect 150970 423922 151026 423978
rect 151094 423922 151150 423978
rect 151218 423922 151274 423978
rect 151342 423922 151398 423978
rect 150970 406294 151026 406350
rect 151094 406294 151150 406350
rect 151218 406294 151274 406350
rect 151342 406294 151398 406350
rect 150970 406170 151026 406226
rect 151094 406170 151150 406226
rect 151218 406170 151274 406226
rect 151342 406170 151398 406226
rect 150970 406046 151026 406102
rect 151094 406046 151150 406102
rect 151218 406046 151274 406102
rect 151342 406046 151398 406102
rect 150970 405922 151026 405978
rect 151094 405922 151150 405978
rect 151218 405922 151274 405978
rect 151342 405922 151398 405978
rect 150970 388294 151026 388350
rect 151094 388294 151150 388350
rect 151218 388294 151274 388350
rect 151342 388294 151398 388350
rect 150970 388170 151026 388226
rect 151094 388170 151150 388226
rect 151218 388170 151274 388226
rect 151342 388170 151398 388226
rect 150970 388046 151026 388102
rect 151094 388046 151150 388102
rect 151218 388046 151274 388102
rect 151342 388046 151398 388102
rect 150970 387922 151026 387978
rect 151094 387922 151150 387978
rect 151218 387922 151274 387978
rect 151342 387922 151398 387978
rect 150970 370294 151026 370350
rect 151094 370294 151150 370350
rect 151218 370294 151274 370350
rect 151342 370294 151398 370350
rect 150970 370170 151026 370226
rect 151094 370170 151150 370226
rect 151218 370170 151274 370226
rect 151342 370170 151398 370226
rect 150970 370046 151026 370102
rect 151094 370046 151150 370102
rect 151218 370046 151274 370102
rect 151342 370046 151398 370102
rect 150970 369922 151026 369978
rect 151094 369922 151150 369978
rect 151218 369922 151274 369978
rect 151342 369922 151398 369978
rect 150970 352294 151026 352350
rect 151094 352294 151150 352350
rect 151218 352294 151274 352350
rect 151342 352294 151398 352350
rect 150970 352170 151026 352226
rect 151094 352170 151150 352226
rect 151218 352170 151274 352226
rect 151342 352170 151398 352226
rect 150970 352046 151026 352102
rect 151094 352046 151150 352102
rect 151218 352046 151274 352102
rect 151342 352046 151398 352102
rect 150970 351922 151026 351978
rect 151094 351922 151150 351978
rect 151218 351922 151274 351978
rect 151342 351922 151398 351978
rect 150970 334294 151026 334350
rect 151094 334294 151150 334350
rect 151218 334294 151274 334350
rect 151342 334294 151398 334350
rect 150970 334170 151026 334226
rect 151094 334170 151150 334226
rect 151218 334170 151274 334226
rect 151342 334170 151398 334226
rect 150970 334046 151026 334102
rect 151094 334046 151150 334102
rect 151218 334046 151274 334102
rect 151342 334046 151398 334102
rect 150970 333922 151026 333978
rect 151094 333922 151150 333978
rect 151218 333922 151274 333978
rect 151342 333922 151398 333978
rect 150970 316294 151026 316350
rect 151094 316294 151150 316350
rect 151218 316294 151274 316350
rect 151342 316294 151398 316350
rect 150970 316170 151026 316226
rect 151094 316170 151150 316226
rect 151218 316170 151274 316226
rect 151342 316170 151398 316226
rect 150970 316046 151026 316102
rect 151094 316046 151150 316102
rect 151218 316046 151274 316102
rect 151342 316046 151398 316102
rect 150970 315922 151026 315978
rect 151094 315922 151150 315978
rect 151218 315922 151274 315978
rect 151342 315922 151398 315978
rect 150970 298294 151026 298350
rect 151094 298294 151150 298350
rect 151218 298294 151274 298350
rect 151342 298294 151398 298350
rect 150970 298170 151026 298226
rect 151094 298170 151150 298226
rect 151218 298170 151274 298226
rect 151342 298170 151398 298226
rect 150970 298046 151026 298102
rect 151094 298046 151150 298102
rect 151218 298046 151274 298102
rect 151342 298046 151398 298102
rect 150970 297922 151026 297978
rect 151094 297922 151150 297978
rect 151218 297922 151274 297978
rect 151342 297922 151398 297978
rect 150970 280294 151026 280350
rect 151094 280294 151150 280350
rect 151218 280294 151274 280350
rect 151342 280294 151398 280350
rect 150970 280170 151026 280226
rect 151094 280170 151150 280226
rect 151218 280170 151274 280226
rect 151342 280170 151398 280226
rect 150970 280046 151026 280102
rect 151094 280046 151150 280102
rect 151218 280046 151274 280102
rect 151342 280046 151398 280102
rect 150970 279922 151026 279978
rect 151094 279922 151150 279978
rect 151218 279922 151274 279978
rect 151342 279922 151398 279978
rect 150970 262294 151026 262350
rect 151094 262294 151150 262350
rect 151218 262294 151274 262350
rect 151342 262294 151398 262350
rect 150970 262170 151026 262226
rect 151094 262170 151150 262226
rect 151218 262170 151274 262226
rect 151342 262170 151398 262226
rect 150970 262046 151026 262102
rect 151094 262046 151150 262102
rect 151218 262046 151274 262102
rect 151342 262046 151398 262102
rect 150970 261922 151026 261978
rect 151094 261922 151150 261978
rect 151218 261922 151274 261978
rect 151342 261922 151398 261978
rect 150970 244294 151026 244350
rect 151094 244294 151150 244350
rect 151218 244294 151274 244350
rect 151342 244294 151398 244350
rect 150970 244170 151026 244226
rect 151094 244170 151150 244226
rect 151218 244170 151274 244226
rect 151342 244170 151398 244226
rect 150970 244046 151026 244102
rect 151094 244046 151150 244102
rect 151218 244046 151274 244102
rect 151342 244046 151398 244102
rect 150970 243922 151026 243978
rect 151094 243922 151150 243978
rect 151218 243922 151274 243978
rect 151342 243922 151398 243978
rect 150970 226294 151026 226350
rect 151094 226294 151150 226350
rect 151218 226294 151274 226350
rect 151342 226294 151398 226350
rect 150970 226170 151026 226226
rect 151094 226170 151150 226226
rect 151218 226170 151274 226226
rect 151342 226170 151398 226226
rect 150970 226046 151026 226102
rect 151094 226046 151150 226102
rect 151218 226046 151274 226102
rect 151342 226046 151398 226102
rect 150970 225922 151026 225978
rect 151094 225922 151150 225978
rect 151218 225922 151274 225978
rect 151342 225922 151398 225978
rect 150970 208294 151026 208350
rect 151094 208294 151150 208350
rect 151218 208294 151274 208350
rect 151342 208294 151398 208350
rect 150970 208170 151026 208226
rect 151094 208170 151150 208226
rect 151218 208170 151274 208226
rect 151342 208170 151398 208226
rect 150970 208046 151026 208102
rect 151094 208046 151150 208102
rect 151218 208046 151274 208102
rect 151342 208046 151398 208102
rect 150970 207922 151026 207978
rect 151094 207922 151150 207978
rect 151218 207922 151274 207978
rect 151342 207922 151398 207978
rect 150970 190294 151026 190350
rect 151094 190294 151150 190350
rect 151218 190294 151274 190350
rect 151342 190294 151398 190350
rect 150970 190170 151026 190226
rect 151094 190170 151150 190226
rect 151218 190170 151274 190226
rect 151342 190170 151398 190226
rect 150970 190046 151026 190102
rect 151094 190046 151150 190102
rect 151218 190046 151274 190102
rect 151342 190046 151398 190102
rect 150970 189922 151026 189978
rect 151094 189922 151150 189978
rect 151218 189922 151274 189978
rect 151342 189922 151398 189978
rect 150970 172294 151026 172350
rect 151094 172294 151150 172350
rect 151218 172294 151274 172350
rect 151342 172294 151398 172350
rect 150970 172170 151026 172226
rect 151094 172170 151150 172226
rect 151218 172170 151274 172226
rect 151342 172170 151398 172226
rect 150970 172046 151026 172102
rect 151094 172046 151150 172102
rect 151218 172046 151274 172102
rect 151342 172046 151398 172102
rect 150970 171922 151026 171978
rect 151094 171922 151150 171978
rect 151218 171922 151274 171978
rect 151342 171922 151398 171978
rect 150970 154294 151026 154350
rect 151094 154294 151150 154350
rect 151218 154294 151274 154350
rect 151342 154294 151398 154350
rect 150970 154170 151026 154226
rect 151094 154170 151150 154226
rect 151218 154170 151274 154226
rect 151342 154170 151398 154226
rect 150970 154046 151026 154102
rect 151094 154046 151150 154102
rect 151218 154046 151274 154102
rect 151342 154046 151398 154102
rect 150970 153922 151026 153978
rect 151094 153922 151150 153978
rect 151218 153922 151274 153978
rect 151342 153922 151398 153978
rect 150970 136294 151026 136350
rect 151094 136294 151150 136350
rect 151218 136294 151274 136350
rect 151342 136294 151398 136350
rect 150970 136170 151026 136226
rect 151094 136170 151150 136226
rect 151218 136170 151274 136226
rect 151342 136170 151398 136226
rect 150970 136046 151026 136102
rect 151094 136046 151150 136102
rect 151218 136046 151274 136102
rect 151342 136046 151398 136102
rect 150970 135922 151026 135978
rect 151094 135922 151150 135978
rect 151218 135922 151274 135978
rect 151342 135922 151398 135978
rect 150970 118294 151026 118350
rect 151094 118294 151150 118350
rect 151218 118294 151274 118350
rect 151342 118294 151398 118350
rect 150970 118170 151026 118226
rect 151094 118170 151150 118226
rect 151218 118170 151274 118226
rect 151342 118170 151398 118226
rect 150970 118046 151026 118102
rect 151094 118046 151150 118102
rect 151218 118046 151274 118102
rect 151342 118046 151398 118102
rect 150970 117922 151026 117978
rect 151094 117922 151150 117978
rect 151218 117922 151274 117978
rect 151342 117922 151398 117978
rect 150970 100294 151026 100350
rect 151094 100294 151150 100350
rect 151218 100294 151274 100350
rect 151342 100294 151398 100350
rect 150970 100170 151026 100226
rect 151094 100170 151150 100226
rect 151218 100170 151274 100226
rect 151342 100170 151398 100226
rect 150970 100046 151026 100102
rect 151094 100046 151150 100102
rect 151218 100046 151274 100102
rect 151342 100046 151398 100102
rect 150970 99922 151026 99978
rect 151094 99922 151150 99978
rect 151218 99922 151274 99978
rect 151342 99922 151398 99978
rect 150970 82294 151026 82350
rect 151094 82294 151150 82350
rect 151218 82294 151274 82350
rect 151342 82294 151398 82350
rect 150970 82170 151026 82226
rect 151094 82170 151150 82226
rect 151218 82170 151274 82226
rect 151342 82170 151398 82226
rect 150970 82046 151026 82102
rect 151094 82046 151150 82102
rect 151218 82046 151274 82102
rect 151342 82046 151398 82102
rect 150970 81922 151026 81978
rect 151094 81922 151150 81978
rect 151218 81922 151274 81978
rect 151342 81922 151398 81978
rect 150970 64294 151026 64350
rect 151094 64294 151150 64350
rect 151218 64294 151274 64350
rect 151342 64294 151398 64350
rect 150970 64170 151026 64226
rect 151094 64170 151150 64226
rect 151218 64170 151274 64226
rect 151342 64170 151398 64226
rect 150970 64046 151026 64102
rect 151094 64046 151150 64102
rect 151218 64046 151274 64102
rect 151342 64046 151398 64102
rect 150970 63922 151026 63978
rect 151094 63922 151150 63978
rect 151218 63922 151274 63978
rect 151342 63922 151398 63978
rect 150970 46294 151026 46350
rect 151094 46294 151150 46350
rect 151218 46294 151274 46350
rect 151342 46294 151398 46350
rect 150970 46170 151026 46226
rect 151094 46170 151150 46226
rect 151218 46170 151274 46226
rect 151342 46170 151398 46226
rect 150970 46046 151026 46102
rect 151094 46046 151150 46102
rect 151218 46046 151274 46102
rect 151342 46046 151398 46102
rect 150970 45922 151026 45978
rect 151094 45922 151150 45978
rect 151218 45922 151274 45978
rect 151342 45922 151398 45978
rect 150970 28294 151026 28350
rect 151094 28294 151150 28350
rect 151218 28294 151274 28350
rect 151342 28294 151398 28350
rect 150970 28170 151026 28226
rect 151094 28170 151150 28226
rect 151218 28170 151274 28226
rect 151342 28170 151398 28226
rect 150970 28046 151026 28102
rect 151094 28046 151150 28102
rect 151218 28046 151274 28102
rect 151342 28046 151398 28102
rect 150970 27922 151026 27978
rect 151094 27922 151150 27978
rect 151218 27922 151274 27978
rect 151342 27922 151398 27978
rect 150970 10294 151026 10350
rect 151094 10294 151150 10350
rect 151218 10294 151274 10350
rect 151342 10294 151398 10350
rect 150970 10170 151026 10226
rect 151094 10170 151150 10226
rect 151218 10170 151274 10226
rect 151342 10170 151398 10226
rect 150970 10046 151026 10102
rect 151094 10046 151150 10102
rect 151218 10046 151274 10102
rect 151342 10046 151398 10102
rect 150970 9922 151026 9978
rect 151094 9922 151150 9978
rect 151218 9922 151274 9978
rect 151342 9922 151398 9978
rect 150970 -1176 151026 -1120
rect 151094 -1176 151150 -1120
rect 151218 -1176 151274 -1120
rect 151342 -1176 151398 -1120
rect 150970 -1300 151026 -1244
rect 151094 -1300 151150 -1244
rect 151218 -1300 151274 -1244
rect 151342 -1300 151398 -1244
rect 150970 -1424 151026 -1368
rect 151094 -1424 151150 -1368
rect 151218 -1424 151274 -1368
rect 151342 -1424 151398 -1368
rect 150970 -1548 151026 -1492
rect 151094 -1548 151150 -1492
rect 151218 -1548 151274 -1492
rect 151342 -1548 151398 -1492
rect 165250 597156 165306 597212
rect 165374 597156 165430 597212
rect 165498 597156 165554 597212
rect 165622 597156 165678 597212
rect 165250 597032 165306 597088
rect 165374 597032 165430 597088
rect 165498 597032 165554 597088
rect 165622 597032 165678 597088
rect 165250 596908 165306 596964
rect 165374 596908 165430 596964
rect 165498 596908 165554 596964
rect 165622 596908 165678 596964
rect 165250 596784 165306 596840
rect 165374 596784 165430 596840
rect 165498 596784 165554 596840
rect 165622 596784 165678 596840
rect 165250 580294 165306 580350
rect 165374 580294 165430 580350
rect 165498 580294 165554 580350
rect 165622 580294 165678 580350
rect 165250 580170 165306 580226
rect 165374 580170 165430 580226
rect 165498 580170 165554 580226
rect 165622 580170 165678 580226
rect 165250 580046 165306 580102
rect 165374 580046 165430 580102
rect 165498 580046 165554 580102
rect 165622 580046 165678 580102
rect 165250 579922 165306 579978
rect 165374 579922 165430 579978
rect 165498 579922 165554 579978
rect 165622 579922 165678 579978
rect 165250 562294 165306 562350
rect 165374 562294 165430 562350
rect 165498 562294 165554 562350
rect 165622 562294 165678 562350
rect 165250 562170 165306 562226
rect 165374 562170 165430 562226
rect 165498 562170 165554 562226
rect 165622 562170 165678 562226
rect 165250 562046 165306 562102
rect 165374 562046 165430 562102
rect 165498 562046 165554 562102
rect 165622 562046 165678 562102
rect 165250 561922 165306 561978
rect 165374 561922 165430 561978
rect 165498 561922 165554 561978
rect 165622 561922 165678 561978
rect 165250 544294 165306 544350
rect 165374 544294 165430 544350
rect 165498 544294 165554 544350
rect 165622 544294 165678 544350
rect 165250 544170 165306 544226
rect 165374 544170 165430 544226
rect 165498 544170 165554 544226
rect 165622 544170 165678 544226
rect 165250 544046 165306 544102
rect 165374 544046 165430 544102
rect 165498 544046 165554 544102
rect 165622 544046 165678 544102
rect 165250 543922 165306 543978
rect 165374 543922 165430 543978
rect 165498 543922 165554 543978
rect 165622 543922 165678 543978
rect 165250 526294 165306 526350
rect 165374 526294 165430 526350
rect 165498 526294 165554 526350
rect 165622 526294 165678 526350
rect 165250 526170 165306 526226
rect 165374 526170 165430 526226
rect 165498 526170 165554 526226
rect 165622 526170 165678 526226
rect 165250 526046 165306 526102
rect 165374 526046 165430 526102
rect 165498 526046 165554 526102
rect 165622 526046 165678 526102
rect 165250 525922 165306 525978
rect 165374 525922 165430 525978
rect 165498 525922 165554 525978
rect 165622 525922 165678 525978
rect 165250 508294 165306 508350
rect 165374 508294 165430 508350
rect 165498 508294 165554 508350
rect 165622 508294 165678 508350
rect 165250 508170 165306 508226
rect 165374 508170 165430 508226
rect 165498 508170 165554 508226
rect 165622 508170 165678 508226
rect 165250 508046 165306 508102
rect 165374 508046 165430 508102
rect 165498 508046 165554 508102
rect 165622 508046 165678 508102
rect 165250 507922 165306 507978
rect 165374 507922 165430 507978
rect 165498 507922 165554 507978
rect 165622 507922 165678 507978
rect 165250 490294 165306 490350
rect 165374 490294 165430 490350
rect 165498 490294 165554 490350
rect 165622 490294 165678 490350
rect 165250 490170 165306 490226
rect 165374 490170 165430 490226
rect 165498 490170 165554 490226
rect 165622 490170 165678 490226
rect 165250 490046 165306 490102
rect 165374 490046 165430 490102
rect 165498 490046 165554 490102
rect 165622 490046 165678 490102
rect 165250 489922 165306 489978
rect 165374 489922 165430 489978
rect 165498 489922 165554 489978
rect 165622 489922 165678 489978
rect 165250 472294 165306 472350
rect 165374 472294 165430 472350
rect 165498 472294 165554 472350
rect 165622 472294 165678 472350
rect 165250 472170 165306 472226
rect 165374 472170 165430 472226
rect 165498 472170 165554 472226
rect 165622 472170 165678 472226
rect 165250 472046 165306 472102
rect 165374 472046 165430 472102
rect 165498 472046 165554 472102
rect 165622 472046 165678 472102
rect 165250 471922 165306 471978
rect 165374 471922 165430 471978
rect 165498 471922 165554 471978
rect 165622 471922 165678 471978
rect 165250 454294 165306 454350
rect 165374 454294 165430 454350
rect 165498 454294 165554 454350
rect 165622 454294 165678 454350
rect 165250 454170 165306 454226
rect 165374 454170 165430 454226
rect 165498 454170 165554 454226
rect 165622 454170 165678 454226
rect 165250 454046 165306 454102
rect 165374 454046 165430 454102
rect 165498 454046 165554 454102
rect 165622 454046 165678 454102
rect 165250 453922 165306 453978
rect 165374 453922 165430 453978
rect 165498 453922 165554 453978
rect 165622 453922 165678 453978
rect 165250 436294 165306 436350
rect 165374 436294 165430 436350
rect 165498 436294 165554 436350
rect 165622 436294 165678 436350
rect 165250 436170 165306 436226
rect 165374 436170 165430 436226
rect 165498 436170 165554 436226
rect 165622 436170 165678 436226
rect 165250 436046 165306 436102
rect 165374 436046 165430 436102
rect 165498 436046 165554 436102
rect 165622 436046 165678 436102
rect 165250 435922 165306 435978
rect 165374 435922 165430 435978
rect 165498 435922 165554 435978
rect 165622 435922 165678 435978
rect 165250 418294 165306 418350
rect 165374 418294 165430 418350
rect 165498 418294 165554 418350
rect 165622 418294 165678 418350
rect 165250 418170 165306 418226
rect 165374 418170 165430 418226
rect 165498 418170 165554 418226
rect 165622 418170 165678 418226
rect 165250 418046 165306 418102
rect 165374 418046 165430 418102
rect 165498 418046 165554 418102
rect 165622 418046 165678 418102
rect 165250 417922 165306 417978
rect 165374 417922 165430 417978
rect 165498 417922 165554 417978
rect 165622 417922 165678 417978
rect 165250 400294 165306 400350
rect 165374 400294 165430 400350
rect 165498 400294 165554 400350
rect 165622 400294 165678 400350
rect 165250 400170 165306 400226
rect 165374 400170 165430 400226
rect 165498 400170 165554 400226
rect 165622 400170 165678 400226
rect 165250 400046 165306 400102
rect 165374 400046 165430 400102
rect 165498 400046 165554 400102
rect 165622 400046 165678 400102
rect 165250 399922 165306 399978
rect 165374 399922 165430 399978
rect 165498 399922 165554 399978
rect 165622 399922 165678 399978
rect 165250 382294 165306 382350
rect 165374 382294 165430 382350
rect 165498 382294 165554 382350
rect 165622 382294 165678 382350
rect 165250 382170 165306 382226
rect 165374 382170 165430 382226
rect 165498 382170 165554 382226
rect 165622 382170 165678 382226
rect 165250 382046 165306 382102
rect 165374 382046 165430 382102
rect 165498 382046 165554 382102
rect 165622 382046 165678 382102
rect 165250 381922 165306 381978
rect 165374 381922 165430 381978
rect 165498 381922 165554 381978
rect 165622 381922 165678 381978
rect 165250 364294 165306 364350
rect 165374 364294 165430 364350
rect 165498 364294 165554 364350
rect 165622 364294 165678 364350
rect 165250 364170 165306 364226
rect 165374 364170 165430 364226
rect 165498 364170 165554 364226
rect 165622 364170 165678 364226
rect 165250 364046 165306 364102
rect 165374 364046 165430 364102
rect 165498 364046 165554 364102
rect 165622 364046 165678 364102
rect 165250 363922 165306 363978
rect 165374 363922 165430 363978
rect 165498 363922 165554 363978
rect 165622 363922 165678 363978
rect 165250 346294 165306 346350
rect 165374 346294 165430 346350
rect 165498 346294 165554 346350
rect 165622 346294 165678 346350
rect 165250 346170 165306 346226
rect 165374 346170 165430 346226
rect 165498 346170 165554 346226
rect 165622 346170 165678 346226
rect 165250 346046 165306 346102
rect 165374 346046 165430 346102
rect 165498 346046 165554 346102
rect 165622 346046 165678 346102
rect 165250 345922 165306 345978
rect 165374 345922 165430 345978
rect 165498 345922 165554 345978
rect 165622 345922 165678 345978
rect 165250 328294 165306 328350
rect 165374 328294 165430 328350
rect 165498 328294 165554 328350
rect 165622 328294 165678 328350
rect 165250 328170 165306 328226
rect 165374 328170 165430 328226
rect 165498 328170 165554 328226
rect 165622 328170 165678 328226
rect 165250 328046 165306 328102
rect 165374 328046 165430 328102
rect 165498 328046 165554 328102
rect 165622 328046 165678 328102
rect 165250 327922 165306 327978
rect 165374 327922 165430 327978
rect 165498 327922 165554 327978
rect 165622 327922 165678 327978
rect 165250 310294 165306 310350
rect 165374 310294 165430 310350
rect 165498 310294 165554 310350
rect 165622 310294 165678 310350
rect 165250 310170 165306 310226
rect 165374 310170 165430 310226
rect 165498 310170 165554 310226
rect 165622 310170 165678 310226
rect 165250 310046 165306 310102
rect 165374 310046 165430 310102
rect 165498 310046 165554 310102
rect 165622 310046 165678 310102
rect 165250 309922 165306 309978
rect 165374 309922 165430 309978
rect 165498 309922 165554 309978
rect 165622 309922 165678 309978
rect 165250 292294 165306 292350
rect 165374 292294 165430 292350
rect 165498 292294 165554 292350
rect 165622 292294 165678 292350
rect 165250 292170 165306 292226
rect 165374 292170 165430 292226
rect 165498 292170 165554 292226
rect 165622 292170 165678 292226
rect 165250 292046 165306 292102
rect 165374 292046 165430 292102
rect 165498 292046 165554 292102
rect 165622 292046 165678 292102
rect 165250 291922 165306 291978
rect 165374 291922 165430 291978
rect 165498 291922 165554 291978
rect 165622 291922 165678 291978
rect 165250 274294 165306 274350
rect 165374 274294 165430 274350
rect 165498 274294 165554 274350
rect 165622 274294 165678 274350
rect 165250 274170 165306 274226
rect 165374 274170 165430 274226
rect 165498 274170 165554 274226
rect 165622 274170 165678 274226
rect 165250 274046 165306 274102
rect 165374 274046 165430 274102
rect 165498 274046 165554 274102
rect 165622 274046 165678 274102
rect 165250 273922 165306 273978
rect 165374 273922 165430 273978
rect 165498 273922 165554 273978
rect 165622 273922 165678 273978
rect 165250 256294 165306 256350
rect 165374 256294 165430 256350
rect 165498 256294 165554 256350
rect 165622 256294 165678 256350
rect 165250 256170 165306 256226
rect 165374 256170 165430 256226
rect 165498 256170 165554 256226
rect 165622 256170 165678 256226
rect 165250 256046 165306 256102
rect 165374 256046 165430 256102
rect 165498 256046 165554 256102
rect 165622 256046 165678 256102
rect 165250 255922 165306 255978
rect 165374 255922 165430 255978
rect 165498 255922 165554 255978
rect 165622 255922 165678 255978
rect 165250 238294 165306 238350
rect 165374 238294 165430 238350
rect 165498 238294 165554 238350
rect 165622 238294 165678 238350
rect 165250 238170 165306 238226
rect 165374 238170 165430 238226
rect 165498 238170 165554 238226
rect 165622 238170 165678 238226
rect 165250 238046 165306 238102
rect 165374 238046 165430 238102
rect 165498 238046 165554 238102
rect 165622 238046 165678 238102
rect 165250 237922 165306 237978
rect 165374 237922 165430 237978
rect 165498 237922 165554 237978
rect 165622 237922 165678 237978
rect 165250 220294 165306 220350
rect 165374 220294 165430 220350
rect 165498 220294 165554 220350
rect 165622 220294 165678 220350
rect 165250 220170 165306 220226
rect 165374 220170 165430 220226
rect 165498 220170 165554 220226
rect 165622 220170 165678 220226
rect 165250 220046 165306 220102
rect 165374 220046 165430 220102
rect 165498 220046 165554 220102
rect 165622 220046 165678 220102
rect 165250 219922 165306 219978
rect 165374 219922 165430 219978
rect 165498 219922 165554 219978
rect 165622 219922 165678 219978
rect 165250 202294 165306 202350
rect 165374 202294 165430 202350
rect 165498 202294 165554 202350
rect 165622 202294 165678 202350
rect 165250 202170 165306 202226
rect 165374 202170 165430 202226
rect 165498 202170 165554 202226
rect 165622 202170 165678 202226
rect 165250 202046 165306 202102
rect 165374 202046 165430 202102
rect 165498 202046 165554 202102
rect 165622 202046 165678 202102
rect 165250 201922 165306 201978
rect 165374 201922 165430 201978
rect 165498 201922 165554 201978
rect 165622 201922 165678 201978
rect 165250 184294 165306 184350
rect 165374 184294 165430 184350
rect 165498 184294 165554 184350
rect 165622 184294 165678 184350
rect 165250 184170 165306 184226
rect 165374 184170 165430 184226
rect 165498 184170 165554 184226
rect 165622 184170 165678 184226
rect 165250 184046 165306 184102
rect 165374 184046 165430 184102
rect 165498 184046 165554 184102
rect 165622 184046 165678 184102
rect 165250 183922 165306 183978
rect 165374 183922 165430 183978
rect 165498 183922 165554 183978
rect 165622 183922 165678 183978
rect 165250 166294 165306 166350
rect 165374 166294 165430 166350
rect 165498 166294 165554 166350
rect 165622 166294 165678 166350
rect 165250 166170 165306 166226
rect 165374 166170 165430 166226
rect 165498 166170 165554 166226
rect 165622 166170 165678 166226
rect 165250 166046 165306 166102
rect 165374 166046 165430 166102
rect 165498 166046 165554 166102
rect 165622 166046 165678 166102
rect 165250 165922 165306 165978
rect 165374 165922 165430 165978
rect 165498 165922 165554 165978
rect 165622 165922 165678 165978
rect 165250 148294 165306 148350
rect 165374 148294 165430 148350
rect 165498 148294 165554 148350
rect 165622 148294 165678 148350
rect 165250 148170 165306 148226
rect 165374 148170 165430 148226
rect 165498 148170 165554 148226
rect 165622 148170 165678 148226
rect 165250 148046 165306 148102
rect 165374 148046 165430 148102
rect 165498 148046 165554 148102
rect 165622 148046 165678 148102
rect 165250 147922 165306 147978
rect 165374 147922 165430 147978
rect 165498 147922 165554 147978
rect 165622 147922 165678 147978
rect 165250 130294 165306 130350
rect 165374 130294 165430 130350
rect 165498 130294 165554 130350
rect 165622 130294 165678 130350
rect 165250 130170 165306 130226
rect 165374 130170 165430 130226
rect 165498 130170 165554 130226
rect 165622 130170 165678 130226
rect 165250 130046 165306 130102
rect 165374 130046 165430 130102
rect 165498 130046 165554 130102
rect 165622 130046 165678 130102
rect 165250 129922 165306 129978
rect 165374 129922 165430 129978
rect 165498 129922 165554 129978
rect 165622 129922 165678 129978
rect 165250 112294 165306 112350
rect 165374 112294 165430 112350
rect 165498 112294 165554 112350
rect 165622 112294 165678 112350
rect 165250 112170 165306 112226
rect 165374 112170 165430 112226
rect 165498 112170 165554 112226
rect 165622 112170 165678 112226
rect 165250 112046 165306 112102
rect 165374 112046 165430 112102
rect 165498 112046 165554 112102
rect 165622 112046 165678 112102
rect 165250 111922 165306 111978
rect 165374 111922 165430 111978
rect 165498 111922 165554 111978
rect 165622 111922 165678 111978
rect 165250 94294 165306 94350
rect 165374 94294 165430 94350
rect 165498 94294 165554 94350
rect 165622 94294 165678 94350
rect 165250 94170 165306 94226
rect 165374 94170 165430 94226
rect 165498 94170 165554 94226
rect 165622 94170 165678 94226
rect 165250 94046 165306 94102
rect 165374 94046 165430 94102
rect 165498 94046 165554 94102
rect 165622 94046 165678 94102
rect 165250 93922 165306 93978
rect 165374 93922 165430 93978
rect 165498 93922 165554 93978
rect 165622 93922 165678 93978
rect 165250 76294 165306 76350
rect 165374 76294 165430 76350
rect 165498 76294 165554 76350
rect 165622 76294 165678 76350
rect 165250 76170 165306 76226
rect 165374 76170 165430 76226
rect 165498 76170 165554 76226
rect 165622 76170 165678 76226
rect 165250 76046 165306 76102
rect 165374 76046 165430 76102
rect 165498 76046 165554 76102
rect 165622 76046 165678 76102
rect 165250 75922 165306 75978
rect 165374 75922 165430 75978
rect 165498 75922 165554 75978
rect 165622 75922 165678 75978
rect 165250 58294 165306 58350
rect 165374 58294 165430 58350
rect 165498 58294 165554 58350
rect 165622 58294 165678 58350
rect 165250 58170 165306 58226
rect 165374 58170 165430 58226
rect 165498 58170 165554 58226
rect 165622 58170 165678 58226
rect 165250 58046 165306 58102
rect 165374 58046 165430 58102
rect 165498 58046 165554 58102
rect 165622 58046 165678 58102
rect 165250 57922 165306 57978
rect 165374 57922 165430 57978
rect 165498 57922 165554 57978
rect 165622 57922 165678 57978
rect 165250 40294 165306 40350
rect 165374 40294 165430 40350
rect 165498 40294 165554 40350
rect 165622 40294 165678 40350
rect 165250 40170 165306 40226
rect 165374 40170 165430 40226
rect 165498 40170 165554 40226
rect 165622 40170 165678 40226
rect 165250 40046 165306 40102
rect 165374 40046 165430 40102
rect 165498 40046 165554 40102
rect 165622 40046 165678 40102
rect 165250 39922 165306 39978
rect 165374 39922 165430 39978
rect 165498 39922 165554 39978
rect 165622 39922 165678 39978
rect 165250 22294 165306 22350
rect 165374 22294 165430 22350
rect 165498 22294 165554 22350
rect 165622 22294 165678 22350
rect 165250 22170 165306 22226
rect 165374 22170 165430 22226
rect 165498 22170 165554 22226
rect 165622 22170 165678 22226
rect 165250 22046 165306 22102
rect 165374 22046 165430 22102
rect 165498 22046 165554 22102
rect 165622 22046 165678 22102
rect 165250 21922 165306 21978
rect 165374 21922 165430 21978
rect 165498 21922 165554 21978
rect 165622 21922 165678 21978
rect 165250 4294 165306 4350
rect 165374 4294 165430 4350
rect 165498 4294 165554 4350
rect 165622 4294 165678 4350
rect 165250 4170 165306 4226
rect 165374 4170 165430 4226
rect 165498 4170 165554 4226
rect 165622 4170 165678 4226
rect 165250 4046 165306 4102
rect 165374 4046 165430 4102
rect 165498 4046 165554 4102
rect 165622 4046 165678 4102
rect 165250 3922 165306 3978
rect 165374 3922 165430 3978
rect 165498 3922 165554 3978
rect 165622 3922 165678 3978
rect 165250 -216 165306 -160
rect 165374 -216 165430 -160
rect 165498 -216 165554 -160
rect 165622 -216 165678 -160
rect 165250 -340 165306 -284
rect 165374 -340 165430 -284
rect 165498 -340 165554 -284
rect 165622 -340 165678 -284
rect 165250 -464 165306 -408
rect 165374 -464 165430 -408
rect 165498 -464 165554 -408
rect 165622 -464 165678 -408
rect 165250 -588 165306 -532
rect 165374 -588 165430 -532
rect 165498 -588 165554 -532
rect 165622 -588 165678 -532
rect 168970 598116 169026 598172
rect 169094 598116 169150 598172
rect 169218 598116 169274 598172
rect 169342 598116 169398 598172
rect 168970 597992 169026 598048
rect 169094 597992 169150 598048
rect 169218 597992 169274 598048
rect 169342 597992 169398 598048
rect 168970 597868 169026 597924
rect 169094 597868 169150 597924
rect 169218 597868 169274 597924
rect 169342 597868 169398 597924
rect 168970 597744 169026 597800
rect 169094 597744 169150 597800
rect 169218 597744 169274 597800
rect 169342 597744 169398 597800
rect 168970 586294 169026 586350
rect 169094 586294 169150 586350
rect 169218 586294 169274 586350
rect 169342 586294 169398 586350
rect 168970 586170 169026 586226
rect 169094 586170 169150 586226
rect 169218 586170 169274 586226
rect 169342 586170 169398 586226
rect 168970 586046 169026 586102
rect 169094 586046 169150 586102
rect 169218 586046 169274 586102
rect 169342 586046 169398 586102
rect 168970 585922 169026 585978
rect 169094 585922 169150 585978
rect 169218 585922 169274 585978
rect 169342 585922 169398 585978
rect 168970 568294 169026 568350
rect 169094 568294 169150 568350
rect 169218 568294 169274 568350
rect 169342 568294 169398 568350
rect 168970 568170 169026 568226
rect 169094 568170 169150 568226
rect 169218 568170 169274 568226
rect 169342 568170 169398 568226
rect 168970 568046 169026 568102
rect 169094 568046 169150 568102
rect 169218 568046 169274 568102
rect 169342 568046 169398 568102
rect 168970 567922 169026 567978
rect 169094 567922 169150 567978
rect 169218 567922 169274 567978
rect 169342 567922 169398 567978
rect 168970 550294 169026 550350
rect 169094 550294 169150 550350
rect 169218 550294 169274 550350
rect 169342 550294 169398 550350
rect 168970 550170 169026 550226
rect 169094 550170 169150 550226
rect 169218 550170 169274 550226
rect 169342 550170 169398 550226
rect 168970 550046 169026 550102
rect 169094 550046 169150 550102
rect 169218 550046 169274 550102
rect 169342 550046 169398 550102
rect 168970 549922 169026 549978
rect 169094 549922 169150 549978
rect 169218 549922 169274 549978
rect 169342 549922 169398 549978
rect 168970 532294 169026 532350
rect 169094 532294 169150 532350
rect 169218 532294 169274 532350
rect 169342 532294 169398 532350
rect 168970 532170 169026 532226
rect 169094 532170 169150 532226
rect 169218 532170 169274 532226
rect 169342 532170 169398 532226
rect 168970 532046 169026 532102
rect 169094 532046 169150 532102
rect 169218 532046 169274 532102
rect 169342 532046 169398 532102
rect 168970 531922 169026 531978
rect 169094 531922 169150 531978
rect 169218 531922 169274 531978
rect 169342 531922 169398 531978
rect 168970 514294 169026 514350
rect 169094 514294 169150 514350
rect 169218 514294 169274 514350
rect 169342 514294 169398 514350
rect 168970 514170 169026 514226
rect 169094 514170 169150 514226
rect 169218 514170 169274 514226
rect 169342 514170 169398 514226
rect 168970 514046 169026 514102
rect 169094 514046 169150 514102
rect 169218 514046 169274 514102
rect 169342 514046 169398 514102
rect 168970 513922 169026 513978
rect 169094 513922 169150 513978
rect 169218 513922 169274 513978
rect 169342 513922 169398 513978
rect 168970 496294 169026 496350
rect 169094 496294 169150 496350
rect 169218 496294 169274 496350
rect 169342 496294 169398 496350
rect 168970 496170 169026 496226
rect 169094 496170 169150 496226
rect 169218 496170 169274 496226
rect 169342 496170 169398 496226
rect 168970 496046 169026 496102
rect 169094 496046 169150 496102
rect 169218 496046 169274 496102
rect 169342 496046 169398 496102
rect 168970 495922 169026 495978
rect 169094 495922 169150 495978
rect 169218 495922 169274 495978
rect 169342 495922 169398 495978
rect 168970 478294 169026 478350
rect 169094 478294 169150 478350
rect 169218 478294 169274 478350
rect 169342 478294 169398 478350
rect 168970 478170 169026 478226
rect 169094 478170 169150 478226
rect 169218 478170 169274 478226
rect 169342 478170 169398 478226
rect 168970 478046 169026 478102
rect 169094 478046 169150 478102
rect 169218 478046 169274 478102
rect 169342 478046 169398 478102
rect 168970 477922 169026 477978
rect 169094 477922 169150 477978
rect 169218 477922 169274 477978
rect 169342 477922 169398 477978
rect 168970 460294 169026 460350
rect 169094 460294 169150 460350
rect 169218 460294 169274 460350
rect 169342 460294 169398 460350
rect 168970 460170 169026 460226
rect 169094 460170 169150 460226
rect 169218 460170 169274 460226
rect 169342 460170 169398 460226
rect 168970 460046 169026 460102
rect 169094 460046 169150 460102
rect 169218 460046 169274 460102
rect 169342 460046 169398 460102
rect 168970 459922 169026 459978
rect 169094 459922 169150 459978
rect 169218 459922 169274 459978
rect 169342 459922 169398 459978
rect 168970 442294 169026 442350
rect 169094 442294 169150 442350
rect 169218 442294 169274 442350
rect 169342 442294 169398 442350
rect 168970 442170 169026 442226
rect 169094 442170 169150 442226
rect 169218 442170 169274 442226
rect 169342 442170 169398 442226
rect 168970 442046 169026 442102
rect 169094 442046 169150 442102
rect 169218 442046 169274 442102
rect 169342 442046 169398 442102
rect 168970 441922 169026 441978
rect 169094 441922 169150 441978
rect 169218 441922 169274 441978
rect 169342 441922 169398 441978
rect 168970 424294 169026 424350
rect 169094 424294 169150 424350
rect 169218 424294 169274 424350
rect 169342 424294 169398 424350
rect 168970 424170 169026 424226
rect 169094 424170 169150 424226
rect 169218 424170 169274 424226
rect 169342 424170 169398 424226
rect 168970 424046 169026 424102
rect 169094 424046 169150 424102
rect 169218 424046 169274 424102
rect 169342 424046 169398 424102
rect 168970 423922 169026 423978
rect 169094 423922 169150 423978
rect 169218 423922 169274 423978
rect 169342 423922 169398 423978
rect 168970 406294 169026 406350
rect 169094 406294 169150 406350
rect 169218 406294 169274 406350
rect 169342 406294 169398 406350
rect 168970 406170 169026 406226
rect 169094 406170 169150 406226
rect 169218 406170 169274 406226
rect 169342 406170 169398 406226
rect 168970 406046 169026 406102
rect 169094 406046 169150 406102
rect 169218 406046 169274 406102
rect 169342 406046 169398 406102
rect 168970 405922 169026 405978
rect 169094 405922 169150 405978
rect 169218 405922 169274 405978
rect 169342 405922 169398 405978
rect 168970 388294 169026 388350
rect 169094 388294 169150 388350
rect 169218 388294 169274 388350
rect 169342 388294 169398 388350
rect 168970 388170 169026 388226
rect 169094 388170 169150 388226
rect 169218 388170 169274 388226
rect 169342 388170 169398 388226
rect 168970 388046 169026 388102
rect 169094 388046 169150 388102
rect 169218 388046 169274 388102
rect 169342 388046 169398 388102
rect 168970 387922 169026 387978
rect 169094 387922 169150 387978
rect 169218 387922 169274 387978
rect 169342 387922 169398 387978
rect 168970 370294 169026 370350
rect 169094 370294 169150 370350
rect 169218 370294 169274 370350
rect 169342 370294 169398 370350
rect 168970 370170 169026 370226
rect 169094 370170 169150 370226
rect 169218 370170 169274 370226
rect 169342 370170 169398 370226
rect 168970 370046 169026 370102
rect 169094 370046 169150 370102
rect 169218 370046 169274 370102
rect 169342 370046 169398 370102
rect 168970 369922 169026 369978
rect 169094 369922 169150 369978
rect 169218 369922 169274 369978
rect 169342 369922 169398 369978
rect 168970 352294 169026 352350
rect 169094 352294 169150 352350
rect 169218 352294 169274 352350
rect 169342 352294 169398 352350
rect 168970 352170 169026 352226
rect 169094 352170 169150 352226
rect 169218 352170 169274 352226
rect 169342 352170 169398 352226
rect 168970 352046 169026 352102
rect 169094 352046 169150 352102
rect 169218 352046 169274 352102
rect 169342 352046 169398 352102
rect 168970 351922 169026 351978
rect 169094 351922 169150 351978
rect 169218 351922 169274 351978
rect 169342 351922 169398 351978
rect 168970 334294 169026 334350
rect 169094 334294 169150 334350
rect 169218 334294 169274 334350
rect 169342 334294 169398 334350
rect 168970 334170 169026 334226
rect 169094 334170 169150 334226
rect 169218 334170 169274 334226
rect 169342 334170 169398 334226
rect 168970 334046 169026 334102
rect 169094 334046 169150 334102
rect 169218 334046 169274 334102
rect 169342 334046 169398 334102
rect 168970 333922 169026 333978
rect 169094 333922 169150 333978
rect 169218 333922 169274 333978
rect 169342 333922 169398 333978
rect 168970 316294 169026 316350
rect 169094 316294 169150 316350
rect 169218 316294 169274 316350
rect 169342 316294 169398 316350
rect 168970 316170 169026 316226
rect 169094 316170 169150 316226
rect 169218 316170 169274 316226
rect 169342 316170 169398 316226
rect 168970 316046 169026 316102
rect 169094 316046 169150 316102
rect 169218 316046 169274 316102
rect 169342 316046 169398 316102
rect 168970 315922 169026 315978
rect 169094 315922 169150 315978
rect 169218 315922 169274 315978
rect 169342 315922 169398 315978
rect 168970 298294 169026 298350
rect 169094 298294 169150 298350
rect 169218 298294 169274 298350
rect 169342 298294 169398 298350
rect 168970 298170 169026 298226
rect 169094 298170 169150 298226
rect 169218 298170 169274 298226
rect 169342 298170 169398 298226
rect 168970 298046 169026 298102
rect 169094 298046 169150 298102
rect 169218 298046 169274 298102
rect 169342 298046 169398 298102
rect 168970 297922 169026 297978
rect 169094 297922 169150 297978
rect 169218 297922 169274 297978
rect 169342 297922 169398 297978
rect 168970 280294 169026 280350
rect 169094 280294 169150 280350
rect 169218 280294 169274 280350
rect 169342 280294 169398 280350
rect 168970 280170 169026 280226
rect 169094 280170 169150 280226
rect 169218 280170 169274 280226
rect 169342 280170 169398 280226
rect 168970 280046 169026 280102
rect 169094 280046 169150 280102
rect 169218 280046 169274 280102
rect 169342 280046 169398 280102
rect 168970 279922 169026 279978
rect 169094 279922 169150 279978
rect 169218 279922 169274 279978
rect 169342 279922 169398 279978
rect 168970 262294 169026 262350
rect 169094 262294 169150 262350
rect 169218 262294 169274 262350
rect 169342 262294 169398 262350
rect 168970 262170 169026 262226
rect 169094 262170 169150 262226
rect 169218 262170 169274 262226
rect 169342 262170 169398 262226
rect 168970 262046 169026 262102
rect 169094 262046 169150 262102
rect 169218 262046 169274 262102
rect 169342 262046 169398 262102
rect 168970 261922 169026 261978
rect 169094 261922 169150 261978
rect 169218 261922 169274 261978
rect 169342 261922 169398 261978
rect 168970 244294 169026 244350
rect 169094 244294 169150 244350
rect 169218 244294 169274 244350
rect 169342 244294 169398 244350
rect 168970 244170 169026 244226
rect 169094 244170 169150 244226
rect 169218 244170 169274 244226
rect 169342 244170 169398 244226
rect 168970 244046 169026 244102
rect 169094 244046 169150 244102
rect 169218 244046 169274 244102
rect 169342 244046 169398 244102
rect 168970 243922 169026 243978
rect 169094 243922 169150 243978
rect 169218 243922 169274 243978
rect 169342 243922 169398 243978
rect 168970 226294 169026 226350
rect 169094 226294 169150 226350
rect 169218 226294 169274 226350
rect 169342 226294 169398 226350
rect 168970 226170 169026 226226
rect 169094 226170 169150 226226
rect 169218 226170 169274 226226
rect 169342 226170 169398 226226
rect 168970 226046 169026 226102
rect 169094 226046 169150 226102
rect 169218 226046 169274 226102
rect 169342 226046 169398 226102
rect 168970 225922 169026 225978
rect 169094 225922 169150 225978
rect 169218 225922 169274 225978
rect 169342 225922 169398 225978
rect 168970 208294 169026 208350
rect 169094 208294 169150 208350
rect 169218 208294 169274 208350
rect 169342 208294 169398 208350
rect 168970 208170 169026 208226
rect 169094 208170 169150 208226
rect 169218 208170 169274 208226
rect 169342 208170 169398 208226
rect 168970 208046 169026 208102
rect 169094 208046 169150 208102
rect 169218 208046 169274 208102
rect 169342 208046 169398 208102
rect 168970 207922 169026 207978
rect 169094 207922 169150 207978
rect 169218 207922 169274 207978
rect 169342 207922 169398 207978
rect 168970 190294 169026 190350
rect 169094 190294 169150 190350
rect 169218 190294 169274 190350
rect 169342 190294 169398 190350
rect 168970 190170 169026 190226
rect 169094 190170 169150 190226
rect 169218 190170 169274 190226
rect 169342 190170 169398 190226
rect 168970 190046 169026 190102
rect 169094 190046 169150 190102
rect 169218 190046 169274 190102
rect 169342 190046 169398 190102
rect 168970 189922 169026 189978
rect 169094 189922 169150 189978
rect 169218 189922 169274 189978
rect 169342 189922 169398 189978
rect 168970 172294 169026 172350
rect 169094 172294 169150 172350
rect 169218 172294 169274 172350
rect 169342 172294 169398 172350
rect 168970 172170 169026 172226
rect 169094 172170 169150 172226
rect 169218 172170 169274 172226
rect 169342 172170 169398 172226
rect 168970 172046 169026 172102
rect 169094 172046 169150 172102
rect 169218 172046 169274 172102
rect 169342 172046 169398 172102
rect 168970 171922 169026 171978
rect 169094 171922 169150 171978
rect 169218 171922 169274 171978
rect 169342 171922 169398 171978
rect 168970 154294 169026 154350
rect 169094 154294 169150 154350
rect 169218 154294 169274 154350
rect 169342 154294 169398 154350
rect 168970 154170 169026 154226
rect 169094 154170 169150 154226
rect 169218 154170 169274 154226
rect 169342 154170 169398 154226
rect 168970 154046 169026 154102
rect 169094 154046 169150 154102
rect 169218 154046 169274 154102
rect 169342 154046 169398 154102
rect 168970 153922 169026 153978
rect 169094 153922 169150 153978
rect 169218 153922 169274 153978
rect 169342 153922 169398 153978
rect 168970 136294 169026 136350
rect 169094 136294 169150 136350
rect 169218 136294 169274 136350
rect 169342 136294 169398 136350
rect 168970 136170 169026 136226
rect 169094 136170 169150 136226
rect 169218 136170 169274 136226
rect 169342 136170 169398 136226
rect 168970 136046 169026 136102
rect 169094 136046 169150 136102
rect 169218 136046 169274 136102
rect 169342 136046 169398 136102
rect 168970 135922 169026 135978
rect 169094 135922 169150 135978
rect 169218 135922 169274 135978
rect 169342 135922 169398 135978
rect 168970 118294 169026 118350
rect 169094 118294 169150 118350
rect 169218 118294 169274 118350
rect 169342 118294 169398 118350
rect 168970 118170 169026 118226
rect 169094 118170 169150 118226
rect 169218 118170 169274 118226
rect 169342 118170 169398 118226
rect 168970 118046 169026 118102
rect 169094 118046 169150 118102
rect 169218 118046 169274 118102
rect 169342 118046 169398 118102
rect 168970 117922 169026 117978
rect 169094 117922 169150 117978
rect 169218 117922 169274 117978
rect 169342 117922 169398 117978
rect 168970 100294 169026 100350
rect 169094 100294 169150 100350
rect 169218 100294 169274 100350
rect 169342 100294 169398 100350
rect 168970 100170 169026 100226
rect 169094 100170 169150 100226
rect 169218 100170 169274 100226
rect 169342 100170 169398 100226
rect 168970 100046 169026 100102
rect 169094 100046 169150 100102
rect 169218 100046 169274 100102
rect 169342 100046 169398 100102
rect 168970 99922 169026 99978
rect 169094 99922 169150 99978
rect 169218 99922 169274 99978
rect 169342 99922 169398 99978
rect 168970 82294 169026 82350
rect 169094 82294 169150 82350
rect 169218 82294 169274 82350
rect 169342 82294 169398 82350
rect 168970 82170 169026 82226
rect 169094 82170 169150 82226
rect 169218 82170 169274 82226
rect 169342 82170 169398 82226
rect 168970 82046 169026 82102
rect 169094 82046 169150 82102
rect 169218 82046 169274 82102
rect 169342 82046 169398 82102
rect 168970 81922 169026 81978
rect 169094 81922 169150 81978
rect 169218 81922 169274 81978
rect 169342 81922 169398 81978
rect 168970 64294 169026 64350
rect 169094 64294 169150 64350
rect 169218 64294 169274 64350
rect 169342 64294 169398 64350
rect 168970 64170 169026 64226
rect 169094 64170 169150 64226
rect 169218 64170 169274 64226
rect 169342 64170 169398 64226
rect 168970 64046 169026 64102
rect 169094 64046 169150 64102
rect 169218 64046 169274 64102
rect 169342 64046 169398 64102
rect 168970 63922 169026 63978
rect 169094 63922 169150 63978
rect 169218 63922 169274 63978
rect 169342 63922 169398 63978
rect 168970 46294 169026 46350
rect 169094 46294 169150 46350
rect 169218 46294 169274 46350
rect 169342 46294 169398 46350
rect 168970 46170 169026 46226
rect 169094 46170 169150 46226
rect 169218 46170 169274 46226
rect 169342 46170 169398 46226
rect 168970 46046 169026 46102
rect 169094 46046 169150 46102
rect 169218 46046 169274 46102
rect 169342 46046 169398 46102
rect 168970 45922 169026 45978
rect 169094 45922 169150 45978
rect 169218 45922 169274 45978
rect 169342 45922 169398 45978
rect 168970 28294 169026 28350
rect 169094 28294 169150 28350
rect 169218 28294 169274 28350
rect 169342 28294 169398 28350
rect 168970 28170 169026 28226
rect 169094 28170 169150 28226
rect 169218 28170 169274 28226
rect 169342 28170 169398 28226
rect 168970 28046 169026 28102
rect 169094 28046 169150 28102
rect 169218 28046 169274 28102
rect 169342 28046 169398 28102
rect 168970 27922 169026 27978
rect 169094 27922 169150 27978
rect 169218 27922 169274 27978
rect 169342 27922 169398 27978
rect 168970 10294 169026 10350
rect 169094 10294 169150 10350
rect 169218 10294 169274 10350
rect 169342 10294 169398 10350
rect 168970 10170 169026 10226
rect 169094 10170 169150 10226
rect 169218 10170 169274 10226
rect 169342 10170 169398 10226
rect 168970 10046 169026 10102
rect 169094 10046 169150 10102
rect 169218 10046 169274 10102
rect 169342 10046 169398 10102
rect 168970 9922 169026 9978
rect 169094 9922 169150 9978
rect 169218 9922 169274 9978
rect 169342 9922 169398 9978
rect 168970 -1176 169026 -1120
rect 169094 -1176 169150 -1120
rect 169218 -1176 169274 -1120
rect 169342 -1176 169398 -1120
rect 168970 -1300 169026 -1244
rect 169094 -1300 169150 -1244
rect 169218 -1300 169274 -1244
rect 169342 -1300 169398 -1244
rect 168970 -1424 169026 -1368
rect 169094 -1424 169150 -1368
rect 169218 -1424 169274 -1368
rect 169342 -1424 169398 -1368
rect 168970 -1548 169026 -1492
rect 169094 -1548 169150 -1492
rect 169218 -1548 169274 -1492
rect 169342 -1548 169398 -1492
rect 183250 597156 183306 597212
rect 183374 597156 183430 597212
rect 183498 597156 183554 597212
rect 183622 597156 183678 597212
rect 183250 597032 183306 597088
rect 183374 597032 183430 597088
rect 183498 597032 183554 597088
rect 183622 597032 183678 597088
rect 183250 596908 183306 596964
rect 183374 596908 183430 596964
rect 183498 596908 183554 596964
rect 183622 596908 183678 596964
rect 183250 596784 183306 596840
rect 183374 596784 183430 596840
rect 183498 596784 183554 596840
rect 183622 596784 183678 596840
rect 183250 580294 183306 580350
rect 183374 580294 183430 580350
rect 183498 580294 183554 580350
rect 183622 580294 183678 580350
rect 183250 580170 183306 580226
rect 183374 580170 183430 580226
rect 183498 580170 183554 580226
rect 183622 580170 183678 580226
rect 183250 580046 183306 580102
rect 183374 580046 183430 580102
rect 183498 580046 183554 580102
rect 183622 580046 183678 580102
rect 183250 579922 183306 579978
rect 183374 579922 183430 579978
rect 183498 579922 183554 579978
rect 183622 579922 183678 579978
rect 183250 562294 183306 562350
rect 183374 562294 183430 562350
rect 183498 562294 183554 562350
rect 183622 562294 183678 562350
rect 183250 562170 183306 562226
rect 183374 562170 183430 562226
rect 183498 562170 183554 562226
rect 183622 562170 183678 562226
rect 183250 562046 183306 562102
rect 183374 562046 183430 562102
rect 183498 562046 183554 562102
rect 183622 562046 183678 562102
rect 183250 561922 183306 561978
rect 183374 561922 183430 561978
rect 183498 561922 183554 561978
rect 183622 561922 183678 561978
rect 183250 544294 183306 544350
rect 183374 544294 183430 544350
rect 183498 544294 183554 544350
rect 183622 544294 183678 544350
rect 183250 544170 183306 544226
rect 183374 544170 183430 544226
rect 183498 544170 183554 544226
rect 183622 544170 183678 544226
rect 183250 544046 183306 544102
rect 183374 544046 183430 544102
rect 183498 544046 183554 544102
rect 183622 544046 183678 544102
rect 183250 543922 183306 543978
rect 183374 543922 183430 543978
rect 183498 543922 183554 543978
rect 183622 543922 183678 543978
rect 183250 526294 183306 526350
rect 183374 526294 183430 526350
rect 183498 526294 183554 526350
rect 183622 526294 183678 526350
rect 183250 526170 183306 526226
rect 183374 526170 183430 526226
rect 183498 526170 183554 526226
rect 183622 526170 183678 526226
rect 183250 526046 183306 526102
rect 183374 526046 183430 526102
rect 183498 526046 183554 526102
rect 183622 526046 183678 526102
rect 183250 525922 183306 525978
rect 183374 525922 183430 525978
rect 183498 525922 183554 525978
rect 183622 525922 183678 525978
rect 183250 508294 183306 508350
rect 183374 508294 183430 508350
rect 183498 508294 183554 508350
rect 183622 508294 183678 508350
rect 183250 508170 183306 508226
rect 183374 508170 183430 508226
rect 183498 508170 183554 508226
rect 183622 508170 183678 508226
rect 183250 508046 183306 508102
rect 183374 508046 183430 508102
rect 183498 508046 183554 508102
rect 183622 508046 183678 508102
rect 183250 507922 183306 507978
rect 183374 507922 183430 507978
rect 183498 507922 183554 507978
rect 183622 507922 183678 507978
rect 183250 490294 183306 490350
rect 183374 490294 183430 490350
rect 183498 490294 183554 490350
rect 183622 490294 183678 490350
rect 183250 490170 183306 490226
rect 183374 490170 183430 490226
rect 183498 490170 183554 490226
rect 183622 490170 183678 490226
rect 183250 490046 183306 490102
rect 183374 490046 183430 490102
rect 183498 490046 183554 490102
rect 183622 490046 183678 490102
rect 183250 489922 183306 489978
rect 183374 489922 183430 489978
rect 183498 489922 183554 489978
rect 183622 489922 183678 489978
rect 183250 472294 183306 472350
rect 183374 472294 183430 472350
rect 183498 472294 183554 472350
rect 183622 472294 183678 472350
rect 183250 472170 183306 472226
rect 183374 472170 183430 472226
rect 183498 472170 183554 472226
rect 183622 472170 183678 472226
rect 183250 472046 183306 472102
rect 183374 472046 183430 472102
rect 183498 472046 183554 472102
rect 183622 472046 183678 472102
rect 183250 471922 183306 471978
rect 183374 471922 183430 471978
rect 183498 471922 183554 471978
rect 183622 471922 183678 471978
rect 183250 454294 183306 454350
rect 183374 454294 183430 454350
rect 183498 454294 183554 454350
rect 183622 454294 183678 454350
rect 183250 454170 183306 454226
rect 183374 454170 183430 454226
rect 183498 454170 183554 454226
rect 183622 454170 183678 454226
rect 183250 454046 183306 454102
rect 183374 454046 183430 454102
rect 183498 454046 183554 454102
rect 183622 454046 183678 454102
rect 183250 453922 183306 453978
rect 183374 453922 183430 453978
rect 183498 453922 183554 453978
rect 183622 453922 183678 453978
rect 183250 436294 183306 436350
rect 183374 436294 183430 436350
rect 183498 436294 183554 436350
rect 183622 436294 183678 436350
rect 183250 436170 183306 436226
rect 183374 436170 183430 436226
rect 183498 436170 183554 436226
rect 183622 436170 183678 436226
rect 183250 436046 183306 436102
rect 183374 436046 183430 436102
rect 183498 436046 183554 436102
rect 183622 436046 183678 436102
rect 183250 435922 183306 435978
rect 183374 435922 183430 435978
rect 183498 435922 183554 435978
rect 183622 435922 183678 435978
rect 183250 418294 183306 418350
rect 183374 418294 183430 418350
rect 183498 418294 183554 418350
rect 183622 418294 183678 418350
rect 183250 418170 183306 418226
rect 183374 418170 183430 418226
rect 183498 418170 183554 418226
rect 183622 418170 183678 418226
rect 183250 418046 183306 418102
rect 183374 418046 183430 418102
rect 183498 418046 183554 418102
rect 183622 418046 183678 418102
rect 183250 417922 183306 417978
rect 183374 417922 183430 417978
rect 183498 417922 183554 417978
rect 183622 417922 183678 417978
rect 183250 400294 183306 400350
rect 183374 400294 183430 400350
rect 183498 400294 183554 400350
rect 183622 400294 183678 400350
rect 183250 400170 183306 400226
rect 183374 400170 183430 400226
rect 183498 400170 183554 400226
rect 183622 400170 183678 400226
rect 183250 400046 183306 400102
rect 183374 400046 183430 400102
rect 183498 400046 183554 400102
rect 183622 400046 183678 400102
rect 183250 399922 183306 399978
rect 183374 399922 183430 399978
rect 183498 399922 183554 399978
rect 183622 399922 183678 399978
rect 183250 382294 183306 382350
rect 183374 382294 183430 382350
rect 183498 382294 183554 382350
rect 183622 382294 183678 382350
rect 183250 382170 183306 382226
rect 183374 382170 183430 382226
rect 183498 382170 183554 382226
rect 183622 382170 183678 382226
rect 183250 382046 183306 382102
rect 183374 382046 183430 382102
rect 183498 382046 183554 382102
rect 183622 382046 183678 382102
rect 183250 381922 183306 381978
rect 183374 381922 183430 381978
rect 183498 381922 183554 381978
rect 183622 381922 183678 381978
rect 183250 364294 183306 364350
rect 183374 364294 183430 364350
rect 183498 364294 183554 364350
rect 183622 364294 183678 364350
rect 183250 364170 183306 364226
rect 183374 364170 183430 364226
rect 183498 364170 183554 364226
rect 183622 364170 183678 364226
rect 183250 364046 183306 364102
rect 183374 364046 183430 364102
rect 183498 364046 183554 364102
rect 183622 364046 183678 364102
rect 183250 363922 183306 363978
rect 183374 363922 183430 363978
rect 183498 363922 183554 363978
rect 183622 363922 183678 363978
rect 183250 346294 183306 346350
rect 183374 346294 183430 346350
rect 183498 346294 183554 346350
rect 183622 346294 183678 346350
rect 183250 346170 183306 346226
rect 183374 346170 183430 346226
rect 183498 346170 183554 346226
rect 183622 346170 183678 346226
rect 183250 346046 183306 346102
rect 183374 346046 183430 346102
rect 183498 346046 183554 346102
rect 183622 346046 183678 346102
rect 183250 345922 183306 345978
rect 183374 345922 183430 345978
rect 183498 345922 183554 345978
rect 183622 345922 183678 345978
rect 183250 328294 183306 328350
rect 183374 328294 183430 328350
rect 183498 328294 183554 328350
rect 183622 328294 183678 328350
rect 183250 328170 183306 328226
rect 183374 328170 183430 328226
rect 183498 328170 183554 328226
rect 183622 328170 183678 328226
rect 183250 328046 183306 328102
rect 183374 328046 183430 328102
rect 183498 328046 183554 328102
rect 183622 328046 183678 328102
rect 183250 327922 183306 327978
rect 183374 327922 183430 327978
rect 183498 327922 183554 327978
rect 183622 327922 183678 327978
rect 183250 310294 183306 310350
rect 183374 310294 183430 310350
rect 183498 310294 183554 310350
rect 183622 310294 183678 310350
rect 183250 310170 183306 310226
rect 183374 310170 183430 310226
rect 183498 310170 183554 310226
rect 183622 310170 183678 310226
rect 183250 310046 183306 310102
rect 183374 310046 183430 310102
rect 183498 310046 183554 310102
rect 183622 310046 183678 310102
rect 183250 309922 183306 309978
rect 183374 309922 183430 309978
rect 183498 309922 183554 309978
rect 183622 309922 183678 309978
rect 183250 292294 183306 292350
rect 183374 292294 183430 292350
rect 183498 292294 183554 292350
rect 183622 292294 183678 292350
rect 183250 292170 183306 292226
rect 183374 292170 183430 292226
rect 183498 292170 183554 292226
rect 183622 292170 183678 292226
rect 183250 292046 183306 292102
rect 183374 292046 183430 292102
rect 183498 292046 183554 292102
rect 183622 292046 183678 292102
rect 183250 291922 183306 291978
rect 183374 291922 183430 291978
rect 183498 291922 183554 291978
rect 183622 291922 183678 291978
rect 183250 274294 183306 274350
rect 183374 274294 183430 274350
rect 183498 274294 183554 274350
rect 183622 274294 183678 274350
rect 183250 274170 183306 274226
rect 183374 274170 183430 274226
rect 183498 274170 183554 274226
rect 183622 274170 183678 274226
rect 183250 274046 183306 274102
rect 183374 274046 183430 274102
rect 183498 274046 183554 274102
rect 183622 274046 183678 274102
rect 183250 273922 183306 273978
rect 183374 273922 183430 273978
rect 183498 273922 183554 273978
rect 183622 273922 183678 273978
rect 183250 256294 183306 256350
rect 183374 256294 183430 256350
rect 183498 256294 183554 256350
rect 183622 256294 183678 256350
rect 183250 256170 183306 256226
rect 183374 256170 183430 256226
rect 183498 256170 183554 256226
rect 183622 256170 183678 256226
rect 183250 256046 183306 256102
rect 183374 256046 183430 256102
rect 183498 256046 183554 256102
rect 183622 256046 183678 256102
rect 183250 255922 183306 255978
rect 183374 255922 183430 255978
rect 183498 255922 183554 255978
rect 183622 255922 183678 255978
rect 183250 238294 183306 238350
rect 183374 238294 183430 238350
rect 183498 238294 183554 238350
rect 183622 238294 183678 238350
rect 183250 238170 183306 238226
rect 183374 238170 183430 238226
rect 183498 238170 183554 238226
rect 183622 238170 183678 238226
rect 183250 238046 183306 238102
rect 183374 238046 183430 238102
rect 183498 238046 183554 238102
rect 183622 238046 183678 238102
rect 183250 237922 183306 237978
rect 183374 237922 183430 237978
rect 183498 237922 183554 237978
rect 183622 237922 183678 237978
rect 183250 220294 183306 220350
rect 183374 220294 183430 220350
rect 183498 220294 183554 220350
rect 183622 220294 183678 220350
rect 183250 220170 183306 220226
rect 183374 220170 183430 220226
rect 183498 220170 183554 220226
rect 183622 220170 183678 220226
rect 183250 220046 183306 220102
rect 183374 220046 183430 220102
rect 183498 220046 183554 220102
rect 183622 220046 183678 220102
rect 183250 219922 183306 219978
rect 183374 219922 183430 219978
rect 183498 219922 183554 219978
rect 183622 219922 183678 219978
rect 183250 202294 183306 202350
rect 183374 202294 183430 202350
rect 183498 202294 183554 202350
rect 183622 202294 183678 202350
rect 183250 202170 183306 202226
rect 183374 202170 183430 202226
rect 183498 202170 183554 202226
rect 183622 202170 183678 202226
rect 183250 202046 183306 202102
rect 183374 202046 183430 202102
rect 183498 202046 183554 202102
rect 183622 202046 183678 202102
rect 183250 201922 183306 201978
rect 183374 201922 183430 201978
rect 183498 201922 183554 201978
rect 183622 201922 183678 201978
rect 183250 184294 183306 184350
rect 183374 184294 183430 184350
rect 183498 184294 183554 184350
rect 183622 184294 183678 184350
rect 183250 184170 183306 184226
rect 183374 184170 183430 184226
rect 183498 184170 183554 184226
rect 183622 184170 183678 184226
rect 183250 184046 183306 184102
rect 183374 184046 183430 184102
rect 183498 184046 183554 184102
rect 183622 184046 183678 184102
rect 183250 183922 183306 183978
rect 183374 183922 183430 183978
rect 183498 183922 183554 183978
rect 183622 183922 183678 183978
rect 183250 166294 183306 166350
rect 183374 166294 183430 166350
rect 183498 166294 183554 166350
rect 183622 166294 183678 166350
rect 183250 166170 183306 166226
rect 183374 166170 183430 166226
rect 183498 166170 183554 166226
rect 183622 166170 183678 166226
rect 183250 166046 183306 166102
rect 183374 166046 183430 166102
rect 183498 166046 183554 166102
rect 183622 166046 183678 166102
rect 183250 165922 183306 165978
rect 183374 165922 183430 165978
rect 183498 165922 183554 165978
rect 183622 165922 183678 165978
rect 183250 148294 183306 148350
rect 183374 148294 183430 148350
rect 183498 148294 183554 148350
rect 183622 148294 183678 148350
rect 183250 148170 183306 148226
rect 183374 148170 183430 148226
rect 183498 148170 183554 148226
rect 183622 148170 183678 148226
rect 183250 148046 183306 148102
rect 183374 148046 183430 148102
rect 183498 148046 183554 148102
rect 183622 148046 183678 148102
rect 183250 147922 183306 147978
rect 183374 147922 183430 147978
rect 183498 147922 183554 147978
rect 183622 147922 183678 147978
rect 183250 130294 183306 130350
rect 183374 130294 183430 130350
rect 183498 130294 183554 130350
rect 183622 130294 183678 130350
rect 183250 130170 183306 130226
rect 183374 130170 183430 130226
rect 183498 130170 183554 130226
rect 183622 130170 183678 130226
rect 183250 130046 183306 130102
rect 183374 130046 183430 130102
rect 183498 130046 183554 130102
rect 183622 130046 183678 130102
rect 183250 129922 183306 129978
rect 183374 129922 183430 129978
rect 183498 129922 183554 129978
rect 183622 129922 183678 129978
rect 183250 112294 183306 112350
rect 183374 112294 183430 112350
rect 183498 112294 183554 112350
rect 183622 112294 183678 112350
rect 183250 112170 183306 112226
rect 183374 112170 183430 112226
rect 183498 112170 183554 112226
rect 183622 112170 183678 112226
rect 183250 112046 183306 112102
rect 183374 112046 183430 112102
rect 183498 112046 183554 112102
rect 183622 112046 183678 112102
rect 183250 111922 183306 111978
rect 183374 111922 183430 111978
rect 183498 111922 183554 111978
rect 183622 111922 183678 111978
rect 183250 94294 183306 94350
rect 183374 94294 183430 94350
rect 183498 94294 183554 94350
rect 183622 94294 183678 94350
rect 183250 94170 183306 94226
rect 183374 94170 183430 94226
rect 183498 94170 183554 94226
rect 183622 94170 183678 94226
rect 183250 94046 183306 94102
rect 183374 94046 183430 94102
rect 183498 94046 183554 94102
rect 183622 94046 183678 94102
rect 183250 93922 183306 93978
rect 183374 93922 183430 93978
rect 183498 93922 183554 93978
rect 183622 93922 183678 93978
rect 183250 76294 183306 76350
rect 183374 76294 183430 76350
rect 183498 76294 183554 76350
rect 183622 76294 183678 76350
rect 183250 76170 183306 76226
rect 183374 76170 183430 76226
rect 183498 76170 183554 76226
rect 183622 76170 183678 76226
rect 183250 76046 183306 76102
rect 183374 76046 183430 76102
rect 183498 76046 183554 76102
rect 183622 76046 183678 76102
rect 183250 75922 183306 75978
rect 183374 75922 183430 75978
rect 183498 75922 183554 75978
rect 183622 75922 183678 75978
rect 183250 58294 183306 58350
rect 183374 58294 183430 58350
rect 183498 58294 183554 58350
rect 183622 58294 183678 58350
rect 183250 58170 183306 58226
rect 183374 58170 183430 58226
rect 183498 58170 183554 58226
rect 183622 58170 183678 58226
rect 183250 58046 183306 58102
rect 183374 58046 183430 58102
rect 183498 58046 183554 58102
rect 183622 58046 183678 58102
rect 183250 57922 183306 57978
rect 183374 57922 183430 57978
rect 183498 57922 183554 57978
rect 183622 57922 183678 57978
rect 183250 40294 183306 40350
rect 183374 40294 183430 40350
rect 183498 40294 183554 40350
rect 183622 40294 183678 40350
rect 183250 40170 183306 40226
rect 183374 40170 183430 40226
rect 183498 40170 183554 40226
rect 183622 40170 183678 40226
rect 183250 40046 183306 40102
rect 183374 40046 183430 40102
rect 183498 40046 183554 40102
rect 183622 40046 183678 40102
rect 183250 39922 183306 39978
rect 183374 39922 183430 39978
rect 183498 39922 183554 39978
rect 183622 39922 183678 39978
rect 183250 22294 183306 22350
rect 183374 22294 183430 22350
rect 183498 22294 183554 22350
rect 183622 22294 183678 22350
rect 183250 22170 183306 22226
rect 183374 22170 183430 22226
rect 183498 22170 183554 22226
rect 183622 22170 183678 22226
rect 183250 22046 183306 22102
rect 183374 22046 183430 22102
rect 183498 22046 183554 22102
rect 183622 22046 183678 22102
rect 183250 21922 183306 21978
rect 183374 21922 183430 21978
rect 183498 21922 183554 21978
rect 183622 21922 183678 21978
rect 183250 4294 183306 4350
rect 183374 4294 183430 4350
rect 183498 4294 183554 4350
rect 183622 4294 183678 4350
rect 183250 4170 183306 4226
rect 183374 4170 183430 4226
rect 183498 4170 183554 4226
rect 183622 4170 183678 4226
rect 183250 4046 183306 4102
rect 183374 4046 183430 4102
rect 183498 4046 183554 4102
rect 183622 4046 183678 4102
rect 183250 3922 183306 3978
rect 183374 3922 183430 3978
rect 183498 3922 183554 3978
rect 183622 3922 183678 3978
rect 183250 -216 183306 -160
rect 183374 -216 183430 -160
rect 183498 -216 183554 -160
rect 183622 -216 183678 -160
rect 183250 -340 183306 -284
rect 183374 -340 183430 -284
rect 183498 -340 183554 -284
rect 183622 -340 183678 -284
rect 183250 -464 183306 -408
rect 183374 -464 183430 -408
rect 183498 -464 183554 -408
rect 183622 -464 183678 -408
rect 183250 -588 183306 -532
rect 183374 -588 183430 -532
rect 183498 -588 183554 -532
rect 183622 -588 183678 -532
rect 186970 598116 187026 598172
rect 187094 598116 187150 598172
rect 187218 598116 187274 598172
rect 187342 598116 187398 598172
rect 186970 597992 187026 598048
rect 187094 597992 187150 598048
rect 187218 597992 187274 598048
rect 187342 597992 187398 598048
rect 186970 597868 187026 597924
rect 187094 597868 187150 597924
rect 187218 597868 187274 597924
rect 187342 597868 187398 597924
rect 186970 597744 187026 597800
rect 187094 597744 187150 597800
rect 187218 597744 187274 597800
rect 187342 597744 187398 597800
rect 186970 586294 187026 586350
rect 187094 586294 187150 586350
rect 187218 586294 187274 586350
rect 187342 586294 187398 586350
rect 186970 586170 187026 586226
rect 187094 586170 187150 586226
rect 187218 586170 187274 586226
rect 187342 586170 187398 586226
rect 186970 586046 187026 586102
rect 187094 586046 187150 586102
rect 187218 586046 187274 586102
rect 187342 586046 187398 586102
rect 186970 585922 187026 585978
rect 187094 585922 187150 585978
rect 187218 585922 187274 585978
rect 187342 585922 187398 585978
rect 186970 568294 187026 568350
rect 187094 568294 187150 568350
rect 187218 568294 187274 568350
rect 187342 568294 187398 568350
rect 186970 568170 187026 568226
rect 187094 568170 187150 568226
rect 187218 568170 187274 568226
rect 187342 568170 187398 568226
rect 186970 568046 187026 568102
rect 187094 568046 187150 568102
rect 187218 568046 187274 568102
rect 187342 568046 187398 568102
rect 186970 567922 187026 567978
rect 187094 567922 187150 567978
rect 187218 567922 187274 567978
rect 187342 567922 187398 567978
rect 186970 550294 187026 550350
rect 187094 550294 187150 550350
rect 187218 550294 187274 550350
rect 187342 550294 187398 550350
rect 186970 550170 187026 550226
rect 187094 550170 187150 550226
rect 187218 550170 187274 550226
rect 187342 550170 187398 550226
rect 186970 550046 187026 550102
rect 187094 550046 187150 550102
rect 187218 550046 187274 550102
rect 187342 550046 187398 550102
rect 186970 549922 187026 549978
rect 187094 549922 187150 549978
rect 187218 549922 187274 549978
rect 187342 549922 187398 549978
rect 186970 532294 187026 532350
rect 187094 532294 187150 532350
rect 187218 532294 187274 532350
rect 187342 532294 187398 532350
rect 186970 532170 187026 532226
rect 187094 532170 187150 532226
rect 187218 532170 187274 532226
rect 187342 532170 187398 532226
rect 186970 532046 187026 532102
rect 187094 532046 187150 532102
rect 187218 532046 187274 532102
rect 187342 532046 187398 532102
rect 186970 531922 187026 531978
rect 187094 531922 187150 531978
rect 187218 531922 187274 531978
rect 187342 531922 187398 531978
rect 186970 514294 187026 514350
rect 187094 514294 187150 514350
rect 187218 514294 187274 514350
rect 187342 514294 187398 514350
rect 186970 514170 187026 514226
rect 187094 514170 187150 514226
rect 187218 514170 187274 514226
rect 187342 514170 187398 514226
rect 186970 514046 187026 514102
rect 187094 514046 187150 514102
rect 187218 514046 187274 514102
rect 187342 514046 187398 514102
rect 186970 513922 187026 513978
rect 187094 513922 187150 513978
rect 187218 513922 187274 513978
rect 187342 513922 187398 513978
rect 186970 496294 187026 496350
rect 187094 496294 187150 496350
rect 187218 496294 187274 496350
rect 187342 496294 187398 496350
rect 186970 496170 187026 496226
rect 187094 496170 187150 496226
rect 187218 496170 187274 496226
rect 187342 496170 187398 496226
rect 186970 496046 187026 496102
rect 187094 496046 187150 496102
rect 187218 496046 187274 496102
rect 187342 496046 187398 496102
rect 186970 495922 187026 495978
rect 187094 495922 187150 495978
rect 187218 495922 187274 495978
rect 187342 495922 187398 495978
rect 186970 478294 187026 478350
rect 187094 478294 187150 478350
rect 187218 478294 187274 478350
rect 187342 478294 187398 478350
rect 186970 478170 187026 478226
rect 187094 478170 187150 478226
rect 187218 478170 187274 478226
rect 187342 478170 187398 478226
rect 186970 478046 187026 478102
rect 187094 478046 187150 478102
rect 187218 478046 187274 478102
rect 187342 478046 187398 478102
rect 186970 477922 187026 477978
rect 187094 477922 187150 477978
rect 187218 477922 187274 477978
rect 187342 477922 187398 477978
rect 186970 460294 187026 460350
rect 187094 460294 187150 460350
rect 187218 460294 187274 460350
rect 187342 460294 187398 460350
rect 186970 460170 187026 460226
rect 187094 460170 187150 460226
rect 187218 460170 187274 460226
rect 187342 460170 187398 460226
rect 186970 460046 187026 460102
rect 187094 460046 187150 460102
rect 187218 460046 187274 460102
rect 187342 460046 187398 460102
rect 186970 459922 187026 459978
rect 187094 459922 187150 459978
rect 187218 459922 187274 459978
rect 187342 459922 187398 459978
rect 186970 442294 187026 442350
rect 187094 442294 187150 442350
rect 187218 442294 187274 442350
rect 187342 442294 187398 442350
rect 186970 442170 187026 442226
rect 187094 442170 187150 442226
rect 187218 442170 187274 442226
rect 187342 442170 187398 442226
rect 186970 442046 187026 442102
rect 187094 442046 187150 442102
rect 187218 442046 187274 442102
rect 187342 442046 187398 442102
rect 186970 441922 187026 441978
rect 187094 441922 187150 441978
rect 187218 441922 187274 441978
rect 187342 441922 187398 441978
rect 186970 424294 187026 424350
rect 187094 424294 187150 424350
rect 187218 424294 187274 424350
rect 187342 424294 187398 424350
rect 186970 424170 187026 424226
rect 187094 424170 187150 424226
rect 187218 424170 187274 424226
rect 187342 424170 187398 424226
rect 186970 424046 187026 424102
rect 187094 424046 187150 424102
rect 187218 424046 187274 424102
rect 187342 424046 187398 424102
rect 186970 423922 187026 423978
rect 187094 423922 187150 423978
rect 187218 423922 187274 423978
rect 187342 423922 187398 423978
rect 186970 406294 187026 406350
rect 187094 406294 187150 406350
rect 187218 406294 187274 406350
rect 187342 406294 187398 406350
rect 186970 406170 187026 406226
rect 187094 406170 187150 406226
rect 187218 406170 187274 406226
rect 187342 406170 187398 406226
rect 186970 406046 187026 406102
rect 187094 406046 187150 406102
rect 187218 406046 187274 406102
rect 187342 406046 187398 406102
rect 186970 405922 187026 405978
rect 187094 405922 187150 405978
rect 187218 405922 187274 405978
rect 187342 405922 187398 405978
rect 186970 388294 187026 388350
rect 187094 388294 187150 388350
rect 187218 388294 187274 388350
rect 187342 388294 187398 388350
rect 186970 388170 187026 388226
rect 187094 388170 187150 388226
rect 187218 388170 187274 388226
rect 187342 388170 187398 388226
rect 186970 388046 187026 388102
rect 187094 388046 187150 388102
rect 187218 388046 187274 388102
rect 187342 388046 187398 388102
rect 186970 387922 187026 387978
rect 187094 387922 187150 387978
rect 187218 387922 187274 387978
rect 187342 387922 187398 387978
rect 186970 370294 187026 370350
rect 187094 370294 187150 370350
rect 187218 370294 187274 370350
rect 187342 370294 187398 370350
rect 186970 370170 187026 370226
rect 187094 370170 187150 370226
rect 187218 370170 187274 370226
rect 187342 370170 187398 370226
rect 186970 370046 187026 370102
rect 187094 370046 187150 370102
rect 187218 370046 187274 370102
rect 187342 370046 187398 370102
rect 186970 369922 187026 369978
rect 187094 369922 187150 369978
rect 187218 369922 187274 369978
rect 187342 369922 187398 369978
rect 186970 352294 187026 352350
rect 187094 352294 187150 352350
rect 187218 352294 187274 352350
rect 187342 352294 187398 352350
rect 186970 352170 187026 352226
rect 187094 352170 187150 352226
rect 187218 352170 187274 352226
rect 187342 352170 187398 352226
rect 186970 352046 187026 352102
rect 187094 352046 187150 352102
rect 187218 352046 187274 352102
rect 187342 352046 187398 352102
rect 186970 351922 187026 351978
rect 187094 351922 187150 351978
rect 187218 351922 187274 351978
rect 187342 351922 187398 351978
rect 186970 334294 187026 334350
rect 187094 334294 187150 334350
rect 187218 334294 187274 334350
rect 187342 334294 187398 334350
rect 186970 334170 187026 334226
rect 187094 334170 187150 334226
rect 187218 334170 187274 334226
rect 187342 334170 187398 334226
rect 186970 334046 187026 334102
rect 187094 334046 187150 334102
rect 187218 334046 187274 334102
rect 187342 334046 187398 334102
rect 186970 333922 187026 333978
rect 187094 333922 187150 333978
rect 187218 333922 187274 333978
rect 187342 333922 187398 333978
rect 186970 316294 187026 316350
rect 187094 316294 187150 316350
rect 187218 316294 187274 316350
rect 187342 316294 187398 316350
rect 186970 316170 187026 316226
rect 187094 316170 187150 316226
rect 187218 316170 187274 316226
rect 187342 316170 187398 316226
rect 186970 316046 187026 316102
rect 187094 316046 187150 316102
rect 187218 316046 187274 316102
rect 187342 316046 187398 316102
rect 186970 315922 187026 315978
rect 187094 315922 187150 315978
rect 187218 315922 187274 315978
rect 187342 315922 187398 315978
rect 186970 298294 187026 298350
rect 187094 298294 187150 298350
rect 187218 298294 187274 298350
rect 187342 298294 187398 298350
rect 186970 298170 187026 298226
rect 187094 298170 187150 298226
rect 187218 298170 187274 298226
rect 187342 298170 187398 298226
rect 186970 298046 187026 298102
rect 187094 298046 187150 298102
rect 187218 298046 187274 298102
rect 187342 298046 187398 298102
rect 186970 297922 187026 297978
rect 187094 297922 187150 297978
rect 187218 297922 187274 297978
rect 187342 297922 187398 297978
rect 186970 280294 187026 280350
rect 187094 280294 187150 280350
rect 187218 280294 187274 280350
rect 187342 280294 187398 280350
rect 186970 280170 187026 280226
rect 187094 280170 187150 280226
rect 187218 280170 187274 280226
rect 187342 280170 187398 280226
rect 186970 280046 187026 280102
rect 187094 280046 187150 280102
rect 187218 280046 187274 280102
rect 187342 280046 187398 280102
rect 186970 279922 187026 279978
rect 187094 279922 187150 279978
rect 187218 279922 187274 279978
rect 187342 279922 187398 279978
rect 186970 262294 187026 262350
rect 187094 262294 187150 262350
rect 187218 262294 187274 262350
rect 187342 262294 187398 262350
rect 186970 262170 187026 262226
rect 187094 262170 187150 262226
rect 187218 262170 187274 262226
rect 187342 262170 187398 262226
rect 186970 262046 187026 262102
rect 187094 262046 187150 262102
rect 187218 262046 187274 262102
rect 187342 262046 187398 262102
rect 186970 261922 187026 261978
rect 187094 261922 187150 261978
rect 187218 261922 187274 261978
rect 187342 261922 187398 261978
rect 186970 244294 187026 244350
rect 187094 244294 187150 244350
rect 187218 244294 187274 244350
rect 187342 244294 187398 244350
rect 186970 244170 187026 244226
rect 187094 244170 187150 244226
rect 187218 244170 187274 244226
rect 187342 244170 187398 244226
rect 186970 244046 187026 244102
rect 187094 244046 187150 244102
rect 187218 244046 187274 244102
rect 187342 244046 187398 244102
rect 186970 243922 187026 243978
rect 187094 243922 187150 243978
rect 187218 243922 187274 243978
rect 187342 243922 187398 243978
rect 186970 226294 187026 226350
rect 187094 226294 187150 226350
rect 187218 226294 187274 226350
rect 187342 226294 187398 226350
rect 186970 226170 187026 226226
rect 187094 226170 187150 226226
rect 187218 226170 187274 226226
rect 187342 226170 187398 226226
rect 186970 226046 187026 226102
rect 187094 226046 187150 226102
rect 187218 226046 187274 226102
rect 187342 226046 187398 226102
rect 186970 225922 187026 225978
rect 187094 225922 187150 225978
rect 187218 225922 187274 225978
rect 187342 225922 187398 225978
rect 186970 208294 187026 208350
rect 187094 208294 187150 208350
rect 187218 208294 187274 208350
rect 187342 208294 187398 208350
rect 186970 208170 187026 208226
rect 187094 208170 187150 208226
rect 187218 208170 187274 208226
rect 187342 208170 187398 208226
rect 186970 208046 187026 208102
rect 187094 208046 187150 208102
rect 187218 208046 187274 208102
rect 187342 208046 187398 208102
rect 186970 207922 187026 207978
rect 187094 207922 187150 207978
rect 187218 207922 187274 207978
rect 187342 207922 187398 207978
rect 186970 190294 187026 190350
rect 187094 190294 187150 190350
rect 187218 190294 187274 190350
rect 187342 190294 187398 190350
rect 186970 190170 187026 190226
rect 187094 190170 187150 190226
rect 187218 190170 187274 190226
rect 187342 190170 187398 190226
rect 186970 190046 187026 190102
rect 187094 190046 187150 190102
rect 187218 190046 187274 190102
rect 187342 190046 187398 190102
rect 186970 189922 187026 189978
rect 187094 189922 187150 189978
rect 187218 189922 187274 189978
rect 187342 189922 187398 189978
rect 186970 172294 187026 172350
rect 187094 172294 187150 172350
rect 187218 172294 187274 172350
rect 187342 172294 187398 172350
rect 186970 172170 187026 172226
rect 187094 172170 187150 172226
rect 187218 172170 187274 172226
rect 187342 172170 187398 172226
rect 186970 172046 187026 172102
rect 187094 172046 187150 172102
rect 187218 172046 187274 172102
rect 187342 172046 187398 172102
rect 186970 171922 187026 171978
rect 187094 171922 187150 171978
rect 187218 171922 187274 171978
rect 187342 171922 187398 171978
rect 186970 154294 187026 154350
rect 187094 154294 187150 154350
rect 187218 154294 187274 154350
rect 187342 154294 187398 154350
rect 186970 154170 187026 154226
rect 187094 154170 187150 154226
rect 187218 154170 187274 154226
rect 187342 154170 187398 154226
rect 186970 154046 187026 154102
rect 187094 154046 187150 154102
rect 187218 154046 187274 154102
rect 187342 154046 187398 154102
rect 186970 153922 187026 153978
rect 187094 153922 187150 153978
rect 187218 153922 187274 153978
rect 187342 153922 187398 153978
rect 186970 136294 187026 136350
rect 187094 136294 187150 136350
rect 187218 136294 187274 136350
rect 187342 136294 187398 136350
rect 186970 136170 187026 136226
rect 187094 136170 187150 136226
rect 187218 136170 187274 136226
rect 187342 136170 187398 136226
rect 186970 136046 187026 136102
rect 187094 136046 187150 136102
rect 187218 136046 187274 136102
rect 187342 136046 187398 136102
rect 186970 135922 187026 135978
rect 187094 135922 187150 135978
rect 187218 135922 187274 135978
rect 187342 135922 187398 135978
rect 186970 118294 187026 118350
rect 187094 118294 187150 118350
rect 187218 118294 187274 118350
rect 187342 118294 187398 118350
rect 186970 118170 187026 118226
rect 187094 118170 187150 118226
rect 187218 118170 187274 118226
rect 187342 118170 187398 118226
rect 186970 118046 187026 118102
rect 187094 118046 187150 118102
rect 187218 118046 187274 118102
rect 187342 118046 187398 118102
rect 186970 117922 187026 117978
rect 187094 117922 187150 117978
rect 187218 117922 187274 117978
rect 187342 117922 187398 117978
rect 186970 100294 187026 100350
rect 187094 100294 187150 100350
rect 187218 100294 187274 100350
rect 187342 100294 187398 100350
rect 186970 100170 187026 100226
rect 187094 100170 187150 100226
rect 187218 100170 187274 100226
rect 187342 100170 187398 100226
rect 186970 100046 187026 100102
rect 187094 100046 187150 100102
rect 187218 100046 187274 100102
rect 187342 100046 187398 100102
rect 186970 99922 187026 99978
rect 187094 99922 187150 99978
rect 187218 99922 187274 99978
rect 187342 99922 187398 99978
rect 186970 82294 187026 82350
rect 187094 82294 187150 82350
rect 187218 82294 187274 82350
rect 187342 82294 187398 82350
rect 186970 82170 187026 82226
rect 187094 82170 187150 82226
rect 187218 82170 187274 82226
rect 187342 82170 187398 82226
rect 186970 82046 187026 82102
rect 187094 82046 187150 82102
rect 187218 82046 187274 82102
rect 187342 82046 187398 82102
rect 186970 81922 187026 81978
rect 187094 81922 187150 81978
rect 187218 81922 187274 81978
rect 187342 81922 187398 81978
rect 186970 64294 187026 64350
rect 187094 64294 187150 64350
rect 187218 64294 187274 64350
rect 187342 64294 187398 64350
rect 186970 64170 187026 64226
rect 187094 64170 187150 64226
rect 187218 64170 187274 64226
rect 187342 64170 187398 64226
rect 186970 64046 187026 64102
rect 187094 64046 187150 64102
rect 187218 64046 187274 64102
rect 187342 64046 187398 64102
rect 186970 63922 187026 63978
rect 187094 63922 187150 63978
rect 187218 63922 187274 63978
rect 187342 63922 187398 63978
rect 186970 46294 187026 46350
rect 187094 46294 187150 46350
rect 187218 46294 187274 46350
rect 187342 46294 187398 46350
rect 186970 46170 187026 46226
rect 187094 46170 187150 46226
rect 187218 46170 187274 46226
rect 187342 46170 187398 46226
rect 186970 46046 187026 46102
rect 187094 46046 187150 46102
rect 187218 46046 187274 46102
rect 187342 46046 187398 46102
rect 186970 45922 187026 45978
rect 187094 45922 187150 45978
rect 187218 45922 187274 45978
rect 187342 45922 187398 45978
rect 186970 28294 187026 28350
rect 187094 28294 187150 28350
rect 187218 28294 187274 28350
rect 187342 28294 187398 28350
rect 186970 28170 187026 28226
rect 187094 28170 187150 28226
rect 187218 28170 187274 28226
rect 187342 28170 187398 28226
rect 186970 28046 187026 28102
rect 187094 28046 187150 28102
rect 187218 28046 187274 28102
rect 187342 28046 187398 28102
rect 186970 27922 187026 27978
rect 187094 27922 187150 27978
rect 187218 27922 187274 27978
rect 187342 27922 187398 27978
rect 186970 10294 187026 10350
rect 187094 10294 187150 10350
rect 187218 10294 187274 10350
rect 187342 10294 187398 10350
rect 186970 10170 187026 10226
rect 187094 10170 187150 10226
rect 187218 10170 187274 10226
rect 187342 10170 187398 10226
rect 186970 10046 187026 10102
rect 187094 10046 187150 10102
rect 187218 10046 187274 10102
rect 187342 10046 187398 10102
rect 186970 9922 187026 9978
rect 187094 9922 187150 9978
rect 187218 9922 187274 9978
rect 187342 9922 187398 9978
rect 186970 -1176 187026 -1120
rect 187094 -1176 187150 -1120
rect 187218 -1176 187274 -1120
rect 187342 -1176 187398 -1120
rect 186970 -1300 187026 -1244
rect 187094 -1300 187150 -1244
rect 187218 -1300 187274 -1244
rect 187342 -1300 187398 -1244
rect 186970 -1424 187026 -1368
rect 187094 -1424 187150 -1368
rect 187218 -1424 187274 -1368
rect 187342 -1424 187398 -1368
rect 186970 -1548 187026 -1492
rect 187094 -1548 187150 -1492
rect 187218 -1548 187274 -1492
rect 187342 -1548 187398 -1492
rect 201250 597156 201306 597212
rect 201374 597156 201430 597212
rect 201498 597156 201554 597212
rect 201622 597156 201678 597212
rect 201250 597032 201306 597088
rect 201374 597032 201430 597088
rect 201498 597032 201554 597088
rect 201622 597032 201678 597088
rect 201250 596908 201306 596964
rect 201374 596908 201430 596964
rect 201498 596908 201554 596964
rect 201622 596908 201678 596964
rect 201250 596784 201306 596840
rect 201374 596784 201430 596840
rect 201498 596784 201554 596840
rect 201622 596784 201678 596840
rect 201250 580294 201306 580350
rect 201374 580294 201430 580350
rect 201498 580294 201554 580350
rect 201622 580294 201678 580350
rect 201250 580170 201306 580226
rect 201374 580170 201430 580226
rect 201498 580170 201554 580226
rect 201622 580170 201678 580226
rect 201250 580046 201306 580102
rect 201374 580046 201430 580102
rect 201498 580046 201554 580102
rect 201622 580046 201678 580102
rect 201250 579922 201306 579978
rect 201374 579922 201430 579978
rect 201498 579922 201554 579978
rect 201622 579922 201678 579978
rect 201250 562294 201306 562350
rect 201374 562294 201430 562350
rect 201498 562294 201554 562350
rect 201622 562294 201678 562350
rect 201250 562170 201306 562226
rect 201374 562170 201430 562226
rect 201498 562170 201554 562226
rect 201622 562170 201678 562226
rect 201250 562046 201306 562102
rect 201374 562046 201430 562102
rect 201498 562046 201554 562102
rect 201622 562046 201678 562102
rect 201250 561922 201306 561978
rect 201374 561922 201430 561978
rect 201498 561922 201554 561978
rect 201622 561922 201678 561978
rect 201250 544294 201306 544350
rect 201374 544294 201430 544350
rect 201498 544294 201554 544350
rect 201622 544294 201678 544350
rect 201250 544170 201306 544226
rect 201374 544170 201430 544226
rect 201498 544170 201554 544226
rect 201622 544170 201678 544226
rect 201250 544046 201306 544102
rect 201374 544046 201430 544102
rect 201498 544046 201554 544102
rect 201622 544046 201678 544102
rect 201250 543922 201306 543978
rect 201374 543922 201430 543978
rect 201498 543922 201554 543978
rect 201622 543922 201678 543978
rect 201250 526294 201306 526350
rect 201374 526294 201430 526350
rect 201498 526294 201554 526350
rect 201622 526294 201678 526350
rect 201250 526170 201306 526226
rect 201374 526170 201430 526226
rect 201498 526170 201554 526226
rect 201622 526170 201678 526226
rect 201250 526046 201306 526102
rect 201374 526046 201430 526102
rect 201498 526046 201554 526102
rect 201622 526046 201678 526102
rect 201250 525922 201306 525978
rect 201374 525922 201430 525978
rect 201498 525922 201554 525978
rect 201622 525922 201678 525978
rect 201250 508294 201306 508350
rect 201374 508294 201430 508350
rect 201498 508294 201554 508350
rect 201622 508294 201678 508350
rect 201250 508170 201306 508226
rect 201374 508170 201430 508226
rect 201498 508170 201554 508226
rect 201622 508170 201678 508226
rect 201250 508046 201306 508102
rect 201374 508046 201430 508102
rect 201498 508046 201554 508102
rect 201622 508046 201678 508102
rect 201250 507922 201306 507978
rect 201374 507922 201430 507978
rect 201498 507922 201554 507978
rect 201622 507922 201678 507978
rect 204970 598116 205026 598172
rect 205094 598116 205150 598172
rect 205218 598116 205274 598172
rect 205342 598116 205398 598172
rect 204970 597992 205026 598048
rect 205094 597992 205150 598048
rect 205218 597992 205274 598048
rect 205342 597992 205398 598048
rect 204970 597868 205026 597924
rect 205094 597868 205150 597924
rect 205218 597868 205274 597924
rect 205342 597868 205398 597924
rect 204970 597744 205026 597800
rect 205094 597744 205150 597800
rect 205218 597744 205274 597800
rect 205342 597744 205398 597800
rect 204970 586294 205026 586350
rect 205094 586294 205150 586350
rect 205218 586294 205274 586350
rect 205342 586294 205398 586350
rect 204970 586170 205026 586226
rect 205094 586170 205150 586226
rect 205218 586170 205274 586226
rect 205342 586170 205398 586226
rect 204970 586046 205026 586102
rect 205094 586046 205150 586102
rect 205218 586046 205274 586102
rect 205342 586046 205398 586102
rect 204970 585922 205026 585978
rect 205094 585922 205150 585978
rect 205218 585922 205274 585978
rect 205342 585922 205398 585978
rect 204970 568294 205026 568350
rect 205094 568294 205150 568350
rect 205218 568294 205274 568350
rect 205342 568294 205398 568350
rect 204970 568170 205026 568226
rect 205094 568170 205150 568226
rect 205218 568170 205274 568226
rect 205342 568170 205398 568226
rect 204970 568046 205026 568102
rect 205094 568046 205150 568102
rect 205218 568046 205274 568102
rect 205342 568046 205398 568102
rect 204970 567922 205026 567978
rect 205094 567922 205150 567978
rect 205218 567922 205274 567978
rect 205342 567922 205398 567978
rect 204970 550294 205026 550350
rect 205094 550294 205150 550350
rect 205218 550294 205274 550350
rect 205342 550294 205398 550350
rect 204970 550170 205026 550226
rect 205094 550170 205150 550226
rect 205218 550170 205274 550226
rect 205342 550170 205398 550226
rect 204970 550046 205026 550102
rect 205094 550046 205150 550102
rect 205218 550046 205274 550102
rect 205342 550046 205398 550102
rect 204970 549922 205026 549978
rect 205094 549922 205150 549978
rect 205218 549922 205274 549978
rect 205342 549922 205398 549978
rect 204970 532294 205026 532350
rect 205094 532294 205150 532350
rect 205218 532294 205274 532350
rect 205342 532294 205398 532350
rect 204970 532170 205026 532226
rect 205094 532170 205150 532226
rect 205218 532170 205274 532226
rect 205342 532170 205398 532226
rect 204970 532046 205026 532102
rect 205094 532046 205150 532102
rect 205218 532046 205274 532102
rect 205342 532046 205398 532102
rect 204970 531922 205026 531978
rect 205094 531922 205150 531978
rect 205218 531922 205274 531978
rect 205342 531922 205398 531978
rect 204970 514294 205026 514350
rect 205094 514294 205150 514350
rect 205218 514294 205274 514350
rect 205342 514294 205398 514350
rect 204970 514170 205026 514226
rect 205094 514170 205150 514226
rect 205218 514170 205274 514226
rect 205342 514170 205398 514226
rect 204970 514046 205026 514102
rect 205094 514046 205150 514102
rect 205218 514046 205274 514102
rect 205342 514046 205398 514102
rect 204970 513922 205026 513978
rect 205094 513922 205150 513978
rect 205218 513922 205274 513978
rect 205342 513922 205398 513978
rect 219250 597156 219306 597212
rect 219374 597156 219430 597212
rect 219498 597156 219554 597212
rect 219622 597156 219678 597212
rect 219250 597032 219306 597088
rect 219374 597032 219430 597088
rect 219498 597032 219554 597088
rect 219622 597032 219678 597088
rect 219250 596908 219306 596964
rect 219374 596908 219430 596964
rect 219498 596908 219554 596964
rect 219622 596908 219678 596964
rect 219250 596784 219306 596840
rect 219374 596784 219430 596840
rect 219498 596784 219554 596840
rect 219622 596784 219678 596840
rect 219250 580294 219306 580350
rect 219374 580294 219430 580350
rect 219498 580294 219554 580350
rect 219622 580294 219678 580350
rect 219250 580170 219306 580226
rect 219374 580170 219430 580226
rect 219498 580170 219554 580226
rect 219622 580170 219678 580226
rect 219250 580046 219306 580102
rect 219374 580046 219430 580102
rect 219498 580046 219554 580102
rect 219622 580046 219678 580102
rect 219250 579922 219306 579978
rect 219374 579922 219430 579978
rect 219498 579922 219554 579978
rect 219622 579922 219678 579978
rect 219250 562294 219306 562350
rect 219374 562294 219430 562350
rect 219498 562294 219554 562350
rect 219622 562294 219678 562350
rect 219250 562170 219306 562226
rect 219374 562170 219430 562226
rect 219498 562170 219554 562226
rect 219622 562170 219678 562226
rect 219250 562046 219306 562102
rect 219374 562046 219430 562102
rect 219498 562046 219554 562102
rect 219622 562046 219678 562102
rect 219250 561922 219306 561978
rect 219374 561922 219430 561978
rect 219498 561922 219554 561978
rect 219622 561922 219678 561978
rect 219250 544294 219306 544350
rect 219374 544294 219430 544350
rect 219498 544294 219554 544350
rect 219622 544294 219678 544350
rect 219250 544170 219306 544226
rect 219374 544170 219430 544226
rect 219498 544170 219554 544226
rect 219622 544170 219678 544226
rect 219250 544046 219306 544102
rect 219374 544046 219430 544102
rect 219498 544046 219554 544102
rect 219622 544046 219678 544102
rect 219250 543922 219306 543978
rect 219374 543922 219430 543978
rect 219498 543922 219554 543978
rect 219622 543922 219678 543978
rect 219250 526294 219306 526350
rect 219374 526294 219430 526350
rect 219498 526294 219554 526350
rect 219622 526294 219678 526350
rect 219250 526170 219306 526226
rect 219374 526170 219430 526226
rect 219498 526170 219554 526226
rect 219622 526170 219678 526226
rect 219250 526046 219306 526102
rect 219374 526046 219430 526102
rect 219498 526046 219554 526102
rect 219622 526046 219678 526102
rect 219250 525922 219306 525978
rect 219374 525922 219430 525978
rect 219498 525922 219554 525978
rect 219622 525922 219678 525978
rect 219250 508294 219306 508350
rect 219374 508294 219430 508350
rect 219498 508294 219554 508350
rect 219622 508294 219678 508350
rect 219250 508170 219306 508226
rect 219374 508170 219430 508226
rect 219498 508170 219554 508226
rect 219622 508170 219678 508226
rect 219250 508046 219306 508102
rect 219374 508046 219430 508102
rect 219498 508046 219554 508102
rect 219622 508046 219678 508102
rect 219250 507922 219306 507978
rect 219374 507922 219430 507978
rect 219498 507922 219554 507978
rect 219622 507922 219678 507978
rect 222970 598116 223026 598172
rect 223094 598116 223150 598172
rect 223218 598116 223274 598172
rect 223342 598116 223398 598172
rect 222970 597992 223026 598048
rect 223094 597992 223150 598048
rect 223218 597992 223274 598048
rect 223342 597992 223398 598048
rect 222970 597868 223026 597924
rect 223094 597868 223150 597924
rect 223218 597868 223274 597924
rect 223342 597868 223398 597924
rect 222970 597744 223026 597800
rect 223094 597744 223150 597800
rect 223218 597744 223274 597800
rect 223342 597744 223398 597800
rect 222970 586294 223026 586350
rect 223094 586294 223150 586350
rect 223218 586294 223274 586350
rect 223342 586294 223398 586350
rect 222970 586170 223026 586226
rect 223094 586170 223150 586226
rect 223218 586170 223274 586226
rect 223342 586170 223398 586226
rect 222970 586046 223026 586102
rect 223094 586046 223150 586102
rect 223218 586046 223274 586102
rect 223342 586046 223398 586102
rect 222970 585922 223026 585978
rect 223094 585922 223150 585978
rect 223218 585922 223274 585978
rect 223342 585922 223398 585978
rect 222970 568294 223026 568350
rect 223094 568294 223150 568350
rect 223218 568294 223274 568350
rect 223342 568294 223398 568350
rect 222970 568170 223026 568226
rect 223094 568170 223150 568226
rect 223218 568170 223274 568226
rect 223342 568170 223398 568226
rect 222970 568046 223026 568102
rect 223094 568046 223150 568102
rect 223218 568046 223274 568102
rect 223342 568046 223398 568102
rect 222970 567922 223026 567978
rect 223094 567922 223150 567978
rect 223218 567922 223274 567978
rect 223342 567922 223398 567978
rect 222970 550294 223026 550350
rect 223094 550294 223150 550350
rect 223218 550294 223274 550350
rect 223342 550294 223398 550350
rect 222970 550170 223026 550226
rect 223094 550170 223150 550226
rect 223218 550170 223274 550226
rect 223342 550170 223398 550226
rect 222970 550046 223026 550102
rect 223094 550046 223150 550102
rect 223218 550046 223274 550102
rect 223342 550046 223398 550102
rect 222970 549922 223026 549978
rect 223094 549922 223150 549978
rect 223218 549922 223274 549978
rect 223342 549922 223398 549978
rect 222970 532294 223026 532350
rect 223094 532294 223150 532350
rect 223218 532294 223274 532350
rect 223342 532294 223398 532350
rect 222970 532170 223026 532226
rect 223094 532170 223150 532226
rect 223218 532170 223274 532226
rect 223342 532170 223398 532226
rect 222970 532046 223026 532102
rect 223094 532046 223150 532102
rect 223218 532046 223274 532102
rect 223342 532046 223398 532102
rect 222970 531922 223026 531978
rect 223094 531922 223150 531978
rect 223218 531922 223274 531978
rect 223342 531922 223398 531978
rect 222970 514294 223026 514350
rect 223094 514294 223150 514350
rect 223218 514294 223274 514350
rect 223342 514294 223398 514350
rect 222970 514170 223026 514226
rect 223094 514170 223150 514226
rect 223218 514170 223274 514226
rect 223342 514170 223398 514226
rect 222970 514046 223026 514102
rect 223094 514046 223150 514102
rect 223218 514046 223274 514102
rect 223342 514046 223398 514102
rect 222970 513922 223026 513978
rect 223094 513922 223150 513978
rect 223218 513922 223274 513978
rect 223342 513922 223398 513978
rect 237250 597156 237306 597212
rect 237374 597156 237430 597212
rect 237498 597156 237554 597212
rect 237622 597156 237678 597212
rect 237250 597032 237306 597088
rect 237374 597032 237430 597088
rect 237498 597032 237554 597088
rect 237622 597032 237678 597088
rect 237250 596908 237306 596964
rect 237374 596908 237430 596964
rect 237498 596908 237554 596964
rect 237622 596908 237678 596964
rect 237250 596784 237306 596840
rect 237374 596784 237430 596840
rect 237498 596784 237554 596840
rect 237622 596784 237678 596840
rect 237250 580294 237306 580350
rect 237374 580294 237430 580350
rect 237498 580294 237554 580350
rect 237622 580294 237678 580350
rect 237250 580170 237306 580226
rect 237374 580170 237430 580226
rect 237498 580170 237554 580226
rect 237622 580170 237678 580226
rect 237250 580046 237306 580102
rect 237374 580046 237430 580102
rect 237498 580046 237554 580102
rect 237622 580046 237678 580102
rect 237250 579922 237306 579978
rect 237374 579922 237430 579978
rect 237498 579922 237554 579978
rect 237622 579922 237678 579978
rect 237250 562294 237306 562350
rect 237374 562294 237430 562350
rect 237498 562294 237554 562350
rect 237622 562294 237678 562350
rect 237250 562170 237306 562226
rect 237374 562170 237430 562226
rect 237498 562170 237554 562226
rect 237622 562170 237678 562226
rect 237250 562046 237306 562102
rect 237374 562046 237430 562102
rect 237498 562046 237554 562102
rect 237622 562046 237678 562102
rect 237250 561922 237306 561978
rect 237374 561922 237430 561978
rect 237498 561922 237554 561978
rect 237622 561922 237678 561978
rect 237250 544294 237306 544350
rect 237374 544294 237430 544350
rect 237498 544294 237554 544350
rect 237622 544294 237678 544350
rect 237250 544170 237306 544226
rect 237374 544170 237430 544226
rect 237498 544170 237554 544226
rect 237622 544170 237678 544226
rect 237250 544046 237306 544102
rect 237374 544046 237430 544102
rect 237498 544046 237554 544102
rect 237622 544046 237678 544102
rect 237250 543922 237306 543978
rect 237374 543922 237430 543978
rect 237498 543922 237554 543978
rect 237622 543922 237678 543978
rect 237250 526294 237306 526350
rect 237374 526294 237430 526350
rect 237498 526294 237554 526350
rect 237622 526294 237678 526350
rect 237250 526170 237306 526226
rect 237374 526170 237430 526226
rect 237498 526170 237554 526226
rect 237622 526170 237678 526226
rect 237250 526046 237306 526102
rect 237374 526046 237430 526102
rect 237498 526046 237554 526102
rect 237622 526046 237678 526102
rect 237250 525922 237306 525978
rect 237374 525922 237430 525978
rect 237498 525922 237554 525978
rect 237622 525922 237678 525978
rect 237250 508294 237306 508350
rect 237374 508294 237430 508350
rect 237498 508294 237554 508350
rect 237622 508294 237678 508350
rect 237250 508170 237306 508226
rect 237374 508170 237430 508226
rect 237498 508170 237554 508226
rect 237622 508170 237678 508226
rect 237250 508046 237306 508102
rect 237374 508046 237430 508102
rect 237498 508046 237554 508102
rect 237622 508046 237678 508102
rect 237250 507922 237306 507978
rect 237374 507922 237430 507978
rect 237498 507922 237554 507978
rect 237622 507922 237678 507978
rect 240970 598116 241026 598172
rect 241094 598116 241150 598172
rect 241218 598116 241274 598172
rect 241342 598116 241398 598172
rect 240970 597992 241026 598048
rect 241094 597992 241150 598048
rect 241218 597992 241274 598048
rect 241342 597992 241398 598048
rect 240970 597868 241026 597924
rect 241094 597868 241150 597924
rect 241218 597868 241274 597924
rect 241342 597868 241398 597924
rect 240970 597744 241026 597800
rect 241094 597744 241150 597800
rect 241218 597744 241274 597800
rect 241342 597744 241398 597800
rect 240970 586294 241026 586350
rect 241094 586294 241150 586350
rect 241218 586294 241274 586350
rect 241342 586294 241398 586350
rect 240970 586170 241026 586226
rect 241094 586170 241150 586226
rect 241218 586170 241274 586226
rect 241342 586170 241398 586226
rect 240970 586046 241026 586102
rect 241094 586046 241150 586102
rect 241218 586046 241274 586102
rect 241342 586046 241398 586102
rect 240970 585922 241026 585978
rect 241094 585922 241150 585978
rect 241218 585922 241274 585978
rect 241342 585922 241398 585978
rect 240970 568294 241026 568350
rect 241094 568294 241150 568350
rect 241218 568294 241274 568350
rect 241342 568294 241398 568350
rect 240970 568170 241026 568226
rect 241094 568170 241150 568226
rect 241218 568170 241274 568226
rect 241342 568170 241398 568226
rect 240970 568046 241026 568102
rect 241094 568046 241150 568102
rect 241218 568046 241274 568102
rect 241342 568046 241398 568102
rect 240970 567922 241026 567978
rect 241094 567922 241150 567978
rect 241218 567922 241274 567978
rect 241342 567922 241398 567978
rect 240970 550294 241026 550350
rect 241094 550294 241150 550350
rect 241218 550294 241274 550350
rect 241342 550294 241398 550350
rect 240970 550170 241026 550226
rect 241094 550170 241150 550226
rect 241218 550170 241274 550226
rect 241342 550170 241398 550226
rect 240970 550046 241026 550102
rect 241094 550046 241150 550102
rect 241218 550046 241274 550102
rect 241342 550046 241398 550102
rect 240970 549922 241026 549978
rect 241094 549922 241150 549978
rect 241218 549922 241274 549978
rect 241342 549922 241398 549978
rect 240970 532294 241026 532350
rect 241094 532294 241150 532350
rect 241218 532294 241274 532350
rect 241342 532294 241398 532350
rect 240970 532170 241026 532226
rect 241094 532170 241150 532226
rect 241218 532170 241274 532226
rect 241342 532170 241398 532226
rect 240970 532046 241026 532102
rect 241094 532046 241150 532102
rect 241218 532046 241274 532102
rect 241342 532046 241398 532102
rect 240970 531922 241026 531978
rect 241094 531922 241150 531978
rect 241218 531922 241274 531978
rect 241342 531922 241398 531978
rect 240970 514294 241026 514350
rect 241094 514294 241150 514350
rect 241218 514294 241274 514350
rect 241342 514294 241398 514350
rect 240970 514170 241026 514226
rect 241094 514170 241150 514226
rect 241218 514170 241274 514226
rect 241342 514170 241398 514226
rect 240970 514046 241026 514102
rect 241094 514046 241150 514102
rect 241218 514046 241274 514102
rect 241342 514046 241398 514102
rect 240970 513922 241026 513978
rect 241094 513922 241150 513978
rect 241218 513922 241274 513978
rect 241342 513922 241398 513978
rect 255250 597156 255306 597212
rect 255374 597156 255430 597212
rect 255498 597156 255554 597212
rect 255622 597156 255678 597212
rect 255250 597032 255306 597088
rect 255374 597032 255430 597088
rect 255498 597032 255554 597088
rect 255622 597032 255678 597088
rect 255250 596908 255306 596964
rect 255374 596908 255430 596964
rect 255498 596908 255554 596964
rect 255622 596908 255678 596964
rect 255250 596784 255306 596840
rect 255374 596784 255430 596840
rect 255498 596784 255554 596840
rect 255622 596784 255678 596840
rect 255250 580294 255306 580350
rect 255374 580294 255430 580350
rect 255498 580294 255554 580350
rect 255622 580294 255678 580350
rect 255250 580170 255306 580226
rect 255374 580170 255430 580226
rect 255498 580170 255554 580226
rect 255622 580170 255678 580226
rect 255250 580046 255306 580102
rect 255374 580046 255430 580102
rect 255498 580046 255554 580102
rect 255622 580046 255678 580102
rect 255250 579922 255306 579978
rect 255374 579922 255430 579978
rect 255498 579922 255554 579978
rect 255622 579922 255678 579978
rect 255250 562294 255306 562350
rect 255374 562294 255430 562350
rect 255498 562294 255554 562350
rect 255622 562294 255678 562350
rect 255250 562170 255306 562226
rect 255374 562170 255430 562226
rect 255498 562170 255554 562226
rect 255622 562170 255678 562226
rect 255250 562046 255306 562102
rect 255374 562046 255430 562102
rect 255498 562046 255554 562102
rect 255622 562046 255678 562102
rect 255250 561922 255306 561978
rect 255374 561922 255430 561978
rect 255498 561922 255554 561978
rect 255622 561922 255678 561978
rect 255250 544294 255306 544350
rect 255374 544294 255430 544350
rect 255498 544294 255554 544350
rect 255622 544294 255678 544350
rect 255250 544170 255306 544226
rect 255374 544170 255430 544226
rect 255498 544170 255554 544226
rect 255622 544170 255678 544226
rect 255250 544046 255306 544102
rect 255374 544046 255430 544102
rect 255498 544046 255554 544102
rect 255622 544046 255678 544102
rect 255250 543922 255306 543978
rect 255374 543922 255430 543978
rect 255498 543922 255554 543978
rect 255622 543922 255678 543978
rect 255250 526294 255306 526350
rect 255374 526294 255430 526350
rect 255498 526294 255554 526350
rect 255622 526294 255678 526350
rect 255250 526170 255306 526226
rect 255374 526170 255430 526226
rect 255498 526170 255554 526226
rect 255622 526170 255678 526226
rect 255250 526046 255306 526102
rect 255374 526046 255430 526102
rect 255498 526046 255554 526102
rect 255622 526046 255678 526102
rect 255250 525922 255306 525978
rect 255374 525922 255430 525978
rect 255498 525922 255554 525978
rect 255622 525922 255678 525978
rect 255250 508294 255306 508350
rect 255374 508294 255430 508350
rect 255498 508294 255554 508350
rect 255622 508294 255678 508350
rect 255250 508170 255306 508226
rect 255374 508170 255430 508226
rect 255498 508170 255554 508226
rect 255622 508170 255678 508226
rect 255250 508046 255306 508102
rect 255374 508046 255430 508102
rect 255498 508046 255554 508102
rect 255622 508046 255678 508102
rect 255250 507922 255306 507978
rect 255374 507922 255430 507978
rect 255498 507922 255554 507978
rect 255622 507922 255678 507978
rect 258970 598116 259026 598172
rect 259094 598116 259150 598172
rect 259218 598116 259274 598172
rect 259342 598116 259398 598172
rect 258970 597992 259026 598048
rect 259094 597992 259150 598048
rect 259218 597992 259274 598048
rect 259342 597992 259398 598048
rect 258970 597868 259026 597924
rect 259094 597868 259150 597924
rect 259218 597868 259274 597924
rect 259342 597868 259398 597924
rect 258970 597744 259026 597800
rect 259094 597744 259150 597800
rect 259218 597744 259274 597800
rect 259342 597744 259398 597800
rect 258970 586294 259026 586350
rect 259094 586294 259150 586350
rect 259218 586294 259274 586350
rect 259342 586294 259398 586350
rect 258970 586170 259026 586226
rect 259094 586170 259150 586226
rect 259218 586170 259274 586226
rect 259342 586170 259398 586226
rect 258970 586046 259026 586102
rect 259094 586046 259150 586102
rect 259218 586046 259274 586102
rect 259342 586046 259398 586102
rect 258970 585922 259026 585978
rect 259094 585922 259150 585978
rect 259218 585922 259274 585978
rect 259342 585922 259398 585978
rect 258970 568294 259026 568350
rect 259094 568294 259150 568350
rect 259218 568294 259274 568350
rect 259342 568294 259398 568350
rect 258970 568170 259026 568226
rect 259094 568170 259150 568226
rect 259218 568170 259274 568226
rect 259342 568170 259398 568226
rect 258970 568046 259026 568102
rect 259094 568046 259150 568102
rect 259218 568046 259274 568102
rect 259342 568046 259398 568102
rect 258970 567922 259026 567978
rect 259094 567922 259150 567978
rect 259218 567922 259274 567978
rect 259342 567922 259398 567978
rect 258970 550294 259026 550350
rect 259094 550294 259150 550350
rect 259218 550294 259274 550350
rect 259342 550294 259398 550350
rect 258970 550170 259026 550226
rect 259094 550170 259150 550226
rect 259218 550170 259274 550226
rect 259342 550170 259398 550226
rect 258970 550046 259026 550102
rect 259094 550046 259150 550102
rect 259218 550046 259274 550102
rect 259342 550046 259398 550102
rect 258970 549922 259026 549978
rect 259094 549922 259150 549978
rect 259218 549922 259274 549978
rect 259342 549922 259398 549978
rect 258970 532294 259026 532350
rect 259094 532294 259150 532350
rect 259218 532294 259274 532350
rect 259342 532294 259398 532350
rect 258970 532170 259026 532226
rect 259094 532170 259150 532226
rect 259218 532170 259274 532226
rect 259342 532170 259398 532226
rect 258970 532046 259026 532102
rect 259094 532046 259150 532102
rect 259218 532046 259274 532102
rect 259342 532046 259398 532102
rect 258970 531922 259026 531978
rect 259094 531922 259150 531978
rect 259218 531922 259274 531978
rect 259342 531922 259398 531978
rect 258970 514294 259026 514350
rect 259094 514294 259150 514350
rect 259218 514294 259274 514350
rect 259342 514294 259398 514350
rect 258970 514170 259026 514226
rect 259094 514170 259150 514226
rect 259218 514170 259274 514226
rect 259342 514170 259398 514226
rect 258970 514046 259026 514102
rect 259094 514046 259150 514102
rect 259218 514046 259274 514102
rect 259342 514046 259398 514102
rect 258970 513922 259026 513978
rect 259094 513922 259150 513978
rect 259218 513922 259274 513978
rect 259342 513922 259398 513978
rect 273250 597156 273306 597212
rect 273374 597156 273430 597212
rect 273498 597156 273554 597212
rect 273622 597156 273678 597212
rect 273250 597032 273306 597088
rect 273374 597032 273430 597088
rect 273498 597032 273554 597088
rect 273622 597032 273678 597088
rect 273250 596908 273306 596964
rect 273374 596908 273430 596964
rect 273498 596908 273554 596964
rect 273622 596908 273678 596964
rect 273250 596784 273306 596840
rect 273374 596784 273430 596840
rect 273498 596784 273554 596840
rect 273622 596784 273678 596840
rect 273250 580294 273306 580350
rect 273374 580294 273430 580350
rect 273498 580294 273554 580350
rect 273622 580294 273678 580350
rect 273250 580170 273306 580226
rect 273374 580170 273430 580226
rect 273498 580170 273554 580226
rect 273622 580170 273678 580226
rect 273250 580046 273306 580102
rect 273374 580046 273430 580102
rect 273498 580046 273554 580102
rect 273622 580046 273678 580102
rect 273250 579922 273306 579978
rect 273374 579922 273430 579978
rect 273498 579922 273554 579978
rect 273622 579922 273678 579978
rect 273250 562294 273306 562350
rect 273374 562294 273430 562350
rect 273498 562294 273554 562350
rect 273622 562294 273678 562350
rect 273250 562170 273306 562226
rect 273374 562170 273430 562226
rect 273498 562170 273554 562226
rect 273622 562170 273678 562226
rect 273250 562046 273306 562102
rect 273374 562046 273430 562102
rect 273498 562046 273554 562102
rect 273622 562046 273678 562102
rect 273250 561922 273306 561978
rect 273374 561922 273430 561978
rect 273498 561922 273554 561978
rect 273622 561922 273678 561978
rect 273250 544294 273306 544350
rect 273374 544294 273430 544350
rect 273498 544294 273554 544350
rect 273622 544294 273678 544350
rect 273250 544170 273306 544226
rect 273374 544170 273430 544226
rect 273498 544170 273554 544226
rect 273622 544170 273678 544226
rect 273250 544046 273306 544102
rect 273374 544046 273430 544102
rect 273498 544046 273554 544102
rect 273622 544046 273678 544102
rect 273250 543922 273306 543978
rect 273374 543922 273430 543978
rect 273498 543922 273554 543978
rect 273622 543922 273678 543978
rect 273250 526294 273306 526350
rect 273374 526294 273430 526350
rect 273498 526294 273554 526350
rect 273622 526294 273678 526350
rect 273250 526170 273306 526226
rect 273374 526170 273430 526226
rect 273498 526170 273554 526226
rect 273622 526170 273678 526226
rect 273250 526046 273306 526102
rect 273374 526046 273430 526102
rect 273498 526046 273554 526102
rect 273622 526046 273678 526102
rect 273250 525922 273306 525978
rect 273374 525922 273430 525978
rect 273498 525922 273554 525978
rect 273622 525922 273678 525978
rect 273250 508294 273306 508350
rect 273374 508294 273430 508350
rect 273498 508294 273554 508350
rect 273622 508294 273678 508350
rect 273250 508170 273306 508226
rect 273374 508170 273430 508226
rect 273498 508170 273554 508226
rect 273622 508170 273678 508226
rect 273250 508046 273306 508102
rect 273374 508046 273430 508102
rect 273498 508046 273554 508102
rect 273622 508046 273678 508102
rect 273250 507922 273306 507978
rect 273374 507922 273430 507978
rect 273498 507922 273554 507978
rect 273622 507922 273678 507978
rect 276970 598116 277026 598172
rect 277094 598116 277150 598172
rect 277218 598116 277274 598172
rect 277342 598116 277398 598172
rect 276970 597992 277026 598048
rect 277094 597992 277150 598048
rect 277218 597992 277274 598048
rect 277342 597992 277398 598048
rect 276970 597868 277026 597924
rect 277094 597868 277150 597924
rect 277218 597868 277274 597924
rect 277342 597868 277398 597924
rect 276970 597744 277026 597800
rect 277094 597744 277150 597800
rect 277218 597744 277274 597800
rect 277342 597744 277398 597800
rect 276970 586294 277026 586350
rect 277094 586294 277150 586350
rect 277218 586294 277274 586350
rect 277342 586294 277398 586350
rect 276970 586170 277026 586226
rect 277094 586170 277150 586226
rect 277218 586170 277274 586226
rect 277342 586170 277398 586226
rect 276970 586046 277026 586102
rect 277094 586046 277150 586102
rect 277218 586046 277274 586102
rect 277342 586046 277398 586102
rect 276970 585922 277026 585978
rect 277094 585922 277150 585978
rect 277218 585922 277274 585978
rect 277342 585922 277398 585978
rect 276970 568294 277026 568350
rect 277094 568294 277150 568350
rect 277218 568294 277274 568350
rect 277342 568294 277398 568350
rect 276970 568170 277026 568226
rect 277094 568170 277150 568226
rect 277218 568170 277274 568226
rect 277342 568170 277398 568226
rect 276970 568046 277026 568102
rect 277094 568046 277150 568102
rect 277218 568046 277274 568102
rect 277342 568046 277398 568102
rect 276970 567922 277026 567978
rect 277094 567922 277150 567978
rect 277218 567922 277274 567978
rect 277342 567922 277398 567978
rect 276970 550294 277026 550350
rect 277094 550294 277150 550350
rect 277218 550294 277274 550350
rect 277342 550294 277398 550350
rect 276970 550170 277026 550226
rect 277094 550170 277150 550226
rect 277218 550170 277274 550226
rect 277342 550170 277398 550226
rect 276970 550046 277026 550102
rect 277094 550046 277150 550102
rect 277218 550046 277274 550102
rect 277342 550046 277398 550102
rect 276970 549922 277026 549978
rect 277094 549922 277150 549978
rect 277218 549922 277274 549978
rect 277342 549922 277398 549978
rect 276970 532294 277026 532350
rect 277094 532294 277150 532350
rect 277218 532294 277274 532350
rect 277342 532294 277398 532350
rect 276970 532170 277026 532226
rect 277094 532170 277150 532226
rect 277218 532170 277274 532226
rect 277342 532170 277398 532226
rect 276970 532046 277026 532102
rect 277094 532046 277150 532102
rect 277218 532046 277274 532102
rect 277342 532046 277398 532102
rect 276970 531922 277026 531978
rect 277094 531922 277150 531978
rect 277218 531922 277274 531978
rect 277342 531922 277398 531978
rect 276970 514294 277026 514350
rect 277094 514294 277150 514350
rect 277218 514294 277274 514350
rect 277342 514294 277398 514350
rect 276970 514170 277026 514226
rect 277094 514170 277150 514226
rect 277218 514170 277274 514226
rect 277342 514170 277398 514226
rect 276970 514046 277026 514102
rect 277094 514046 277150 514102
rect 277218 514046 277274 514102
rect 277342 514046 277398 514102
rect 276970 513922 277026 513978
rect 277094 513922 277150 513978
rect 277218 513922 277274 513978
rect 277342 513922 277398 513978
rect 291250 597156 291306 597212
rect 291374 597156 291430 597212
rect 291498 597156 291554 597212
rect 291622 597156 291678 597212
rect 291250 597032 291306 597088
rect 291374 597032 291430 597088
rect 291498 597032 291554 597088
rect 291622 597032 291678 597088
rect 291250 596908 291306 596964
rect 291374 596908 291430 596964
rect 291498 596908 291554 596964
rect 291622 596908 291678 596964
rect 291250 596784 291306 596840
rect 291374 596784 291430 596840
rect 291498 596784 291554 596840
rect 291622 596784 291678 596840
rect 291250 580294 291306 580350
rect 291374 580294 291430 580350
rect 291498 580294 291554 580350
rect 291622 580294 291678 580350
rect 291250 580170 291306 580226
rect 291374 580170 291430 580226
rect 291498 580170 291554 580226
rect 291622 580170 291678 580226
rect 291250 580046 291306 580102
rect 291374 580046 291430 580102
rect 291498 580046 291554 580102
rect 291622 580046 291678 580102
rect 291250 579922 291306 579978
rect 291374 579922 291430 579978
rect 291498 579922 291554 579978
rect 291622 579922 291678 579978
rect 291250 562294 291306 562350
rect 291374 562294 291430 562350
rect 291498 562294 291554 562350
rect 291622 562294 291678 562350
rect 291250 562170 291306 562226
rect 291374 562170 291430 562226
rect 291498 562170 291554 562226
rect 291622 562170 291678 562226
rect 291250 562046 291306 562102
rect 291374 562046 291430 562102
rect 291498 562046 291554 562102
rect 291622 562046 291678 562102
rect 291250 561922 291306 561978
rect 291374 561922 291430 561978
rect 291498 561922 291554 561978
rect 291622 561922 291678 561978
rect 291250 544294 291306 544350
rect 291374 544294 291430 544350
rect 291498 544294 291554 544350
rect 291622 544294 291678 544350
rect 291250 544170 291306 544226
rect 291374 544170 291430 544226
rect 291498 544170 291554 544226
rect 291622 544170 291678 544226
rect 291250 544046 291306 544102
rect 291374 544046 291430 544102
rect 291498 544046 291554 544102
rect 291622 544046 291678 544102
rect 291250 543922 291306 543978
rect 291374 543922 291430 543978
rect 291498 543922 291554 543978
rect 291622 543922 291678 543978
rect 291250 526294 291306 526350
rect 291374 526294 291430 526350
rect 291498 526294 291554 526350
rect 291622 526294 291678 526350
rect 291250 526170 291306 526226
rect 291374 526170 291430 526226
rect 291498 526170 291554 526226
rect 291622 526170 291678 526226
rect 291250 526046 291306 526102
rect 291374 526046 291430 526102
rect 291498 526046 291554 526102
rect 291622 526046 291678 526102
rect 291250 525922 291306 525978
rect 291374 525922 291430 525978
rect 291498 525922 291554 525978
rect 291622 525922 291678 525978
rect 291250 508294 291306 508350
rect 291374 508294 291430 508350
rect 291498 508294 291554 508350
rect 291622 508294 291678 508350
rect 291250 508170 291306 508226
rect 291374 508170 291430 508226
rect 291498 508170 291554 508226
rect 291622 508170 291678 508226
rect 291250 508046 291306 508102
rect 291374 508046 291430 508102
rect 291498 508046 291554 508102
rect 291622 508046 291678 508102
rect 291250 507922 291306 507978
rect 291374 507922 291430 507978
rect 291498 507922 291554 507978
rect 291622 507922 291678 507978
rect 294970 598116 295026 598172
rect 295094 598116 295150 598172
rect 295218 598116 295274 598172
rect 295342 598116 295398 598172
rect 294970 597992 295026 598048
rect 295094 597992 295150 598048
rect 295218 597992 295274 598048
rect 295342 597992 295398 598048
rect 294970 597868 295026 597924
rect 295094 597868 295150 597924
rect 295218 597868 295274 597924
rect 295342 597868 295398 597924
rect 294970 597744 295026 597800
rect 295094 597744 295150 597800
rect 295218 597744 295274 597800
rect 295342 597744 295398 597800
rect 294970 586294 295026 586350
rect 295094 586294 295150 586350
rect 295218 586294 295274 586350
rect 295342 586294 295398 586350
rect 294970 586170 295026 586226
rect 295094 586170 295150 586226
rect 295218 586170 295274 586226
rect 295342 586170 295398 586226
rect 294970 586046 295026 586102
rect 295094 586046 295150 586102
rect 295218 586046 295274 586102
rect 295342 586046 295398 586102
rect 294970 585922 295026 585978
rect 295094 585922 295150 585978
rect 295218 585922 295274 585978
rect 295342 585922 295398 585978
rect 294970 568294 295026 568350
rect 295094 568294 295150 568350
rect 295218 568294 295274 568350
rect 295342 568294 295398 568350
rect 294970 568170 295026 568226
rect 295094 568170 295150 568226
rect 295218 568170 295274 568226
rect 295342 568170 295398 568226
rect 294970 568046 295026 568102
rect 295094 568046 295150 568102
rect 295218 568046 295274 568102
rect 295342 568046 295398 568102
rect 294970 567922 295026 567978
rect 295094 567922 295150 567978
rect 295218 567922 295274 567978
rect 295342 567922 295398 567978
rect 294970 550294 295026 550350
rect 295094 550294 295150 550350
rect 295218 550294 295274 550350
rect 295342 550294 295398 550350
rect 294970 550170 295026 550226
rect 295094 550170 295150 550226
rect 295218 550170 295274 550226
rect 295342 550170 295398 550226
rect 294970 550046 295026 550102
rect 295094 550046 295150 550102
rect 295218 550046 295274 550102
rect 295342 550046 295398 550102
rect 294970 549922 295026 549978
rect 295094 549922 295150 549978
rect 295218 549922 295274 549978
rect 295342 549922 295398 549978
rect 294970 532294 295026 532350
rect 295094 532294 295150 532350
rect 295218 532294 295274 532350
rect 295342 532294 295398 532350
rect 294970 532170 295026 532226
rect 295094 532170 295150 532226
rect 295218 532170 295274 532226
rect 295342 532170 295398 532226
rect 294970 532046 295026 532102
rect 295094 532046 295150 532102
rect 295218 532046 295274 532102
rect 295342 532046 295398 532102
rect 294970 531922 295026 531978
rect 295094 531922 295150 531978
rect 295218 531922 295274 531978
rect 295342 531922 295398 531978
rect 294970 514294 295026 514350
rect 295094 514294 295150 514350
rect 295218 514294 295274 514350
rect 295342 514294 295398 514350
rect 294970 514170 295026 514226
rect 295094 514170 295150 514226
rect 295218 514170 295274 514226
rect 295342 514170 295398 514226
rect 294970 514046 295026 514102
rect 295094 514046 295150 514102
rect 295218 514046 295274 514102
rect 295342 514046 295398 514102
rect 294970 513922 295026 513978
rect 295094 513922 295150 513978
rect 295218 513922 295274 513978
rect 295342 513922 295398 513978
rect 309250 597156 309306 597212
rect 309374 597156 309430 597212
rect 309498 597156 309554 597212
rect 309622 597156 309678 597212
rect 309250 597032 309306 597088
rect 309374 597032 309430 597088
rect 309498 597032 309554 597088
rect 309622 597032 309678 597088
rect 309250 596908 309306 596964
rect 309374 596908 309430 596964
rect 309498 596908 309554 596964
rect 309622 596908 309678 596964
rect 309250 596784 309306 596840
rect 309374 596784 309430 596840
rect 309498 596784 309554 596840
rect 309622 596784 309678 596840
rect 309250 580294 309306 580350
rect 309374 580294 309430 580350
rect 309498 580294 309554 580350
rect 309622 580294 309678 580350
rect 309250 580170 309306 580226
rect 309374 580170 309430 580226
rect 309498 580170 309554 580226
rect 309622 580170 309678 580226
rect 309250 580046 309306 580102
rect 309374 580046 309430 580102
rect 309498 580046 309554 580102
rect 309622 580046 309678 580102
rect 309250 579922 309306 579978
rect 309374 579922 309430 579978
rect 309498 579922 309554 579978
rect 309622 579922 309678 579978
rect 309250 562294 309306 562350
rect 309374 562294 309430 562350
rect 309498 562294 309554 562350
rect 309622 562294 309678 562350
rect 309250 562170 309306 562226
rect 309374 562170 309430 562226
rect 309498 562170 309554 562226
rect 309622 562170 309678 562226
rect 309250 562046 309306 562102
rect 309374 562046 309430 562102
rect 309498 562046 309554 562102
rect 309622 562046 309678 562102
rect 309250 561922 309306 561978
rect 309374 561922 309430 561978
rect 309498 561922 309554 561978
rect 309622 561922 309678 561978
rect 309250 544294 309306 544350
rect 309374 544294 309430 544350
rect 309498 544294 309554 544350
rect 309622 544294 309678 544350
rect 309250 544170 309306 544226
rect 309374 544170 309430 544226
rect 309498 544170 309554 544226
rect 309622 544170 309678 544226
rect 309250 544046 309306 544102
rect 309374 544046 309430 544102
rect 309498 544046 309554 544102
rect 309622 544046 309678 544102
rect 309250 543922 309306 543978
rect 309374 543922 309430 543978
rect 309498 543922 309554 543978
rect 309622 543922 309678 543978
rect 309250 526294 309306 526350
rect 309374 526294 309430 526350
rect 309498 526294 309554 526350
rect 309622 526294 309678 526350
rect 309250 526170 309306 526226
rect 309374 526170 309430 526226
rect 309498 526170 309554 526226
rect 309622 526170 309678 526226
rect 309250 526046 309306 526102
rect 309374 526046 309430 526102
rect 309498 526046 309554 526102
rect 309622 526046 309678 526102
rect 309250 525922 309306 525978
rect 309374 525922 309430 525978
rect 309498 525922 309554 525978
rect 309622 525922 309678 525978
rect 309250 508294 309306 508350
rect 309374 508294 309430 508350
rect 309498 508294 309554 508350
rect 309622 508294 309678 508350
rect 309250 508170 309306 508226
rect 309374 508170 309430 508226
rect 309498 508170 309554 508226
rect 309622 508170 309678 508226
rect 309250 508046 309306 508102
rect 309374 508046 309430 508102
rect 309498 508046 309554 508102
rect 309622 508046 309678 508102
rect 309250 507922 309306 507978
rect 309374 507922 309430 507978
rect 309498 507922 309554 507978
rect 309622 507922 309678 507978
rect 312970 598116 313026 598172
rect 313094 598116 313150 598172
rect 313218 598116 313274 598172
rect 313342 598116 313398 598172
rect 312970 597992 313026 598048
rect 313094 597992 313150 598048
rect 313218 597992 313274 598048
rect 313342 597992 313398 598048
rect 312970 597868 313026 597924
rect 313094 597868 313150 597924
rect 313218 597868 313274 597924
rect 313342 597868 313398 597924
rect 312970 597744 313026 597800
rect 313094 597744 313150 597800
rect 313218 597744 313274 597800
rect 313342 597744 313398 597800
rect 312970 586294 313026 586350
rect 313094 586294 313150 586350
rect 313218 586294 313274 586350
rect 313342 586294 313398 586350
rect 312970 586170 313026 586226
rect 313094 586170 313150 586226
rect 313218 586170 313274 586226
rect 313342 586170 313398 586226
rect 312970 586046 313026 586102
rect 313094 586046 313150 586102
rect 313218 586046 313274 586102
rect 313342 586046 313398 586102
rect 312970 585922 313026 585978
rect 313094 585922 313150 585978
rect 313218 585922 313274 585978
rect 313342 585922 313398 585978
rect 312970 568294 313026 568350
rect 313094 568294 313150 568350
rect 313218 568294 313274 568350
rect 313342 568294 313398 568350
rect 312970 568170 313026 568226
rect 313094 568170 313150 568226
rect 313218 568170 313274 568226
rect 313342 568170 313398 568226
rect 312970 568046 313026 568102
rect 313094 568046 313150 568102
rect 313218 568046 313274 568102
rect 313342 568046 313398 568102
rect 312970 567922 313026 567978
rect 313094 567922 313150 567978
rect 313218 567922 313274 567978
rect 313342 567922 313398 567978
rect 312970 550294 313026 550350
rect 313094 550294 313150 550350
rect 313218 550294 313274 550350
rect 313342 550294 313398 550350
rect 312970 550170 313026 550226
rect 313094 550170 313150 550226
rect 313218 550170 313274 550226
rect 313342 550170 313398 550226
rect 312970 550046 313026 550102
rect 313094 550046 313150 550102
rect 313218 550046 313274 550102
rect 313342 550046 313398 550102
rect 312970 549922 313026 549978
rect 313094 549922 313150 549978
rect 313218 549922 313274 549978
rect 313342 549922 313398 549978
rect 312970 532294 313026 532350
rect 313094 532294 313150 532350
rect 313218 532294 313274 532350
rect 313342 532294 313398 532350
rect 312970 532170 313026 532226
rect 313094 532170 313150 532226
rect 313218 532170 313274 532226
rect 313342 532170 313398 532226
rect 312970 532046 313026 532102
rect 313094 532046 313150 532102
rect 313218 532046 313274 532102
rect 313342 532046 313398 532102
rect 312970 531922 313026 531978
rect 313094 531922 313150 531978
rect 313218 531922 313274 531978
rect 313342 531922 313398 531978
rect 312970 514294 313026 514350
rect 313094 514294 313150 514350
rect 313218 514294 313274 514350
rect 313342 514294 313398 514350
rect 312970 514170 313026 514226
rect 313094 514170 313150 514226
rect 313218 514170 313274 514226
rect 313342 514170 313398 514226
rect 312970 514046 313026 514102
rect 313094 514046 313150 514102
rect 313218 514046 313274 514102
rect 313342 514046 313398 514102
rect 312970 513922 313026 513978
rect 313094 513922 313150 513978
rect 313218 513922 313274 513978
rect 313342 513922 313398 513978
rect 327250 597156 327306 597212
rect 327374 597156 327430 597212
rect 327498 597156 327554 597212
rect 327622 597156 327678 597212
rect 327250 597032 327306 597088
rect 327374 597032 327430 597088
rect 327498 597032 327554 597088
rect 327622 597032 327678 597088
rect 327250 596908 327306 596964
rect 327374 596908 327430 596964
rect 327498 596908 327554 596964
rect 327622 596908 327678 596964
rect 327250 596784 327306 596840
rect 327374 596784 327430 596840
rect 327498 596784 327554 596840
rect 327622 596784 327678 596840
rect 327250 580294 327306 580350
rect 327374 580294 327430 580350
rect 327498 580294 327554 580350
rect 327622 580294 327678 580350
rect 327250 580170 327306 580226
rect 327374 580170 327430 580226
rect 327498 580170 327554 580226
rect 327622 580170 327678 580226
rect 327250 580046 327306 580102
rect 327374 580046 327430 580102
rect 327498 580046 327554 580102
rect 327622 580046 327678 580102
rect 327250 579922 327306 579978
rect 327374 579922 327430 579978
rect 327498 579922 327554 579978
rect 327622 579922 327678 579978
rect 327250 562294 327306 562350
rect 327374 562294 327430 562350
rect 327498 562294 327554 562350
rect 327622 562294 327678 562350
rect 327250 562170 327306 562226
rect 327374 562170 327430 562226
rect 327498 562170 327554 562226
rect 327622 562170 327678 562226
rect 327250 562046 327306 562102
rect 327374 562046 327430 562102
rect 327498 562046 327554 562102
rect 327622 562046 327678 562102
rect 327250 561922 327306 561978
rect 327374 561922 327430 561978
rect 327498 561922 327554 561978
rect 327622 561922 327678 561978
rect 327250 544294 327306 544350
rect 327374 544294 327430 544350
rect 327498 544294 327554 544350
rect 327622 544294 327678 544350
rect 327250 544170 327306 544226
rect 327374 544170 327430 544226
rect 327498 544170 327554 544226
rect 327622 544170 327678 544226
rect 327250 544046 327306 544102
rect 327374 544046 327430 544102
rect 327498 544046 327554 544102
rect 327622 544046 327678 544102
rect 327250 543922 327306 543978
rect 327374 543922 327430 543978
rect 327498 543922 327554 543978
rect 327622 543922 327678 543978
rect 327250 526294 327306 526350
rect 327374 526294 327430 526350
rect 327498 526294 327554 526350
rect 327622 526294 327678 526350
rect 327250 526170 327306 526226
rect 327374 526170 327430 526226
rect 327498 526170 327554 526226
rect 327622 526170 327678 526226
rect 327250 526046 327306 526102
rect 327374 526046 327430 526102
rect 327498 526046 327554 526102
rect 327622 526046 327678 526102
rect 327250 525922 327306 525978
rect 327374 525922 327430 525978
rect 327498 525922 327554 525978
rect 327622 525922 327678 525978
rect 327250 508294 327306 508350
rect 327374 508294 327430 508350
rect 327498 508294 327554 508350
rect 327622 508294 327678 508350
rect 327250 508170 327306 508226
rect 327374 508170 327430 508226
rect 327498 508170 327554 508226
rect 327622 508170 327678 508226
rect 327250 508046 327306 508102
rect 327374 508046 327430 508102
rect 327498 508046 327554 508102
rect 327622 508046 327678 508102
rect 327250 507922 327306 507978
rect 327374 507922 327430 507978
rect 327498 507922 327554 507978
rect 327622 507922 327678 507978
rect 330970 598116 331026 598172
rect 331094 598116 331150 598172
rect 331218 598116 331274 598172
rect 331342 598116 331398 598172
rect 330970 597992 331026 598048
rect 331094 597992 331150 598048
rect 331218 597992 331274 598048
rect 331342 597992 331398 598048
rect 330970 597868 331026 597924
rect 331094 597868 331150 597924
rect 331218 597868 331274 597924
rect 331342 597868 331398 597924
rect 330970 597744 331026 597800
rect 331094 597744 331150 597800
rect 331218 597744 331274 597800
rect 331342 597744 331398 597800
rect 330970 586294 331026 586350
rect 331094 586294 331150 586350
rect 331218 586294 331274 586350
rect 331342 586294 331398 586350
rect 330970 586170 331026 586226
rect 331094 586170 331150 586226
rect 331218 586170 331274 586226
rect 331342 586170 331398 586226
rect 330970 586046 331026 586102
rect 331094 586046 331150 586102
rect 331218 586046 331274 586102
rect 331342 586046 331398 586102
rect 330970 585922 331026 585978
rect 331094 585922 331150 585978
rect 331218 585922 331274 585978
rect 331342 585922 331398 585978
rect 330970 568294 331026 568350
rect 331094 568294 331150 568350
rect 331218 568294 331274 568350
rect 331342 568294 331398 568350
rect 330970 568170 331026 568226
rect 331094 568170 331150 568226
rect 331218 568170 331274 568226
rect 331342 568170 331398 568226
rect 330970 568046 331026 568102
rect 331094 568046 331150 568102
rect 331218 568046 331274 568102
rect 331342 568046 331398 568102
rect 330970 567922 331026 567978
rect 331094 567922 331150 567978
rect 331218 567922 331274 567978
rect 331342 567922 331398 567978
rect 330970 550294 331026 550350
rect 331094 550294 331150 550350
rect 331218 550294 331274 550350
rect 331342 550294 331398 550350
rect 330970 550170 331026 550226
rect 331094 550170 331150 550226
rect 331218 550170 331274 550226
rect 331342 550170 331398 550226
rect 330970 550046 331026 550102
rect 331094 550046 331150 550102
rect 331218 550046 331274 550102
rect 331342 550046 331398 550102
rect 330970 549922 331026 549978
rect 331094 549922 331150 549978
rect 331218 549922 331274 549978
rect 331342 549922 331398 549978
rect 330970 532294 331026 532350
rect 331094 532294 331150 532350
rect 331218 532294 331274 532350
rect 331342 532294 331398 532350
rect 330970 532170 331026 532226
rect 331094 532170 331150 532226
rect 331218 532170 331274 532226
rect 331342 532170 331398 532226
rect 330970 532046 331026 532102
rect 331094 532046 331150 532102
rect 331218 532046 331274 532102
rect 331342 532046 331398 532102
rect 330970 531922 331026 531978
rect 331094 531922 331150 531978
rect 331218 531922 331274 531978
rect 331342 531922 331398 531978
rect 330970 514294 331026 514350
rect 331094 514294 331150 514350
rect 331218 514294 331274 514350
rect 331342 514294 331398 514350
rect 330970 514170 331026 514226
rect 331094 514170 331150 514226
rect 331218 514170 331274 514226
rect 331342 514170 331398 514226
rect 330970 514046 331026 514102
rect 331094 514046 331150 514102
rect 331218 514046 331274 514102
rect 331342 514046 331398 514102
rect 330970 513922 331026 513978
rect 331094 513922 331150 513978
rect 331218 513922 331274 513978
rect 331342 513922 331398 513978
rect 345250 597156 345306 597212
rect 345374 597156 345430 597212
rect 345498 597156 345554 597212
rect 345622 597156 345678 597212
rect 345250 597032 345306 597088
rect 345374 597032 345430 597088
rect 345498 597032 345554 597088
rect 345622 597032 345678 597088
rect 345250 596908 345306 596964
rect 345374 596908 345430 596964
rect 345498 596908 345554 596964
rect 345622 596908 345678 596964
rect 345250 596784 345306 596840
rect 345374 596784 345430 596840
rect 345498 596784 345554 596840
rect 345622 596784 345678 596840
rect 345250 580294 345306 580350
rect 345374 580294 345430 580350
rect 345498 580294 345554 580350
rect 345622 580294 345678 580350
rect 345250 580170 345306 580226
rect 345374 580170 345430 580226
rect 345498 580170 345554 580226
rect 345622 580170 345678 580226
rect 345250 580046 345306 580102
rect 345374 580046 345430 580102
rect 345498 580046 345554 580102
rect 345622 580046 345678 580102
rect 345250 579922 345306 579978
rect 345374 579922 345430 579978
rect 345498 579922 345554 579978
rect 345622 579922 345678 579978
rect 345250 562294 345306 562350
rect 345374 562294 345430 562350
rect 345498 562294 345554 562350
rect 345622 562294 345678 562350
rect 345250 562170 345306 562226
rect 345374 562170 345430 562226
rect 345498 562170 345554 562226
rect 345622 562170 345678 562226
rect 345250 562046 345306 562102
rect 345374 562046 345430 562102
rect 345498 562046 345554 562102
rect 345622 562046 345678 562102
rect 345250 561922 345306 561978
rect 345374 561922 345430 561978
rect 345498 561922 345554 561978
rect 345622 561922 345678 561978
rect 345250 544294 345306 544350
rect 345374 544294 345430 544350
rect 345498 544294 345554 544350
rect 345622 544294 345678 544350
rect 345250 544170 345306 544226
rect 345374 544170 345430 544226
rect 345498 544170 345554 544226
rect 345622 544170 345678 544226
rect 345250 544046 345306 544102
rect 345374 544046 345430 544102
rect 345498 544046 345554 544102
rect 345622 544046 345678 544102
rect 345250 543922 345306 543978
rect 345374 543922 345430 543978
rect 345498 543922 345554 543978
rect 345622 543922 345678 543978
rect 345250 526294 345306 526350
rect 345374 526294 345430 526350
rect 345498 526294 345554 526350
rect 345622 526294 345678 526350
rect 345250 526170 345306 526226
rect 345374 526170 345430 526226
rect 345498 526170 345554 526226
rect 345622 526170 345678 526226
rect 345250 526046 345306 526102
rect 345374 526046 345430 526102
rect 345498 526046 345554 526102
rect 345622 526046 345678 526102
rect 345250 525922 345306 525978
rect 345374 525922 345430 525978
rect 345498 525922 345554 525978
rect 345622 525922 345678 525978
rect 345250 508294 345306 508350
rect 345374 508294 345430 508350
rect 345498 508294 345554 508350
rect 345622 508294 345678 508350
rect 345250 508170 345306 508226
rect 345374 508170 345430 508226
rect 345498 508170 345554 508226
rect 345622 508170 345678 508226
rect 345250 508046 345306 508102
rect 345374 508046 345430 508102
rect 345498 508046 345554 508102
rect 345622 508046 345678 508102
rect 345250 507922 345306 507978
rect 345374 507922 345430 507978
rect 345498 507922 345554 507978
rect 345622 507922 345678 507978
rect 348970 598116 349026 598172
rect 349094 598116 349150 598172
rect 349218 598116 349274 598172
rect 349342 598116 349398 598172
rect 348970 597992 349026 598048
rect 349094 597992 349150 598048
rect 349218 597992 349274 598048
rect 349342 597992 349398 598048
rect 348970 597868 349026 597924
rect 349094 597868 349150 597924
rect 349218 597868 349274 597924
rect 349342 597868 349398 597924
rect 348970 597744 349026 597800
rect 349094 597744 349150 597800
rect 349218 597744 349274 597800
rect 349342 597744 349398 597800
rect 348970 586294 349026 586350
rect 349094 586294 349150 586350
rect 349218 586294 349274 586350
rect 349342 586294 349398 586350
rect 348970 586170 349026 586226
rect 349094 586170 349150 586226
rect 349218 586170 349274 586226
rect 349342 586170 349398 586226
rect 348970 586046 349026 586102
rect 349094 586046 349150 586102
rect 349218 586046 349274 586102
rect 349342 586046 349398 586102
rect 348970 585922 349026 585978
rect 349094 585922 349150 585978
rect 349218 585922 349274 585978
rect 349342 585922 349398 585978
rect 348970 568294 349026 568350
rect 349094 568294 349150 568350
rect 349218 568294 349274 568350
rect 349342 568294 349398 568350
rect 348970 568170 349026 568226
rect 349094 568170 349150 568226
rect 349218 568170 349274 568226
rect 349342 568170 349398 568226
rect 348970 568046 349026 568102
rect 349094 568046 349150 568102
rect 349218 568046 349274 568102
rect 349342 568046 349398 568102
rect 348970 567922 349026 567978
rect 349094 567922 349150 567978
rect 349218 567922 349274 567978
rect 349342 567922 349398 567978
rect 348970 550294 349026 550350
rect 349094 550294 349150 550350
rect 349218 550294 349274 550350
rect 349342 550294 349398 550350
rect 348970 550170 349026 550226
rect 349094 550170 349150 550226
rect 349218 550170 349274 550226
rect 349342 550170 349398 550226
rect 348970 550046 349026 550102
rect 349094 550046 349150 550102
rect 349218 550046 349274 550102
rect 349342 550046 349398 550102
rect 348970 549922 349026 549978
rect 349094 549922 349150 549978
rect 349218 549922 349274 549978
rect 349342 549922 349398 549978
rect 348970 532294 349026 532350
rect 349094 532294 349150 532350
rect 349218 532294 349274 532350
rect 349342 532294 349398 532350
rect 348970 532170 349026 532226
rect 349094 532170 349150 532226
rect 349218 532170 349274 532226
rect 349342 532170 349398 532226
rect 348970 532046 349026 532102
rect 349094 532046 349150 532102
rect 349218 532046 349274 532102
rect 349342 532046 349398 532102
rect 348970 531922 349026 531978
rect 349094 531922 349150 531978
rect 349218 531922 349274 531978
rect 349342 531922 349398 531978
rect 348970 514294 349026 514350
rect 349094 514294 349150 514350
rect 349218 514294 349274 514350
rect 349342 514294 349398 514350
rect 348970 514170 349026 514226
rect 349094 514170 349150 514226
rect 349218 514170 349274 514226
rect 349342 514170 349398 514226
rect 348970 514046 349026 514102
rect 349094 514046 349150 514102
rect 349218 514046 349274 514102
rect 349342 514046 349398 514102
rect 348970 513922 349026 513978
rect 349094 513922 349150 513978
rect 349218 513922 349274 513978
rect 349342 513922 349398 513978
rect 363250 597156 363306 597212
rect 363374 597156 363430 597212
rect 363498 597156 363554 597212
rect 363622 597156 363678 597212
rect 363250 597032 363306 597088
rect 363374 597032 363430 597088
rect 363498 597032 363554 597088
rect 363622 597032 363678 597088
rect 363250 596908 363306 596964
rect 363374 596908 363430 596964
rect 363498 596908 363554 596964
rect 363622 596908 363678 596964
rect 363250 596784 363306 596840
rect 363374 596784 363430 596840
rect 363498 596784 363554 596840
rect 363622 596784 363678 596840
rect 363250 580294 363306 580350
rect 363374 580294 363430 580350
rect 363498 580294 363554 580350
rect 363622 580294 363678 580350
rect 363250 580170 363306 580226
rect 363374 580170 363430 580226
rect 363498 580170 363554 580226
rect 363622 580170 363678 580226
rect 363250 580046 363306 580102
rect 363374 580046 363430 580102
rect 363498 580046 363554 580102
rect 363622 580046 363678 580102
rect 363250 579922 363306 579978
rect 363374 579922 363430 579978
rect 363498 579922 363554 579978
rect 363622 579922 363678 579978
rect 363250 562294 363306 562350
rect 363374 562294 363430 562350
rect 363498 562294 363554 562350
rect 363622 562294 363678 562350
rect 363250 562170 363306 562226
rect 363374 562170 363430 562226
rect 363498 562170 363554 562226
rect 363622 562170 363678 562226
rect 363250 562046 363306 562102
rect 363374 562046 363430 562102
rect 363498 562046 363554 562102
rect 363622 562046 363678 562102
rect 363250 561922 363306 561978
rect 363374 561922 363430 561978
rect 363498 561922 363554 561978
rect 363622 561922 363678 561978
rect 363250 544294 363306 544350
rect 363374 544294 363430 544350
rect 363498 544294 363554 544350
rect 363622 544294 363678 544350
rect 363250 544170 363306 544226
rect 363374 544170 363430 544226
rect 363498 544170 363554 544226
rect 363622 544170 363678 544226
rect 363250 544046 363306 544102
rect 363374 544046 363430 544102
rect 363498 544046 363554 544102
rect 363622 544046 363678 544102
rect 363250 543922 363306 543978
rect 363374 543922 363430 543978
rect 363498 543922 363554 543978
rect 363622 543922 363678 543978
rect 363250 526294 363306 526350
rect 363374 526294 363430 526350
rect 363498 526294 363554 526350
rect 363622 526294 363678 526350
rect 363250 526170 363306 526226
rect 363374 526170 363430 526226
rect 363498 526170 363554 526226
rect 363622 526170 363678 526226
rect 363250 526046 363306 526102
rect 363374 526046 363430 526102
rect 363498 526046 363554 526102
rect 363622 526046 363678 526102
rect 363250 525922 363306 525978
rect 363374 525922 363430 525978
rect 363498 525922 363554 525978
rect 363622 525922 363678 525978
rect 363250 508294 363306 508350
rect 363374 508294 363430 508350
rect 363498 508294 363554 508350
rect 363622 508294 363678 508350
rect 363250 508170 363306 508226
rect 363374 508170 363430 508226
rect 363498 508170 363554 508226
rect 363622 508170 363678 508226
rect 363250 508046 363306 508102
rect 363374 508046 363430 508102
rect 363498 508046 363554 508102
rect 363622 508046 363678 508102
rect 363250 507922 363306 507978
rect 363374 507922 363430 507978
rect 363498 507922 363554 507978
rect 363622 507922 363678 507978
rect 366970 598116 367026 598172
rect 367094 598116 367150 598172
rect 367218 598116 367274 598172
rect 367342 598116 367398 598172
rect 366970 597992 367026 598048
rect 367094 597992 367150 598048
rect 367218 597992 367274 598048
rect 367342 597992 367398 598048
rect 366970 597868 367026 597924
rect 367094 597868 367150 597924
rect 367218 597868 367274 597924
rect 367342 597868 367398 597924
rect 366970 597744 367026 597800
rect 367094 597744 367150 597800
rect 367218 597744 367274 597800
rect 367342 597744 367398 597800
rect 366970 586294 367026 586350
rect 367094 586294 367150 586350
rect 367218 586294 367274 586350
rect 367342 586294 367398 586350
rect 366970 586170 367026 586226
rect 367094 586170 367150 586226
rect 367218 586170 367274 586226
rect 367342 586170 367398 586226
rect 366970 586046 367026 586102
rect 367094 586046 367150 586102
rect 367218 586046 367274 586102
rect 367342 586046 367398 586102
rect 366970 585922 367026 585978
rect 367094 585922 367150 585978
rect 367218 585922 367274 585978
rect 367342 585922 367398 585978
rect 366970 568294 367026 568350
rect 367094 568294 367150 568350
rect 367218 568294 367274 568350
rect 367342 568294 367398 568350
rect 366970 568170 367026 568226
rect 367094 568170 367150 568226
rect 367218 568170 367274 568226
rect 367342 568170 367398 568226
rect 366970 568046 367026 568102
rect 367094 568046 367150 568102
rect 367218 568046 367274 568102
rect 367342 568046 367398 568102
rect 366970 567922 367026 567978
rect 367094 567922 367150 567978
rect 367218 567922 367274 567978
rect 367342 567922 367398 567978
rect 366970 550294 367026 550350
rect 367094 550294 367150 550350
rect 367218 550294 367274 550350
rect 367342 550294 367398 550350
rect 366970 550170 367026 550226
rect 367094 550170 367150 550226
rect 367218 550170 367274 550226
rect 367342 550170 367398 550226
rect 366970 550046 367026 550102
rect 367094 550046 367150 550102
rect 367218 550046 367274 550102
rect 367342 550046 367398 550102
rect 366970 549922 367026 549978
rect 367094 549922 367150 549978
rect 367218 549922 367274 549978
rect 367342 549922 367398 549978
rect 366970 532294 367026 532350
rect 367094 532294 367150 532350
rect 367218 532294 367274 532350
rect 367342 532294 367398 532350
rect 366970 532170 367026 532226
rect 367094 532170 367150 532226
rect 367218 532170 367274 532226
rect 367342 532170 367398 532226
rect 366970 532046 367026 532102
rect 367094 532046 367150 532102
rect 367218 532046 367274 532102
rect 367342 532046 367398 532102
rect 366970 531922 367026 531978
rect 367094 531922 367150 531978
rect 367218 531922 367274 531978
rect 367342 531922 367398 531978
rect 366970 514294 367026 514350
rect 367094 514294 367150 514350
rect 367218 514294 367274 514350
rect 367342 514294 367398 514350
rect 366970 514170 367026 514226
rect 367094 514170 367150 514226
rect 367218 514170 367274 514226
rect 367342 514170 367398 514226
rect 366970 514046 367026 514102
rect 367094 514046 367150 514102
rect 367218 514046 367274 514102
rect 367342 514046 367398 514102
rect 366970 513922 367026 513978
rect 367094 513922 367150 513978
rect 367218 513922 367274 513978
rect 367342 513922 367398 513978
rect 381250 597156 381306 597212
rect 381374 597156 381430 597212
rect 381498 597156 381554 597212
rect 381622 597156 381678 597212
rect 381250 597032 381306 597088
rect 381374 597032 381430 597088
rect 381498 597032 381554 597088
rect 381622 597032 381678 597088
rect 381250 596908 381306 596964
rect 381374 596908 381430 596964
rect 381498 596908 381554 596964
rect 381622 596908 381678 596964
rect 381250 596784 381306 596840
rect 381374 596784 381430 596840
rect 381498 596784 381554 596840
rect 381622 596784 381678 596840
rect 381250 580294 381306 580350
rect 381374 580294 381430 580350
rect 381498 580294 381554 580350
rect 381622 580294 381678 580350
rect 381250 580170 381306 580226
rect 381374 580170 381430 580226
rect 381498 580170 381554 580226
rect 381622 580170 381678 580226
rect 381250 580046 381306 580102
rect 381374 580046 381430 580102
rect 381498 580046 381554 580102
rect 381622 580046 381678 580102
rect 381250 579922 381306 579978
rect 381374 579922 381430 579978
rect 381498 579922 381554 579978
rect 381622 579922 381678 579978
rect 381250 562294 381306 562350
rect 381374 562294 381430 562350
rect 381498 562294 381554 562350
rect 381622 562294 381678 562350
rect 381250 562170 381306 562226
rect 381374 562170 381430 562226
rect 381498 562170 381554 562226
rect 381622 562170 381678 562226
rect 381250 562046 381306 562102
rect 381374 562046 381430 562102
rect 381498 562046 381554 562102
rect 381622 562046 381678 562102
rect 381250 561922 381306 561978
rect 381374 561922 381430 561978
rect 381498 561922 381554 561978
rect 381622 561922 381678 561978
rect 381250 544294 381306 544350
rect 381374 544294 381430 544350
rect 381498 544294 381554 544350
rect 381622 544294 381678 544350
rect 381250 544170 381306 544226
rect 381374 544170 381430 544226
rect 381498 544170 381554 544226
rect 381622 544170 381678 544226
rect 381250 544046 381306 544102
rect 381374 544046 381430 544102
rect 381498 544046 381554 544102
rect 381622 544046 381678 544102
rect 381250 543922 381306 543978
rect 381374 543922 381430 543978
rect 381498 543922 381554 543978
rect 381622 543922 381678 543978
rect 381250 526294 381306 526350
rect 381374 526294 381430 526350
rect 381498 526294 381554 526350
rect 381622 526294 381678 526350
rect 381250 526170 381306 526226
rect 381374 526170 381430 526226
rect 381498 526170 381554 526226
rect 381622 526170 381678 526226
rect 381250 526046 381306 526102
rect 381374 526046 381430 526102
rect 381498 526046 381554 526102
rect 381622 526046 381678 526102
rect 381250 525922 381306 525978
rect 381374 525922 381430 525978
rect 381498 525922 381554 525978
rect 381622 525922 381678 525978
rect 381250 508294 381306 508350
rect 381374 508294 381430 508350
rect 381498 508294 381554 508350
rect 381622 508294 381678 508350
rect 381250 508170 381306 508226
rect 381374 508170 381430 508226
rect 381498 508170 381554 508226
rect 381622 508170 381678 508226
rect 381250 508046 381306 508102
rect 381374 508046 381430 508102
rect 381498 508046 381554 508102
rect 381622 508046 381678 508102
rect 381250 507922 381306 507978
rect 381374 507922 381430 507978
rect 381498 507922 381554 507978
rect 381622 507922 381678 507978
rect 384970 598116 385026 598172
rect 385094 598116 385150 598172
rect 385218 598116 385274 598172
rect 385342 598116 385398 598172
rect 384970 597992 385026 598048
rect 385094 597992 385150 598048
rect 385218 597992 385274 598048
rect 385342 597992 385398 598048
rect 384970 597868 385026 597924
rect 385094 597868 385150 597924
rect 385218 597868 385274 597924
rect 385342 597868 385398 597924
rect 384970 597744 385026 597800
rect 385094 597744 385150 597800
rect 385218 597744 385274 597800
rect 385342 597744 385398 597800
rect 384970 586294 385026 586350
rect 385094 586294 385150 586350
rect 385218 586294 385274 586350
rect 385342 586294 385398 586350
rect 384970 586170 385026 586226
rect 385094 586170 385150 586226
rect 385218 586170 385274 586226
rect 385342 586170 385398 586226
rect 384970 586046 385026 586102
rect 385094 586046 385150 586102
rect 385218 586046 385274 586102
rect 385342 586046 385398 586102
rect 384970 585922 385026 585978
rect 385094 585922 385150 585978
rect 385218 585922 385274 585978
rect 385342 585922 385398 585978
rect 384970 568294 385026 568350
rect 385094 568294 385150 568350
rect 385218 568294 385274 568350
rect 385342 568294 385398 568350
rect 384970 568170 385026 568226
rect 385094 568170 385150 568226
rect 385218 568170 385274 568226
rect 385342 568170 385398 568226
rect 384970 568046 385026 568102
rect 385094 568046 385150 568102
rect 385218 568046 385274 568102
rect 385342 568046 385398 568102
rect 384970 567922 385026 567978
rect 385094 567922 385150 567978
rect 385218 567922 385274 567978
rect 385342 567922 385398 567978
rect 384970 550294 385026 550350
rect 385094 550294 385150 550350
rect 385218 550294 385274 550350
rect 385342 550294 385398 550350
rect 384970 550170 385026 550226
rect 385094 550170 385150 550226
rect 385218 550170 385274 550226
rect 385342 550170 385398 550226
rect 384970 550046 385026 550102
rect 385094 550046 385150 550102
rect 385218 550046 385274 550102
rect 385342 550046 385398 550102
rect 384970 549922 385026 549978
rect 385094 549922 385150 549978
rect 385218 549922 385274 549978
rect 385342 549922 385398 549978
rect 384970 532294 385026 532350
rect 385094 532294 385150 532350
rect 385218 532294 385274 532350
rect 385342 532294 385398 532350
rect 384970 532170 385026 532226
rect 385094 532170 385150 532226
rect 385218 532170 385274 532226
rect 385342 532170 385398 532226
rect 384970 532046 385026 532102
rect 385094 532046 385150 532102
rect 385218 532046 385274 532102
rect 385342 532046 385398 532102
rect 384970 531922 385026 531978
rect 385094 531922 385150 531978
rect 385218 531922 385274 531978
rect 385342 531922 385398 531978
rect 384970 514294 385026 514350
rect 385094 514294 385150 514350
rect 385218 514294 385274 514350
rect 385342 514294 385398 514350
rect 384970 514170 385026 514226
rect 385094 514170 385150 514226
rect 385218 514170 385274 514226
rect 385342 514170 385398 514226
rect 384970 514046 385026 514102
rect 385094 514046 385150 514102
rect 385218 514046 385274 514102
rect 385342 514046 385398 514102
rect 384970 513922 385026 513978
rect 385094 513922 385150 513978
rect 385218 513922 385274 513978
rect 385342 513922 385398 513978
rect 399250 597156 399306 597212
rect 399374 597156 399430 597212
rect 399498 597156 399554 597212
rect 399622 597156 399678 597212
rect 399250 597032 399306 597088
rect 399374 597032 399430 597088
rect 399498 597032 399554 597088
rect 399622 597032 399678 597088
rect 399250 596908 399306 596964
rect 399374 596908 399430 596964
rect 399498 596908 399554 596964
rect 399622 596908 399678 596964
rect 399250 596784 399306 596840
rect 399374 596784 399430 596840
rect 399498 596784 399554 596840
rect 399622 596784 399678 596840
rect 399250 580294 399306 580350
rect 399374 580294 399430 580350
rect 399498 580294 399554 580350
rect 399622 580294 399678 580350
rect 399250 580170 399306 580226
rect 399374 580170 399430 580226
rect 399498 580170 399554 580226
rect 399622 580170 399678 580226
rect 399250 580046 399306 580102
rect 399374 580046 399430 580102
rect 399498 580046 399554 580102
rect 399622 580046 399678 580102
rect 399250 579922 399306 579978
rect 399374 579922 399430 579978
rect 399498 579922 399554 579978
rect 399622 579922 399678 579978
rect 399250 562294 399306 562350
rect 399374 562294 399430 562350
rect 399498 562294 399554 562350
rect 399622 562294 399678 562350
rect 399250 562170 399306 562226
rect 399374 562170 399430 562226
rect 399498 562170 399554 562226
rect 399622 562170 399678 562226
rect 399250 562046 399306 562102
rect 399374 562046 399430 562102
rect 399498 562046 399554 562102
rect 399622 562046 399678 562102
rect 399250 561922 399306 561978
rect 399374 561922 399430 561978
rect 399498 561922 399554 561978
rect 399622 561922 399678 561978
rect 399250 544294 399306 544350
rect 399374 544294 399430 544350
rect 399498 544294 399554 544350
rect 399622 544294 399678 544350
rect 399250 544170 399306 544226
rect 399374 544170 399430 544226
rect 399498 544170 399554 544226
rect 399622 544170 399678 544226
rect 399250 544046 399306 544102
rect 399374 544046 399430 544102
rect 399498 544046 399554 544102
rect 399622 544046 399678 544102
rect 399250 543922 399306 543978
rect 399374 543922 399430 543978
rect 399498 543922 399554 543978
rect 399622 543922 399678 543978
rect 399250 526294 399306 526350
rect 399374 526294 399430 526350
rect 399498 526294 399554 526350
rect 399622 526294 399678 526350
rect 399250 526170 399306 526226
rect 399374 526170 399430 526226
rect 399498 526170 399554 526226
rect 399622 526170 399678 526226
rect 399250 526046 399306 526102
rect 399374 526046 399430 526102
rect 399498 526046 399554 526102
rect 399622 526046 399678 526102
rect 399250 525922 399306 525978
rect 399374 525922 399430 525978
rect 399498 525922 399554 525978
rect 399622 525922 399678 525978
rect 399250 508294 399306 508350
rect 399374 508294 399430 508350
rect 399498 508294 399554 508350
rect 399622 508294 399678 508350
rect 399250 508170 399306 508226
rect 399374 508170 399430 508226
rect 399498 508170 399554 508226
rect 399622 508170 399678 508226
rect 399250 508046 399306 508102
rect 399374 508046 399430 508102
rect 399498 508046 399554 508102
rect 399622 508046 399678 508102
rect 399250 507922 399306 507978
rect 399374 507922 399430 507978
rect 399498 507922 399554 507978
rect 399622 507922 399678 507978
rect 402970 598116 403026 598172
rect 403094 598116 403150 598172
rect 403218 598116 403274 598172
rect 403342 598116 403398 598172
rect 402970 597992 403026 598048
rect 403094 597992 403150 598048
rect 403218 597992 403274 598048
rect 403342 597992 403398 598048
rect 402970 597868 403026 597924
rect 403094 597868 403150 597924
rect 403218 597868 403274 597924
rect 403342 597868 403398 597924
rect 402970 597744 403026 597800
rect 403094 597744 403150 597800
rect 403218 597744 403274 597800
rect 403342 597744 403398 597800
rect 402970 586294 403026 586350
rect 403094 586294 403150 586350
rect 403218 586294 403274 586350
rect 403342 586294 403398 586350
rect 402970 586170 403026 586226
rect 403094 586170 403150 586226
rect 403218 586170 403274 586226
rect 403342 586170 403398 586226
rect 402970 586046 403026 586102
rect 403094 586046 403150 586102
rect 403218 586046 403274 586102
rect 403342 586046 403398 586102
rect 402970 585922 403026 585978
rect 403094 585922 403150 585978
rect 403218 585922 403274 585978
rect 403342 585922 403398 585978
rect 402970 568294 403026 568350
rect 403094 568294 403150 568350
rect 403218 568294 403274 568350
rect 403342 568294 403398 568350
rect 402970 568170 403026 568226
rect 403094 568170 403150 568226
rect 403218 568170 403274 568226
rect 403342 568170 403398 568226
rect 402970 568046 403026 568102
rect 403094 568046 403150 568102
rect 403218 568046 403274 568102
rect 403342 568046 403398 568102
rect 402970 567922 403026 567978
rect 403094 567922 403150 567978
rect 403218 567922 403274 567978
rect 403342 567922 403398 567978
rect 402970 550294 403026 550350
rect 403094 550294 403150 550350
rect 403218 550294 403274 550350
rect 403342 550294 403398 550350
rect 402970 550170 403026 550226
rect 403094 550170 403150 550226
rect 403218 550170 403274 550226
rect 403342 550170 403398 550226
rect 402970 550046 403026 550102
rect 403094 550046 403150 550102
rect 403218 550046 403274 550102
rect 403342 550046 403398 550102
rect 402970 549922 403026 549978
rect 403094 549922 403150 549978
rect 403218 549922 403274 549978
rect 403342 549922 403398 549978
rect 402970 532294 403026 532350
rect 403094 532294 403150 532350
rect 403218 532294 403274 532350
rect 403342 532294 403398 532350
rect 402970 532170 403026 532226
rect 403094 532170 403150 532226
rect 403218 532170 403274 532226
rect 403342 532170 403398 532226
rect 402970 532046 403026 532102
rect 403094 532046 403150 532102
rect 403218 532046 403274 532102
rect 403342 532046 403398 532102
rect 402970 531922 403026 531978
rect 403094 531922 403150 531978
rect 403218 531922 403274 531978
rect 403342 531922 403398 531978
rect 402970 514294 403026 514350
rect 403094 514294 403150 514350
rect 403218 514294 403274 514350
rect 403342 514294 403398 514350
rect 402970 514170 403026 514226
rect 403094 514170 403150 514226
rect 403218 514170 403274 514226
rect 403342 514170 403398 514226
rect 402970 514046 403026 514102
rect 403094 514046 403150 514102
rect 403218 514046 403274 514102
rect 403342 514046 403398 514102
rect 402970 513922 403026 513978
rect 403094 513922 403150 513978
rect 403218 513922 403274 513978
rect 403342 513922 403398 513978
rect 417250 597156 417306 597212
rect 417374 597156 417430 597212
rect 417498 597156 417554 597212
rect 417622 597156 417678 597212
rect 417250 597032 417306 597088
rect 417374 597032 417430 597088
rect 417498 597032 417554 597088
rect 417622 597032 417678 597088
rect 417250 596908 417306 596964
rect 417374 596908 417430 596964
rect 417498 596908 417554 596964
rect 417622 596908 417678 596964
rect 417250 596784 417306 596840
rect 417374 596784 417430 596840
rect 417498 596784 417554 596840
rect 417622 596784 417678 596840
rect 417250 580294 417306 580350
rect 417374 580294 417430 580350
rect 417498 580294 417554 580350
rect 417622 580294 417678 580350
rect 417250 580170 417306 580226
rect 417374 580170 417430 580226
rect 417498 580170 417554 580226
rect 417622 580170 417678 580226
rect 417250 580046 417306 580102
rect 417374 580046 417430 580102
rect 417498 580046 417554 580102
rect 417622 580046 417678 580102
rect 417250 579922 417306 579978
rect 417374 579922 417430 579978
rect 417498 579922 417554 579978
rect 417622 579922 417678 579978
rect 417250 562294 417306 562350
rect 417374 562294 417430 562350
rect 417498 562294 417554 562350
rect 417622 562294 417678 562350
rect 417250 562170 417306 562226
rect 417374 562170 417430 562226
rect 417498 562170 417554 562226
rect 417622 562170 417678 562226
rect 417250 562046 417306 562102
rect 417374 562046 417430 562102
rect 417498 562046 417554 562102
rect 417622 562046 417678 562102
rect 417250 561922 417306 561978
rect 417374 561922 417430 561978
rect 417498 561922 417554 561978
rect 417622 561922 417678 561978
rect 417250 544294 417306 544350
rect 417374 544294 417430 544350
rect 417498 544294 417554 544350
rect 417622 544294 417678 544350
rect 417250 544170 417306 544226
rect 417374 544170 417430 544226
rect 417498 544170 417554 544226
rect 417622 544170 417678 544226
rect 417250 544046 417306 544102
rect 417374 544046 417430 544102
rect 417498 544046 417554 544102
rect 417622 544046 417678 544102
rect 417250 543922 417306 543978
rect 417374 543922 417430 543978
rect 417498 543922 417554 543978
rect 417622 543922 417678 543978
rect 417250 526294 417306 526350
rect 417374 526294 417430 526350
rect 417498 526294 417554 526350
rect 417622 526294 417678 526350
rect 417250 526170 417306 526226
rect 417374 526170 417430 526226
rect 417498 526170 417554 526226
rect 417622 526170 417678 526226
rect 417250 526046 417306 526102
rect 417374 526046 417430 526102
rect 417498 526046 417554 526102
rect 417622 526046 417678 526102
rect 417250 525922 417306 525978
rect 417374 525922 417430 525978
rect 417498 525922 417554 525978
rect 417622 525922 417678 525978
rect 417250 508294 417306 508350
rect 417374 508294 417430 508350
rect 417498 508294 417554 508350
rect 417622 508294 417678 508350
rect 417250 508170 417306 508226
rect 417374 508170 417430 508226
rect 417498 508170 417554 508226
rect 417622 508170 417678 508226
rect 417250 508046 417306 508102
rect 417374 508046 417430 508102
rect 417498 508046 417554 508102
rect 417622 508046 417678 508102
rect 417250 507922 417306 507978
rect 417374 507922 417430 507978
rect 417498 507922 417554 507978
rect 417622 507922 417678 507978
rect 420970 598116 421026 598172
rect 421094 598116 421150 598172
rect 421218 598116 421274 598172
rect 421342 598116 421398 598172
rect 420970 597992 421026 598048
rect 421094 597992 421150 598048
rect 421218 597992 421274 598048
rect 421342 597992 421398 598048
rect 420970 597868 421026 597924
rect 421094 597868 421150 597924
rect 421218 597868 421274 597924
rect 421342 597868 421398 597924
rect 420970 597744 421026 597800
rect 421094 597744 421150 597800
rect 421218 597744 421274 597800
rect 421342 597744 421398 597800
rect 420970 586294 421026 586350
rect 421094 586294 421150 586350
rect 421218 586294 421274 586350
rect 421342 586294 421398 586350
rect 420970 586170 421026 586226
rect 421094 586170 421150 586226
rect 421218 586170 421274 586226
rect 421342 586170 421398 586226
rect 420970 586046 421026 586102
rect 421094 586046 421150 586102
rect 421218 586046 421274 586102
rect 421342 586046 421398 586102
rect 420970 585922 421026 585978
rect 421094 585922 421150 585978
rect 421218 585922 421274 585978
rect 421342 585922 421398 585978
rect 420970 568294 421026 568350
rect 421094 568294 421150 568350
rect 421218 568294 421274 568350
rect 421342 568294 421398 568350
rect 420970 568170 421026 568226
rect 421094 568170 421150 568226
rect 421218 568170 421274 568226
rect 421342 568170 421398 568226
rect 420970 568046 421026 568102
rect 421094 568046 421150 568102
rect 421218 568046 421274 568102
rect 421342 568046 421398 568102
rect 420970 567922 421026 567978
rect 421094 567922 421150 567978
rect 421218 567922 421274 567978
rect 421342 567922 421398 567978
rect 420970 550294 421026 550350
rect 421094 550294 421150 550350
rect 421218 550294 421274 550350
rect 421342 550294 421398 550350
rect 420970 550170 421026 550226
rect 421094 550170 421150 550226
rect 421218 550170 421274 550226
rect 421342 550170 421398 550226
rect 420970 550046 421026 550102
rect 421094 550046 421150 550102
rect 421218 550046 421274 550102
rect 421342 550046 421398 550102
rect 420970 549922 421026 549978
rect 421094 549922 421150 549978
rect 421218 549922 421274 549978
rect 421342 549922 421398 549978
rect 420970 532294 421026 532350
rect 421094 532294 421150 532350
rect 421218 532294 421274 532350
rect 421342 532294 421398 532350
rect 420970 532170 421026 532226
rect 421094 532170 421150 532226
rect 421218 532170 421274 532226
rect 421342 532170 421398 532226
rect 420970 532046 421026 532102
rect 421094 532046 421150 532102
rect 421218 532046 421274 532102
rect 421342 532046 421398 532102
rect 420970 531922 421026 531978
rect 421094 531922 421150 531978
rect 421218 531922 421274 531978
rect 421342 531922 421398 531978
rect 420970 514294 421026 514350
rect 421094 514294 421150 514350
rect 421218 514294 421274 514350
rect 421342 514294 421398 514350
rect 420970 514170 421026 514226
rect 421094 514170 421150 514226
rect 421218 514170 421274 514226
rect 421342 514170 421398 514226
rect 420970 514046 421026 514102
rect 421094 514046 421150 514102
rect 421218 514046 421274 514102
rect 421342 514046 421398 514102
rect 420970 513922 421026 513978
rect 421094 513922 421150 513978
rect 421218 513922 421274 513978
rect 421342 513922 421398 513978
rect 435250 597156 435306 597212
rect 435374 597156 435430 597212
rect 435498 597156 435554 597212
rect 435622 597156 435678 597212
rect 435250 597032 435306 597088
rect 435374 597032 435430 597088
rect 435498 597032 435554 597088
rect 435622 597032 435678 597088
rect 435250 596908 435306 596964
rect 435374 596908 435430 596964
rect 435498 596908 435554 596964
rect 435622 596908 435678 596964
rect 435250 596784 435306 596840
rect 435374 596784 435430 596840
rect 435498 596784 435554 596840
rect 435622 596784 435678 596840
rect 435250 580294 435306 580350
rect 435374 580294 435430 580350
rect 435498 580294 435554 580350
rect 435622 580294 435678 580350
rect 435250 580170 435306 580226
rect 435374 580170 435430 580226
rect 435498 580170 435554 580226
rect 435622 580170 435678 580226
rect 435250 580046 435306 580102
rect 435374 580046 435430 580102
rect 435498 580046 435554 580102
rect 435622 580046 435678 580102
rect 435250 579922 435306 579978
rect 435374 579922 435430 579978
rect 435498 579922 435554 579978
rect 435622 579922 435678 579978
rect 435250 562294 435306 562350
rect 435374 562294 435430 562350
rect 435498 562294 435554 562350
rect 435622 562294 435678 562350
rect 435250 562170 435306 562226
rect 435374 562170 435430 562226
rect 435498 562170 435554 562226
rect 435622 562170 435678 562226
rect 435250 562046 435306 562102
rect 435374 562046 435430 562102
rect 435498 562046 435554 562102
rect 435622 562046 435678 562102
rect 435250 561922 435306 561978
rect 435374 561922 435430 561978
rect 435498 561922 435554 561978
rect 435622 561922 435678 561978
rect 435250 544294 435306 544350
rect 435374 544294 435430 544350
rect 435498 544294 435554 544350
rect 435622 544294 435678 544350
rect 435250 544170 435306 544226
rect 435374 544170 435430 544226
rect 435498 544170 435554 544226
rect 435622 544170 435678 544226
rect 435250 544046 435306 544102
rect 435374 544046 435430 544102
rect 435498 544046 435554 544102
rect 435622 544046 435678 544102
rect 435250 543922 435306 543978
rect 435374 543922 435430 543978
rect 435498 543922 435554 543978
rect 435622 543922 435678 543978
rect 435250 526294 435306 526350
rect 435374 526294 435430 526350
rect 435498 526294 435554 526350
rect 435622 526294 435678 526350
rect 435250 526170 435306 526226
rect 435374 526170 435430 526226
rect 435498 526170 435554 526226
rect 435622 526170 435678 526226
rect 435250 526046 435306 526102
rect 435374 526046 435430 526102
rect 435498 526046 435554 526102
rect 435622 526046 435678 526102
rect 435250 525922 435306 525978
rect 435374 525922 435430 525978
rect 435498 525922 435554 525978
rect 435622 525922 435678 525978
rect 435250 508294 435306 508350
rect 435374 508294 435430 508350
rect 435498 508294 435554 508350
rect 435622 508294 435678 508350
rect 435250 508170 435306 508226
rect 435374 508170 435430 508226
rect 435498 508170 435554 508226
rect 435622 508170 435678 508226
rect 435250 508046 435306 508102
rect 435374 508046 435430 508102
rect 435498 508046 435554 508102
rect 435622 508046 435678 508102
rect 435250 507922 435306 507978
rect 435374 507922 435430 507978
rect 435498 507922 435554 507978
rect 435622 507922 435678 507978
rect 438970 598116 439026 598172
rect 439094 598116 439150 598172
rect 439218 598116 439274 598172
rect 439342 598116 439398 598172
rect 438970 597992 439026 598048
rect 439094 597992 439150 598048
rect 439218 597992 439274 598048
rect 439342 597992 439398 598048
rect 438970 597868 439026 597924
rect 439094 597868 439150 597924
rect 439218 597868 439274 597924
rect 439342 597868 439398 597924
rect 438970 597744 439026 597800
rect 439094 597744 439150 597800
rect 439218 597744 439274 597800
rect 439342 597744 439398 597800
rect 438970 586294 439026 586350
rect 439094 586294 439150 586350
rect 439218 586294 439274 586350
rect 439342 586294 439398 586350
rect 438970 586170 439026 586226
rect 439094 586170 439150 586226
rect 439218 586170 439274 586226
rect 439342 586170 439398 586226
rect 438970 586046 439026 586102
rect 439094 586046 439150 586102
rect 439218 586046 439274 586102
rect 439342 586046 439398 586102
rect 438970 585922 439026 585978
rect 439094 585922 439150 585978
rect 439218 585922 439274 585978
rect 439342 585922 439398 585978
rect 438970 568294 439026 568350
rect 439094 568294 439150 568350
rect 439218 568294 439274 568350
rect 439342 568294 439398 568350
rect 438970 568170 439026 568226
rect 439094 568170 439150 568226
rect 439218 568170 439274 568226
rect 439342 568170 439398 568226
rect 438970 568046 439026 568102
rect 439094 568046 439150 568102
rect 439218 568046 439274 568102
rect 439342 568046 439398 568102
rect 438970 567922 439026 567978
rect 439094 567922 439150 567978
rect 439218 567922 439274 567978
rect 439342 567922 439398 567978
rect 438970 550294 439026 550350
rect 439094 550294 439150 550350
rect 439218 550294 439274 550350
rect 439342 550294 439398 550350
rect 438970 550170 439026 550226
rect 439094 550170 439150 550226
rect 439218 550170 439274 550226
rect 439342 550170 439398 550226
rect 438970 550046 439026 550102
rect 439094 550046 439150 550102
rect 439218 550046 439274 550102
rect 439342 550046 439398 550102
rect 438970 549922 439026 549978
rect 439094 549922 439150 549978
rect 439218 549922 439274 549978
rect 439342 549922 439398 549978
rect 438970 532294 439026 532350
rect 439094 532294 439150 532350
rect 439218 532294 439274 532350
rect 439342 532294 439398 532350
rect 438970 532170 439026 532226
rect 439094 532170 439150 532226
rect 439218 532170 439274 532226
rect 439342 532170 439398 532226
rect 438970 532046 439026 532102
rect 439094 532046 439150 532102
rect 439218 532046 439274 532102
rect 439342 532046 439398 532102
rect 438970 531922 439026 531978
rect 439094 531922 439150 531978
rect 439218 531922 439274 531978
rect 439342 531922 439398 531978
rect 438970 514294 439026 514350
rect 439094 514294 439150 514350
rect 439218 514294 439274 514350
rect 439342 514294 439398 514350
rect 438970 514170 439026 514226
rect 439094 514170 439150 514226
rect 439218 514170 439274 514226
rect 439342 514170 439398 514226
rect 438970 514046 439026 514102
rect 439094 514046 439150 514102
rect 439218 514046 439274 514102
rect 439342 514046 439398 514102
rect 438970 513922 439026 513978
rect 439094 513922 439150 513978
rect 439218 513922 439274 513978
rect 439342 513922 439398 513978
rect 453250 597156 453306 597212
rect 453374 597156 453430 597212
rect 453498 597156 453554 597212
rect 453622 597156 453678 597212
rect 453250 597032 453306 597088
rect 453374 597032 453430 597088
rect 453498 597032 453554 597088
rect 453622 597032 453678 597088
rect 453250 596908 453306 596964
rect 453374 596908 453430 596964
rect 453498 596908 453554 596964
rect 453622 596908 453678 596964
rect 453250 596784 453306 596840
rect 453374 596784 453430 596840
rect 453498 596784 453554 596840
rect 453622 596784 453678 596840
rect 453250 580294 453306 580350
rect 453374 580294 453430 580350
rect 453498 580294 453554 580350
rect 453622 580294 453678 580350
rect 453250 580170 453306 580226
rect 453374 580170 453430 580226
rect 453498 580170 453554 580226
rect 453622 580170 453678 580226
rect 453250 580046 453306 580102
rect 453374 580046 453430 580102
rect 453498 580046 453554 580102
rect 453622 580046 453678 580102
rect 453250 579922 453306 579978
rect 453374 579922 453430 579978
rect 453498 579922 453554 579978
rect 453622 579922 453678 579978
rect 453250 562294 453306 562350
rect 453374 562294 453430 562350
rect 453498 562294 453554 562350
rect 453622 562294 453678 562350
rect 453250 562170 453306 562226
rect 453374 562170 453430 562226
rect 453498 562170 453554 562226
rect 453622 562170 453678 562226
rect 453250 562046 453306 562102
rect 453374 562046 453430 562102
rect 453498 562046 453554 562102
rect 453622 562046 453678 562102
rect 453250 561922 453306 561978
rect 453374 561922 453430 561978
rect 453498 561922 453554 561978
rect 453622 561922 453678 561978
rect 453250 544294 453306 544350
rect 453374 544294 453430 544350
rect 453498 544294 453554 544350
rect 453622 544294 453678 544350
rect 453250 544170 453306 544226
rect 453374 544170 453430 544226
rect 453498 544170 453554 544226
rect 453622 544170 453678 544226
rect 453250 544046 453306 544102
rect 453374 544046 453430 544102
rect 453498 544046 453554 544102
rect 453622 544046 453678 544102
rect 453250 543922 453306 543978
rect 453374 543922 453430 543978
rect 453498 543922 453554 543978
rect 453622 543922 453678 543978
rect 453250 526294 453306 526350
rect 453374 526294 453430 526350
rect 453498 526294 453554 526350
rect 453622 526294 453678 526350
rect 453250 526170 453306 526226
rect 453374 526170 453430 526226
rect 453498 526170 453554 526226
rect 453622 526170 453678 526226
rect 453250 526046 453306 526102
rect 453374 526046 453430 526102
rect 453498 526046 453554 526102
rect 453622 526046 453678 526102
rect 453250 525922 453306 525978
rect 453374 525922 453430 525978
rect 453498 525922 453554 525978
rect 453622 525922 453678 525978
rect 453250 508294 453306 508350
rect 453374 508294 453430 508350
rect 453498 508294 453554 508350
rect 453622 508294 453678 508350
rect 453250 508170 453306 508226
rect 453374 508170 453430 508226
rect 453498 508170 453554 508226
rect 453622 508170 453678 508226
rect 453250 508046 453306 508102
rect 453374 508046 453430 508102
rect 453498 508046 453554 508102
rect 453622 508046 453678 508102
rect 453250 507922 453306 507978
rect 453374 507922 453430 507978
rect 453498 507922 453554 507978
rect 453622 507922 453678 507978
rect 456970 598116 457026 598172
rect 457094 598116 457150 598172
rect 457218 598116 457274 598172
rect 457342 598116 457398 598172
rect 456970 597992 457026 598048
rect 457094 597992 457150 598048
rect 457218 597992 457274 598048
rect 457342 597992 457398 598048
rect 456970 597868 457026 597924
rect 457094 597868 457150 597924
rect 457218 597868 457274 597924
rect 457342 597868 457398 597924
rect 456970 597744 457026 597800
rect 457094 597744 457150 597800
rect 457218 597744 457274 597800
rect 457342 597744 457398 597800
rect 456970 586294 457026 586350
rect 457094 586294 457150 586350
rect 457218 586294 457274 586350
rect 457342 586294 457398 586350
rect 456970 586170 457026 586226
rect 457094 586170 457150 586226
rect 457218 586170 457274 586226
rect 457342 586170 457398 586226
rect 456970 586046 457026 586102
rect 457094 586046 457150 586102
rect 457218 586046 457274 586102
rect 457342 586046 457398 586102
rect 456970 585922 457026 585978
rect 457094 585922 457150 585978
rect 457218 585922 457274 585978
rect 457342 585922 457398 585978
rect 456970 568294 457026 568350
rect 457094 568294 457150 568350
rect 457218 568294 457274 568350
rect 457342 568294 457398 568350
rect 456970 568170 457026 568226
rect 457094 568170 457150 568226
rect 457218 568170 457274 568226
rect 457342 568170 457398 568226
rect 456970 568046 457026 568102
rect 457094 568046 457150 568102
rect 457218 568046 457274 568102
rect 457342 568046 457398 568102
rect 456970 567922 457026 567978
rect 457094 567922 457150 567978
rect 457218 567922 457274 567978
rect 457342 567922 457398 567978
rect 456970 550294 457026 550350
rect 457094 550294 457150 550350
rect 457218 550294 457274 550350
rect 457342 550294 457398 550350
rect 456970 550170 457026 550226
rect 457094 550170 457150 550226
rect 457218 550170 457274 550226
rect 457342 550170 457398 550226
rect 456970 550046 457026 550102
rect 457094 550046 457150 550102
rect 457218 550046 457274 550102
rect 457342 550046 457398 550102
rect 456970 549922 457026 549978
rect 457094 549922 457150 549978
rect 457218 549922 457274 549978
rect 457342 549922 457398 549978
rect 456970 532294 457026 532350
rect 457094 532294 457150 532350
rect 457218 532294 457274 532350
rect 457342 532294 457398 532350
rect 456970 532170 457026 532226
rect 457094 532170 457150 532226
rect 457218 532170 457274 532226
rect 457342 532170 457398 532226
rect 456970 532046 457026 532102
rect 457094 532046 457150 532102
rect 457218 532046 457274 532102
rect 457342 532046 457398 532102
rect 456970 531922 457026 531978
rect 457094 531922 457150 531978
rect 457218 531922 457274 531978
rect 457342 531922 457398 531978
rect 456970 514294 457026 514350
rect 457094 514294 457150 514350
rect 457218 514294 457274 514350
rect 457342 514294 457398 514350
rect 456970 514170 457026 514226
rect 457094 514170 457150 514226
rect 457218 514170 457274 514226
rect 457342 514170 457398 514226
rect 456970 514046 457026 514102
rect 457094 514046 457150 514102
rect 457218 514046 457274 514102
rect 457342 514046 457398 514102
rect 456970 513922 457026 513978
rect 457094 513922 457150 513978
rect 457218 513922 457274 513978
rect 457342 513922 457398 513978
rect 471250 597156 471306 597212
rect 471374 597156 471430 597212
rect 471498 597156 471554 597212
rect 471622 597156 471678 597212
rect 471250 597032 471306 597088
rect 471374 597032 471430 597088
rect 471498 597032 471554 597088
rect 471622 597032 471678 597088
rect 471250 596908 471306 596964
rect 471374 596908 471430 596964
rect 471498 596908 471554 596964
rect 471622 596908 471678 596964
rect 471250 596784 471306 596840
rect 471374 596784 471430 596840
rect 471498 596784 471554 596840
rect 471622 596784 471678 596840
rect 471250 580294 471306 580350
rect 471374 580294 471430 580350
rect 471498 580294 471554 580350
rect 471622 580294 471678 580350
rect 471250 580170 471306 580226
rect 471374 580170 471430 580226
rect 471498 580170 471554 580226
rect 471622 580170 471678 580226
rect 471250 580046 471306 580102
rect 471374 580046 471430 580102
rect 471498 580046 471554 580102
rect 471622 580046 471678 580102
rect 471250 579922 471306 579978
rect 471374 579922 471430 579978
rect 471498 579922 471554 579978
rect 471622 579922 471678 579978
rect 471250 562294 471306 562350
rect 471374 562294 471430 562350
rect 471498 562294 471554 562350
rect 471622 562294 471678 562350
rect 471250 562170 471306 562226
rect 471374 562170 471430 562226
rect 471498 562170 471554 562226
rect 471622 562170 471678 562226
rect 471250 562046 471306 562102
rect 471374 562046 471430 562102
rect 471498 562046 471554 562102
rect 471622 562046 471678 562102
rect 471250 561922 471306 561978
rect 471374 561922 471430 561978
rect 471498 561922 471554 561978
rect 471622 561922 471678 561978
rect 471250 544294 471306 544350
rect 471374 544294 471430 544350
rect 471498 544294 471554 544350
rect 471622 544294 471678 544350
rect 471250 544170 471306 544226
rect 471374 544170 471430 544226
rect 471498 544170 471554 544226
rect 471622 544170 471678 544226
rect 471250 544046 471306 544102
rect 471374 544046 471430 544102
rect 471498 544046 471554 544102
rect 471622 544046 471678 544102
rect 471250 543922 471306 543978
rect 471374 543922 471430 543978
rect 471498 543922 471554 543978
rect 471622 543922 471678 543978
rect 471250 526294 471306 526350
rect 471374 526294 471430 526350
rect 471498 526294 471554 526350
rect 471622 526294 471678 526350
rect 471250 526170 471306 526226
rect 471374 526170 471430 526226
rect 471498 526170 471554 526226
rect 471622 526170 471678 526226
rect 471250 526046 471306 526102
rect 471374 526046 471430 526102
rect 471498 526046 471554 526102
rect 471622 526046 471678 526102
rect 471250 525922 471306 525978
rect 471374 525922 471430 525978
rect 471498 525922 471554 525978
rect 471622 525922 471678 525978
rect 471250 508294 471306 508350
rect 471374 508294 471430 508350
rect 471498 508294 471554 508350
rect 471622 508294 471678 508350
rect 471250 508170 471306 508226
rect 471374 508170 471430 508226
rect 471498 508170 471554 508226
rect 471622 508170 471678 508226
rect 471250 508046 471306 508102
rect 471374 508046 471430 508102
rect 471498 508046 471554 508102
rect 471622 508046 471678 508102
rect 471250 507922 471306 507978
rect 471374 507922 471430 507978
rect 471498 507922 471554 507978
rect 471622 507922 471678 507978
rect 474970 598116 475026 598172
rect 475094 598116 475150 598172
rect 475218 598116 475274 598172
rect 475342 598116 475398 598172
rect 474970 597992 475026 598048
rect 475094 597992 475150 598048
rect 475218 597992 475274 598048
rect 475342 597992 475398 598048
rect 474970 597868 475026 597924
rect 475094 597868 475150 597924
rect 475218 597868 475274 597924
rect 475342 597868 475398 597924
rect 474970 597744 475026 597800
rect 475094 597744 475150 597800
rect 475218 597744 475274 597800
rect 475342 597744 475398 597800
rect 474970 586294 475026 586350
rect 475094 586294 475150 586350
rect 475218 586294 475274 586350
rect 475342 586294 475398 586350
rect 474970 586170 475026 586226
rect 475094 586170 475150 586226
rect 475218 586170 475274 586226
rect 475342 586170 475398 586226
rect 474970 586046 475026 586102
rect 475094 586046 475150 586102
rect 475218 586046 475274 586102
rect 475342 586046 475398 586102
rect 474970 585922 475026 585978
rect 475094 585922 475150 585978
rect 475218 585922 475274 585978
rect 475342 585922 475398 585978
rect 474970 568294 475026 568350
rect 475094 568294 475150 568350
rect 475218 568294 475274 568350
rect 475342 568294 475398 568350
rect 474970 568170 475026 568226
rect 475094 568170 475150 568226
rect 475218 568170 475274 568226
rect 475342 568170 475398 568226
rect 474970 568046 475026 568102
rect 475094 568046 475150 568102
rect 475218 568046 475274 568102
rect 475342 568046 475398 568102
rect 474970 567922 475026 567978
rect 475094 567922 475150 567978
rect 475218 567922 475274 567978
rect 475342 567922 475398 567978
rect 474970 550294 475026 550350
rect 475094 550294 475150 550350
rect 475218 550294 475274 550350
rect 475342 550294 475398 550350
rect 474970 550170 475026 550226
rect 475094 550170 475150 550226
rect 475218 550170 475274 550226
rect 475342 550170 475398 550226
rect 474970 550046 475026 550102
rect 475094 550046 475150 550102
rect 475218 550046 475274 550102
rect 475342 550046 475398 550102
rect 474970 549922 475026 549978
rect 475094 549922 475150 549978
rect 475218 549922 475274 549978
rect 475342 549922 475398 549978
rect 474970 532294 475026 532350
rect 475094 532294 475150 532350
rect 475218 532294 475274 532350
rect 475342 532294 475398 532350
rect 474970 532170 475026 532226
rect 475094 532170 475150 532226
rect 475218 532170 475274 532226
rect 475342 532170 475398 532226
rect 474970 532046 475026 532102
rect 475094 532046 475150 532102
rect 475218 532046 475274 532102
rect 475342 532046 475398 532102
rect 474970 531922 475026 531978
rect 475094 531922 475150 531978
rect 475218 531922 475274 531978
rect 475342 531922 475398 531978
rect 474970 514294 475026 514350
rect 475094 514294 475150 514350
rect 475218 514294 475274 514350
rect 475342 514294 475398 514350
rect 474970 514170 475026 514226
rect 475094 514170 475150 514226
rect 475218 514170 475274 514226
rect 475342 514170 475398 514226
rect 474970 514046 475026 514102
rect 475094 514046 475150 514102
rect 475218 514046 475274 514102
rect 475342 514046 475398 514102
rect 474970 513922 475026 513978
rect 475094 513922 475150 513978
rect 475218 513922 475274 513978
rect 475342 513922 475398 513978
rect 489250 597156 489306 597212
rect 489374 597156 489430 597212
rect 489498 597156 489554 597212
rect 489622 597156 489678 597212
rect 489250 597032 489306 597088
rect 489374 597032 489430 597088
rect 489498 597032 489554 597088
rect 489622 597032 489678 597088
rect 489250 596908 489306 596964
rect 489374 596908 489430 596964
rect 489498 596908 489554 596964
rect 489622 596908 489678 596964
rect 489250 596784 489306 596840
rect 489374 596784 489430 596840
rect 489498 596784 489554 596840
rect 489622 596784 489678 596840
rect 489250 580294 489306 580350
rect 489374 580294 489430 580350
rect 489498 580294 489554 580350
rect 489622 580294 489678 580350
rect 489250 580170 489306 580226
rect 489374 580170 489430 580226
rect 489498 580170 489554 580226
rect 489622 580170 489678 580226
rect 489250 580046 489306 580102
rect 489374 580046 489430 580102
rect 489498 580046 489554 580102
rect 489622 580046 489678 580102
rect 489250 579922 489306 579978
rect 489374 579922 489430 579978
rect 489498 579922 489554 579978
rect 489622 579922 489678 579978
rect 489250 562294 489306 562350
rect 489374 562294 489430 562350
rect 489498 562294 489554 562350
rect 489622 562294 489678 562350
rect 489250 562170 489306 562226
rect 489374 562170 489430 562226
rect 489498 562170 489554 562226
rect 489622 562170 489678 562226
rect 489250 562046 489306 562102
rect 489374 562046 489430 562102
rect 489498 562046 489554 562102
rect 489622 562046 489678 562102
rect 489250 561922 489306 561978
rect 489374 561922 489430 561978
rect 489498 561922 489554 561978
rect 489622 561922 489678 561978
rect 489250 544294 489306 544350
rect 489374 544294 489430 544350
rect 489498 544294 489554 544350
rect 489622 544294 489678 544350
rect 489250 544170 489306 544226
rect 489374 544170 489430 544226
rect 489498 544170 489554 544226
rect 489622 544170 489678 544226
rect 489250 544046 489306 544102
rect 489374 544046 489430 544102
rect 489498 544046 489554 544102
rect 489622 544046 489678 544102
rect 489250 543922 489306 543978
rect 489374 543922 489430 543978
rect 489498 543922 489554 543978
rect 489622 543922 489678 543978
rect 489250 526294 489306 526350
rect 489374 526294 489430 526350
rect 489498 526294 489554 526350
rect 489622 526294 489678 526350
rect 489250 526170 489306 526226
rect 489374 526170 489430 526226
rect 489498 526170 489554 526226
rect 489622 526170 489678 526226
rect 489250 526046 489306 526102
rect 489374 526046 489430 526102
rect 489498 526046 489554 526102
rect 489622 526046 489678 526102
rect 489250 525922 489306 525978
rect 489374 525922 489430 525978
rect 489498 525922 489554 525978
rect 489622 525922 489678 525978
rect 489250 508294 489306 508350
rect 489374 508294 489430 508350
rect 489498 508294 489554 508350
rect 489622 508294 489678 508350
rect 489250 508170 489306 508226
rect 489374 508170 489430 508226
rect 489498 508170 489554 508226
rect 489622 508170 489678 508226
rect 489250 508046 489306 508102
rect 489374 508046 489430 508102
rect 489498 508046 489554 508102
rect 489622 508046 489678 508102
rect 489250 507922 489306 507978
rect 489374 507922 489430 507978
rect 489498 507922 489554 507978
rect 489622 507922 489678 507978
rect 492970 598116 493026 598172
rect 493094 598116 493150 598172
rect 493218 598116 493274 598172
rect 493342 598116 493398 598172
rect 492970 597992 493026 598048
rect 493094 597992 493150 598048
rect 493218 597992 493274 598048
rect 493342 597992 493398 598048
rect 492970 597868 493026 597924
rect 493094 597868 493150 597924
rect 493218 597868 493274 597924
rect 493342 597868 493398 597924
rect 492970 597744 493026 597800
rect 493094 597744 493150 597800
rect 493218 597744 493274 597800
rect 493342 597744 493398 597800
rect 492970 586294 493026 586350
rect 493094 586294 493150 586350
rect 493218 586294 493274 586350
rect 493342 586294 493398 586350
rect 492970 586170 493026 586226
rect 493094 586170 493150 586226
rect 493218 586170 493274 586226
rect 493342 586170 493398 586226
rect 492970 586046 493026 586102
rect 493094 586046 493150 586102
rect 493218 586046 493274 586102
rect 493342 586046 493398 586102
rect 492970 585922 493026 585978
rect 493094 585922 493150 585978
rect 493218 585922 493274 585978
rect 493342 585922 493398 585978
rect 492970 568294 493026 568350
rect 493094 568294 493150 568350
rect 493218 568294 493274 568350
rect 493342 568294 493398 568350
rect 492970 568170 493026 568226
rect 493094 568170 493150 568226
rect 493218 568170 493274 568226
rect 493342 568170 493398 568226
rect 492970 568046 493026 568102
rect 493094 568046 493150 568102
rect 493218 568046 493274 568102
rect 493342 568046 493398 568102
rect 492970 567922 493026 567978
rect 493094 567922 493150 567978
rect 493218 567922 493274 567978
rect 493342 567922 493398 567978
rect 492970 550294 493026 550350
rect 493094 550294 493150 550350
rect 493218 550294 493274 550350
rect 493342 550294 493398 550350
rect 492970 550170 493026 550226
rect 493094 550170 493150 550226
rect 493218 550170 493274 550226
rect 493342 550170 493398 550226
rect 492970 550046 493026 550102
rect 493094 550046 493150 550102
rect 493218 550046 493274 550102
rect 493342 550046 493398 550102
rect 492970 549922 493026 549978
rect 493094 549922 493150 549978
rect 493218 549922 493274 549978
rect 493342 549922 493398 549978
rect 492970 532294 493026 532350
rect 493094 532294 493150 532350
rect 493218 532294 493274 532350
rect 493342 532294 493398 532350
rect 492970 532170 493026 532226
rect 493094 532170 493150 532226
rect 493218 532170 493274 532226
rect 493342 532170 493398 532226
rect 492970 532046 493026 532102
rect 493094 532046 493150 532102
rect 493218 532046 493274 532102
rect 493342 532046 493398 532102
rect 492970 531922 493026 531978
rect 493094 531922 493150 531978
rect 493218 531922 493274 531978
rect 493342 531922 493398 531978
rect 492970 514294 493026 514350
rect 493094 514294 493150 514350
rect 493218 514294 493274 514350
rect 493342 514294 493398 514350
rect 492970 514170 493026 514226
rect 493094 514170 493150 514226
rect 493218 514170 493274 514226
rect 493342 514170 493398 514226
rect 492970 514046 493026 514102
rect 493094 514046 493150 514102
rect 493218 514046 493274 514102
rect 493342 514046 493398 514102
rect 492970 513922 493026 513978
rect 493094 513922 493150 513978
rect 493218 513922 493274 513978
rect 493342 513922 493398 513978
rect 507250 597156 507306 597212
rect 507374 597156 507430 597212
rect 507498 597156 507554 597212
rect 507622 597156 507678 597212
rect 507250 597032 507306 597088
rect 507374 597032 507430 597088
rect 507498 597032 507554 597088
rect 507622 597032 507678 597088
rect 507250 596908 507306 596964
rect 507374 596908 507430 596964
rect 507498 596908 507554 596964
rect 507622 596908 507678 596964
rect 507250 596784 507306 596840
rect 507374 596784 507430 596840
rect 507498 596784 507554 596840
rect 507622 596784 507678 596840
rect 507250 580294 507306 580350
rect 507374 580294 507430 580350
rect 507498 580294 507554 580350
rect 507622 580294 507678 580350
rect 507250 580170 507306 580226
rect 507374 580170 507430 580226
rect 507498 580170 507554 580226
rect 507622 580170 507678 580226
rect 507250 580046 507306 580102
rect 507374 580046 507430 580102
rect 507498 580046 507554 580102
rect 507622 580046 507678 580102
rect 507250 579922 507306 579978
rect 507374 579922 507430 579978
rect 507498 579922 507554 579978
rect 507622 579922 507678 579978
rect 507250 562294 507306 562350
rect 507374 562294 507430 562350
rect 507498 562294 507554 562350
rect 507622 562294 507678 562350
rect 507250 562170 507306 562226
rect 507374 562170 507430 562226
rect 507498 562170 507554 562226
rect 507622 562170 507678 562226
rect 507250 562046 507306 562102
rect 507374 562046 507430 562102
rect 507498 562046 507554 562102
rect 507622 562046 507678 562102
rect 507250 561922 507306 561978
rect 507374 561922 507430 561978
rect 507498 561922 507554 561978
rect 507622 561922 507678 561978
rect 507250 544294 507306 544350
rect 507374 544294 507430 544350
rect 507498 544294 507554 544350
rect 507622 544294 507678 544350
rect 507250 544170 507306 544226
rect 507374 544170 507430 544226
rect 507498 544170 507554 544226
rect 507622 544170 507678 544226
rect 507250 544046 507306 544102
rect 507374 544046 507430 544102
rect 507498 544046 507554 544102
rect 507622 544046 507678 544102
rect 507250 543922 507306 543978
rect 507374 543922 507430 543978
rect 507498 543922 507554 543978
rect 507622 543922 507678 543978
rect 507250 526294 507306 526350
rect 507374 526294 507430 526350
rect 507498 526294 507554 526350
rect 507622 526294 507678 526350
rect 507250 526170 507306 526226
rect 507374 526170 507430 526226
rect 507498 526170 507554 526226
rect 507622 526170 507678 526226
rect 507250 526046 507306 526102
rect 507374 526046 507430 526102
rect 507498 526046 507554 526102
rect 507622 526046 507678 526102
rect 507250 525922 507306 525978
rect 507374 525922 507430 525978
rect 507498 525922 507554 525978
rect 507622 525922 507678 525978
rect 507250 508294 507306 508350
rect 507374 508294 507430 508350
rect 507498 508294 507554 508350
rect 507622 508294 507678 508350
rect 507250 508170 507306 508226
rect 507374 508170 507430 508226
rect 507498 508170 507554 508226
rect 507622 508170 507678 508226
rect 507250 508046 507306 508102
rect 507374 508046 507430 508102
rect 507498 508046 507554 508102
rect 507622 508046 507678 508102
rect 507250 507922 507306 507978
rect 507374 507922 507430 507978
rect 507498 507922 507554 507978
rect 507622 507922 507678 507978
rect 219878 496277 219934 496333
rect 220002 496277 220058 496333
rect 219878 496153 219934 496209
rect 220002 496153 220058 496209
rect 219878 496029 219934 496085
rect 220002 496029 220058 496085
rect 219878 495905 219934 495961
rect 220002 495905 220058 495961
rect 250598 496277 250654 496333
rect 250722 496277 250778 496333
rect 250598 496153 250654 496209
rect 250722 496153 250778 496209
rect 250598 496029 250654 496085
rect 250722 496029 250778 496085
rect 250598 495905 250654 495961
rect 250722 495905 250778 495961
rect 281318 496277 281374 496333
rect 281442 496277 281498 496333
rect 281318 496153 281374 496209
rect 281442 496153 281498 496209
rect 281318 496029 281374 496085
rect 281442 496029 281498 496085
rect 281318 495905 281374 495961
rect 281442 495905 281498 495961
rect 312038 496277 312094 496333
rect 312162 496277 312218 496333
rect 312038 496153 312094 496209
rect 312162 496153 312218 496209
rect 312038 496029 312094 496085
rect 312162 496029 312218 496085
rect 312038 495905 312094 495961
rect 312162 495905 312218 495961
rect 342758 496277 342814 496333
rect 342882 496277 342938 496333
rect 342758 496153 342814 496209
rect 342882 496153 342938 496209
rect 342758 496029 342814 496085
rect 342882 496029 342938 496085
rect 342758 495905 342814 495961
rect 342882 495905 342938 495961
rect 373478 496277 373534 496333
rect 373602 496277 373658 496333
rect 373478 496153 373534 496209
rect 373602 496153 373658 496209
rect 373478 496029 373534 496085
rect 373602 496029 373658 496085
rect 373478 495905 373534 495961
rect 373602 495905 373658 495961
rect 404198 496277 404254 496333
rect 404322 496277 404378 496333
rect 404198 496153 404254 496209
rect 404322 496153 404378 496209
rect 404198 496029 404254 496085
rect 404322 496029 404378 496085
rect 404198 495905 404254 495961
rect 404322 495905 404378 495961
rect 434918 496277 434974 496333
rect 435042 496277 435098 496333
rect 434918 496153 434974 496209
rect 435042 496153 435098 496209
rect 434918 496029 434974 496085
rect 435042 496029 435098 496085
rect 434918 495905 434974 495961
rect 435042 495905 435098 495961
rect 465638 496277 465694 496333
rect 465762 496277 465818 496333
rect 465638 496153 465694 496209
rect 465762 496153 465818 496209
rect 465638 496029 465694 496085
rect 465762 496029 465818 496085
rect 465638 495905 465694 495961
rect 465762 495905 465818 495961
rect 496358 496277 496414 496333
rect 496482 496277 496538 496333
rect 496358 496153 496414 496209
rect 496482 496153 496538 496209
rect 496358 496029 496414 496085
rect 496482 496029 496538 496085
rect 496358 495905 496414 495961
rect 496482 495905 496538 495961
rect 201250 490294 201306 490350
rect 201374 490294 201430 490350
rect 201498 490294 201554 490350
rect 201622 490294 201678 490350
rect 201250 490170 201306 490226
rect 201374 490170 201430 490226
rect 201498 490170 201554 490226
rect 201622 490170 201678 490226
rect 201250 490046 201306 490102
rect 201374 490046 201430 490102
rect 201498 490046 201554 490102
rect 201622 490046 201678 490102
rect 201250 489922 201306 489978
rect 201374 489922 201430 489978
rect 201498 489922 201554 489978
rect 201622 489922 201678 489978
rect 204518 490294 204574 490350
rect 204642 490294 204698 490350
rect 204518 490170 204574 490226
rect 204642 490170 204698 490226
rect 204518 490046 204574 490102
rect 204642 490046 204698 490102
rect 204518 489922 204574 489978
rect 204642 489922 204698 489978
rect 235238 490294 235294 490350
rect 235362 490294 235418 490350
rect 235238 490170 235294 490226
rect 235362 490170 235418 490226
rect 235238 490046 235294 490102
rect 235362 490046 235418 490102
rect 235238 489922 235294 489978
rect 235362 489922 235418 489978
rect 265958 490294 266014 490350
rect 266082 490294 266138 490350
rect 265958 490170 266014 490226
rect 266082 490170 266138 490226
rect 265958 490046 266014 490102
rect 266082 490046 266138 490102
rect 265958 489922 266014 489978
rect 266082 489922 266138 489978
rect 296678 490294 296734 490350
rect 296802 490294 296858 490350
rect 296678 490170 296734 490226
rect 296802 490170 296858 490226
rect 296678 490046 296734 490102
rect 296802 490046 296858 490102
rect 296678 489922 296734 489978
rect 296802 489922 296858 489978
rect 327398 490294 327454 490350
rect 327522 490294 327578 490350
rect 327398 490170 327454 490226
rect 327522 490170 327578 490226
rect 327398 490046 327454 490102
rect 327522 490046 327578 490102
rect 327398 489922 327454 489978
rect 327522 489922 327578 489978
rect 358118 490294 358174 490350
rect 358242 490294 358298 490350
rect 358118 490170 358174 490226
rect 358242 490170 358298 490226
rect 358118 490046 358174 490102
rect 358242 490046 358298 490102
rect 358118 489922 358174 489978
rect 358242 489922 358298 489978
rect 388838 490294 388894 490350
rect 388962 490294 389018 490350
rect 388838 490170 388894 490226
rect 388962 490170 389018 490226
rect 388838 490046 388894 490102
rect 388962 490046 389018 490102
rect 388838 489922 388894 489978
rect 388962 489922 389018 489978
rect 419558 490294 419614 490350
rect 419682 490294 419738 490350
rect 419558 490170 419614 490226
rect 419682 490170 419738 490226
rect 419558 490046 419614 490102
rect 419682 490046 419738 490102
rect 419558 489922 419614 489978
rect 419682 489922 419738 489978
rect 450278 490294 450334 490350
rect 450402 490294 450458 490350
rect 450278 490170 450334 490226
rect 450402 490170 450458 490226
rect 450278 490046 450334 490102
rect 450402 490046 450458 490102
rect 450278 489922 450334 489978
rect 450402 489922 450458 489978
rect 480998 490294 481054 490350
rect 481122 490294 481178 490350
rect 480998 490170 481054 490226
rect 481122 490170 481178 490226
rect 480998 490046 481054 490102
rect 481122 490046 481178 490102
rect 480998 489922 481054 489978
rect 481122 489922 481178 489978
rect 507250 490294 507306 490350
rect 507374 490294 507430 490350
rect 507498 490294 507554 490350
rect 507622 490294 507678 490350
rect 507250 490170 507306 490226
rect 507374 490170 507430 490226
rect 507498 490170 507554 490226
rect 507622 490170 507678 490226
rect 507250 490046 507306 490102
rect 507374 490046 507430 490102
rect 507498 490046 507554 490102
rect 507622 490046 507678 490102
rect 507250 489922 507306 489978
rect 507374 489922 507430 489978
rect 507498 489922 507554 489978
rect 507622 489922 507678 489978
rect 219878 478294 219934 478350
rect 220002 478294 220058 478350
rect 219878 478170 219934 478226
rect 220002 478170 220058 478226
rect 219878 478046 219934 478102
rect 220002 478046 220058 478102
rect 219878 477922 219934 477978
rect 220002 477922 220058 477978
rect 250598 478294 250654 478350
rect 250722 478294 250778 478350
rect 250598 478170 250654 478226
rect 250722 478170 250778 478226
rect 250598 478046 250654 478102
rect 250722 478046 250778 478102
rect 250598 477922 250654 477978
rect 250722 477922 250778 477978
rect 281318 478294 281374 478350
rect 281442 478294 281498 478350
rect 281318 478170 281374 478226
rect 281442 478170 281498 478226
rect 281318 478046 281374 478102
rect 281442 478046 281498 478102
rect 281318 477922 281374 477978
rect 281442 477922 281498 477978
rect 312038 478294 312094 478350
rect 312162 478294 312218 478350
rect 312038 478170 312094 478226
rect 312162 478170 312218 478226
rect 312038 478046 312094 478102
rect 312162 478046 312218 478102
rect 312038 477922 312094 477978
rect 312162 477922 312218 477978
rect 342758 478294 342814 478350
rect 342882 478294 342938 478350
rect 342758 478170 342814 478226
rect 342882 478170 342938 478226
rect 342758 478046 342814 478102
rect 342882 478046 342938 478102
rect 342758 477922 342814 477978
rect 342882 477922 342938 477978
rect 373478 478294 373534 478350
rect 373602 478294 373658 478350
rect 373478 478170 373534 478226
rect 373602 478170 373658 478226
rect 373478 478046 373534 478102
rect 373602 478046 373658 478102
rect 373478 477922 373534 477978
rect 373602 477922 373658 477978
rect 404198 478294 404254 478350
rect 404322 478294 404378 478350
rect 404198 478170 404254 478226
rect 404322 478170 404378 478226
rect 404198 478046 404254 478102
rect 404322 478046 404378 478102
rect 404198 477922 404254 477978
rect 404322 477922 404378 477978
rect 434918 478294 434974 478350
rect 435042 478294 435098 478350
rect 434918 478170 434974 478226
rect 435042 478170 435098 478226
rect 434918 478046 434974 478102
rect 435042 478046 435098 478102
rect 434918 477922 434974 477978
rect 435042 477922 435098 477978
rect 465638 478294 465694 478350
rect 465762 478294 465818 478350
rect 465638 478170 465694 478226
rect 465762 478170 465818 478226
rect 465638 478046 465694 478102
rect 465762 478046 465818 478102
rect 465638 477922 465694 477978
rect 465762 477922 465818 477978
rect 496358 478294 496414 478350
rect 496482 478294 496538 478350
rect 496358 478170 496414 478226
rect 496482 478170 496538 478226
rect 496358 478046 496414 478102
rect 496482 478046 496538 478102
rect 496358 477922 496414 477978
rect 496482 477922 496538 477978
rect 201250 472294 201306 472350
rect 201374 472294 201430 472350
rect 201498 472294 201554 472350
rect 201622 472294 201678 472350
rect 201250 472170 201306 472226
rect 201374 472170 201430 472226
rect 201498 472170 201554 472226
rect 201622 472170 201678 472226
rect 201250 472046 201306 472102
rect 201374 472046 201430 472102
rect 201498 472046 201554 472102
rect 201622 472046 201678 472102
rect 201250 471922 201306 471978
rect 201374 471922 201430 471978
rect 201498 471922 201554 471978
rect 201622 471922 201678 471978
rect 204518 472294 204574 472350
rect 204642 472294 204698 472350
rect 204518 472170 204574 472226
rect 204642 472170 204698 472226
rect 204518 472046 204574 472102
rect 204642 472046 204698 472102
rect 204518 471922 204574 471978
rect 204642 471922 204698 471978
rect 235238 472294 235294 472350
rect 235362 472294 235418 472350
rect 235238 472170 235294 472226
rect 235362 472170 235418 472226
rect 235238 472046 235294 472102
rect 235362 472046 235418 472102
rect 235238 471922 235294 471978
rect 235362 471922 235418 471978
rect 265958 472294 266014 472350
rect 266082 472294 266138 472350
rect 265958 472170 266014 472226
rect 266082 472170 266138 472226
rect 265958 472046 266014 472102
rect 266082 472046 266138 472102
rect 265958 471922 266014 471978
rect 266082 471922 266138 471978
rect 296678 472294 296734 472350
rect 296802 472294 296858 472350
rect 296678 472170 296734 472226
rect 296802 472170 296858 472226
rect 296678 472046 296734 472102
rect 296802 472046 296858 472102
rect 296678 471922 296734 471978
rect 296802 471922 296858 471978
rect 327398 472294 327454 472350
rect 327522 472294 327578 472350
rect 327398 472170 327454 472226
rect 327522 472170 327578 472226
rect 327398 472046 327454 472102
rect 327522 472046 327578 472102
rect 327398 471922 327454 471978
rect 327522 471922 327578 471978
rect 358118 472294 358174 472350
rect 358242 472294 358298 472350
rect 358118 472170 358174 472226
rect 358242 472170 358298 472226
rect 358118 472046 358174 472102
rect 358242 472046 358298 472102
rect 358118 471922 358174 471978
rect 358242 471922 358298 471978
rect 388838 472294 388894 472350
rect 388962 472294 389018 472350
rect 388838 472170 388894 472226
rect 388962 472170 389018 472226
rect 388838 472046 388894 472102
rect 388962 472046 389018 472102
rect 388838 471922 388894 471978
rect 388962 471922 389018 471978
rect 419558 472294 419614 472350
rect 419682 472294 419738 472350
rect 419558 472170 419614 472226
rect 419682 472170 419738 472226
rect 419558 472046 419614 472102
rect 419682 472046 419738 472102
rect 419558 471922 419614 471978
rect 419682 471922 419738 471978
rect 450278 472294 450334 472350
rect 450402 472294 450458 472350
rect 450278 472170 450334 472226
rect 450402 472170 450458 472226
rect 450278 472046 450334 472102
rect 450402 472046 450458 472102
rect 450278 471922 450334 471978
rect 450402 471922 450458 471978
rect 480998 472294 481054 472350
rect 481122 472294 481178 472350
rect 480998 472170 481054 472226
rect 481122 472170 481178 472226
rect 480998 472046 481054 472102
rect 481122 472046 481178 472102
rect 480998 471922 481054 471978
rect 481122 471922 481178 471978
rect 507250 472294 507306 472350
rect 507374 472294 507430 472350
rect 507498 472294 507554 472350
rect 507622 472294 507678 472350
rect 507250 472170 507306 472226
rect 507374 472170 507430 472226
rect 507498 472170 507554 472226
rect 507622 472170 507678 472226
rect 507250 472046 507306 472102
rect 507374 472046 507430 472102
rect 507498 472046 507554 472102
rect 507622 472046 507678 472102
rect 507250 471922 507306 471978
rect 507374 471922 507430 471978
rect 507498 471922 507554 471978
rect 507622 471922 507678 471978
rect 219878 460294 219934 460350
rect 220002 460294 220058 460350
rect 219878 460170 219934 460226
rect 220002 460170 220058 460226
rect 219878 460046 219934 460102
rect 220002 460046 220058 460102
rect 219878 459922 219934 459978
rect 220002 459922 220058 459978
rect 250598 460294 250654 460350
rect 250722 460294 250778 460350
rect 250598 460170 250654 460226
rect 250722 460170 250778 460226
rect 250598 460046 250654 460102
rect 250722 460046 250778 460102
rect 250598 459922 250654 459978
rect 250722 459922 250778 459978
rect 281318 460294 281374 460350
rect 281442 460294 281498 460350
rect 281318 460170 281374 460226
rect 281442 460170 281498 460226
rect 281318 460046 281374 460102
rect 281442 460046 281498 460102
rect 281318 459922 281374 459978
rect 281442 459922 281498 459978
rect 312038 460294 312094 460350
rect 312162 460294 312218 460350
rect 312038 460170 312094 460226
rect 312162 460170 312218 460226
rect 312038 460046 312094 460102
rect 312162 460046 312218 460102
rect 312038 459922 312094 459978
rect 312162 459922 312218 459978
rect 342758 460294 342814 460350
rect 342882 460294 342938 460350
rect 342758 460170 342814 460226
rect 342882 460170 342938 460226
rect 342758 460046 342814 460102
rect 342882 460046 342938 460102
rect 342758 459922 342814 459978
rect 342882 459922 342938 459978
rect 373478 460294 373534 460350
rect 373602 460294 373658 460350
rect 373478 460170 373534 460226
rect 373602 460170 373658 460226
rect 373478 460046 373534 460102
rect 373602 460046 373658 460102
rect 373478 459922 373534 459978
rect 373602 459922 373658 459978
rect 404198 460294 404254 460350
rect 404322 460294 404378 460350
rect 404198 460170 404254 460226
rect 404322 460170 404378 460226
rect 404198 460046 404254 460102
rect 404322 460046 404378 460102
rect 404198 459922 404254 459978
rect 404322 459922 404378 459978
rect 434918 460294 434974 460350
rect 435042 460294 435098 460350
rect 434918 460170 434974 460226
rect 435042 460170 435098 460226
rect 434918 460046 434974 460102
rect 435042 460046 435098 460102
rect 434918 459922 434974 459978
rect 435042 459922 435098 459978
rect 465638 460294 465694 460350
rect 465762 460294 465818 460350
rect 465638 460170 465694 460226
rect 465762 460170 465818 460226
rect 465638 460046 465694 460102
rect 465762 460046 465818 460102
rect 465638 459922 465694 459978
rect 465762 459922 465818 459978
rect 496358 460294 496414 460350
rect 496482 460294 496538 460350
rect 496358 460170 496414 460226
rect 496482 460170 496538 460226
rect 496358 460046 496414 460102
rect 496482 460046 496538 460102
rect 496358 459922 496414 459978
rect 496482 459922 496538 459978
rect 201250 454294 201306 454350
rect 201374 454294 201430 454350
rect 201498 454294 201554 454350
rect 201622 454294 201678 454350
rect 201250 454170 201306 454226
rect 201374 454170 201430 454226
rect 201498 454170 201554 454226
rect 201622 454170 201678 454226
rect 201250 454046 201306 454102
rect 201374 454046 201430 454102
rect 201498 454046 201554 454102
rect 201622 454046 201678 454102
rect 201250 453922 201306 453978
rect 201374 453922 201430 453978
rect 201498 453922 201554 453978
rect 201622 453922 201678 453978
rect 204518 454294 204574 454350
rect 204642 454294 204698 454350
rect 204518 454170 204574 454226
rect 204642 454170 204698 454226
rect 204518 454046 204574 454102
rect 204642 454046 204698 454102
rect 204518 453922 204574 453978
rect 204642 453922 204698 453978
rect 235238 454294 235294 454350
rect 235362 454294 235418 454350
rect 235238 454170 235294 454226
rect 235362 454170 235418 454226
rect 235238 454046 235294 454102
rect 235362 454046 235418 454102
rect 235238 453922 235294 453978
rect 235362 453922 235418 453978
rect 265958 454294 266014 454350
rect 266082 454294 266138 454350
rect 265958 454170 266014 454226
rect 266082 454170 266138 454226
rect 265958 454046 266014 454102
rect 266082 454046 266138 454102
rect 265958 453922 266014 453978
rect 266082 453922 266138 453978
rect 296678 454294 296734 454350
rect 296802 454294 296858 454350
rect 296678 454170 296734 454226
rect 296802 454170 296858 454226
rect 296678 454046 296734 454102
rect 296802 454046 296858 454102
rect 296678 453922 296734 453978
rect 296802 453922 296858 453978
rect 327398 454294 327454 454350
rect 327522 454294 327578 454350
rect 327398 454170 327454 454226
rect 327522 454170 327578 454226
rect 327398 454046 327454 454102
rect 327522 454046 327578 454102
rect 327398 453922 327454 453978
rect 327522 453922 327578 453978
rect 358118 454294 358174 454350
rect 358242 454294 358298 454350
rect 358118 454170 358174 454226
rect 358242 454170 358298 454226
rect 358118 454046 358174 454102
rect 358242 454046 358298 454102
rect 358118 453922 358174 453978
rect 358242 453922 358298 453978
rect 388838 454294 388894 454350
rect 388962 454294 389018 454350
rect 388838 454170 388894 454226
rect 388962 454170 389018 454226
rect 388838 454046 388894 454102
rect 388962 454046 389018 454102
rect 388838 453922 388894 453978
rect 388962 453922 389018 453978
rect 419558 454294 419614 454350
rect 419682 454294 419738 454350
rect 419558 454170 419614 454226
rect 419682 454170 419738 454226
rect 419558 454046 419614 454102
rect 419682 454046 419738 454102
rect 419558 453922 419614 453978
rect 419682 453922 419738 453978
rect 450278 454294 450334 454350
rect 450402 454294 450458 454350
rect 450278 454170 450334 454226
rect 450402 454170 450458 454226
rect 450278 454046 450334 454102
rect 450402 454046 450458 454102
rect 450278 453922 450334 453978
rect 450402 453922 450458 453978
rect 480998 454294 481054 454350
rect 481122 454294 481178 454350
rect 480998 454170 481054 454226
rect 481122 454170 481178 454226
rect 480998 454046 481054 454102
rect 481122 454046 481178 454102
rect 480998 453922 481054 453978
rect 481122 453922 481178 453978
rect 507250 454294 507306 454350
rect 507374 454294 507430 454350
rect 507498 454294 507554 454350
rect 507622 454294 507678 454350
rect 507250 454170 507306 454226
rect 507374 454170 507430 454226
rect 507498 454170 507554 454226
rect 507622 454170 507678 454226
rect 507250 454046 507306 454102
rect 507374 454046 507430 454102
rect 507498 454046 507554 454102
rect 507622 454046 507678 454102
rect 507250 453922 507306 453978
rect 507374 453922 507430 453978
rect 507498 453922 507554 453978
rect 507622 453922 507678 453978
rect 219878 442294 219934 442350
rect 220002 442294 220058 442350
rect 219878 442170 219934 442226
rect 220002 442170 220058 442226
rect 219878 442046 219934 442102
rect 220002 442046 220058 442102
rect 219878 441922 219934 441978
rect 220002 441922 220058 441978
rect 250598 442294 250654 442350
rect 250722 442294 250778 442350
rect 250598 442170 250654 442226
rect 250722 442170 250778 442226
rect 250598 442046 250654 442102
rect 250722 442046 250778 442102
rect 250598 441922 250654 441978
rect 250722 441922 250778 441978
rect 281318 442294 281374 442350
rect 281442 442294 281498 442350
rect 281318 442170 281374 442226
rect 281442 442170 281498 442226
rect 281318 442046 281374 442102
rect 281442 442046 281498 442102
rect 281318 441922 281374 441978
rect 281442 441922 281498 441978
rect 312038 442294 312094 442350
rect 312162 442294 312218 442350
rect 312038 442170 312094 442226
rect 312162 442170 312218 442226
rect 312038 442046 312094 442102
rect 312162 442046 312218 442102
rect 312038 441922 312094 441978
rect 312162 441922 312218 441978
rect 342758 442294 342814 442350
rect 342882 442294 342938 442350
rect 342758 442170 342814 442226
rect 342882 442170 342938 442226
rect 342758 442046 342814 442102
rect 342882 442046 342938 442102
rect 342758 441922 342814 441978
rect 342882 441922 342938 441978
rect 373478 442294 373534 442350
rect 373602 442294 373658 442350
rect 373478 442170 373534 442226
rect 373602 442170 373658 442226
rect 373478 442046 373534 442102
rect 373602 442046 373658 442102
rect 373478 441922 373534 441978
rect 373602 441922 373658 441978
rect 404198 442294 404254 442350
rect 404322 442294 404378 442350
rect 404198 442170 404254 442226
rect 404322 442170 404378 442226
rect 404198 442046 404254 442102
rect 404322 442046 404378 442102
rect 404198 441922 404254 441978
rect 404322 441922 404378 441978
rect 434918 442294 434974 442350
rect 435042 442294 435098 442350
rect 434918 442170 434974 442226
rect 435042 442170 435098 442226
rect 434918 442046 434974 442102
rect 435042 442046 435098 442102
rect 434918 441922 434974 441978
rect 435042 441922 435098 441978
rect 465638 442294 465694 442350
rect 465762 442294 465818 442350
rect 465638 442170 465694 442226
rect 465762 442170 465818 442226
rect 465638 442046 465694 442102
rect 465762 442046 465818 442102
rect 465638 441922 465694 441978
rect 465762 441922 465818 441978
rect 496358 442294 496414 442350
rect 496482 442294 496538 442350
rect 496358 442170 496414 442226
rect 496482 442170 496538 442226
rect 496358 442046 496414 442102
rect 496482 442046 496538 442102
rect 496358 441922 496414 441978
rect 496482 441922 496538 441978
rect 201250 436294 201306 436350
rect 201374 436294 201430 436350
rect 201498 436294 201554 436350
rect 201622 436294 201678 436350
rect 201250 436170 201306 436226
rect 201374 436170 201430 436226
rect 201498 436170 201554 436226
rect 201622 436170 201678 436226
rect 201250 436046 201306 436102
rect 201374 436046 201430 436102
rect 201498 436046 201554 436102
rect 201622 436046 201678 436102
rect 201250 435922 201306 435978
rect 201374 435922 201430 435978
rect 201498 435922 201554 435978
rect 201622 435922 201678 435978
rect 204518 436294 204574 436350
rect 204642 436294 204698 436350
rect 204518 436170 204574 436226
rect 204642 436170 204698 436226
rect 204518 436046 204574 436102
rect 204642 436046 204698 436102
rect 204518 435922 204574 435978
rect 204642 435922 204698 435978
rect 235238 436294 235294 436350
rect 235362 436294 235418 436350
rect 235238 436170 235294 436226
rect 235362 436170 235418 436226
rect 235238 436046 235294 436102
rect 235362 436046 235418 436102
rect 235238 435922 235294 435978
rect 235362 435922 235418 435978
rect 265958 436294 266014 436350
rect 266082 436294 266138 436350
rect 265958 436170 266014 436226
rect 266082 436170 266138 436226
rect 265958 436046 266014 436102
rect 266082 436046 266138 436102
rect 265958 435922 266014 435978
rect 266082 435922 266138 435978
rect 296678 436294 296734 436350
rect 296802 436294 296858 436350
rect 296678 436170 296734 436226
rect 296802 436170 296858 436226
rect 296678 436046 296734 436102
rect 296802 436046 296858 436102
rect 296678 435922 296734 435978
rect 296802 435922 296858 435978
rect 327398 436294 327454 436350
rect 327522 436294 327578 436350
rect 327398 436170 327454 436226
rect 327522 436170 327578 436226
rect 327398 436046 327454 436102
rect 327522 436046 327578 436102
rect 327398 435922 327454 435978
rect 327522 435922 327578 435978
rect 358118 436294 358174 436350
rect 358242 436294 358298 436350
rect 358118 436170 358174 436226
rect 358242 436170 358298 436226
rect 358118 436046 358174 436102
rect 358242 436046 358298 436102
rect 358118 435922 358174 435978
rect 358242 435922 358298 435978
rect 388838 436294 388894 436350
rect 388962 436294 389018 436350
rect 388838 436170 388894 436226
rect 388962 436170 389018 436226
rect 388838 436046 388894 436102
rect 388962 436046 389018 436102
rect 388838 435922 388894 435978
rect 388962 435922 389018 435978
rect 419558 436294 419614 436350
rect 419682 436294 419738 436350
rect 419558 436170 419614 436226
rect 419682 436170 419738 436226
rect 419558 436046 419614 436102
rect 419682 436046 419738 436102
rect 419558 435922 419614 435978
rect 419682 435922 419738 435978
rect 450278 436294 450334 436350
rect 450402 436294 450458 436350
rect 450278 436170 450334 436226
rect 450402 436170 450458 436226
rect 450278 436046 450334 436102
rect 450402 436046 450458 436102
rect 450278 435922 450334 435978
rect 450402 435922 450458 435978
rect 480998 436294 481054 436350
rect 481122 436294 481178 436350
rect 480998 436170 481054 436226
rect 481122 436170 481178 436226
rect 480998 436046 481054 436102
rect 481122 436046 481178 436102
rect 480998 435922 481054 435978
rect 481122 435922 481178 435978
rect 507250 436294 507306 436350
rect 507374 436294 507430 436350
rect 507498 436294 507554 436350
rect 507622 436294 507678 436350
rect 507250 436170 507306 436226
rect 507374 436170 507430 436226
rect 507498 436170 507554 436226
rect 507622 436170 507678 436226
rect 507250 436046 507306 436102
rect 507374 436046 507430 436102
rect 507498 436046 507554 436102
rect 507622 436046 507678 436102
rect 507250 435922 507306 435978
rect 507374 435922 507430 435978
rect 507498 435922 507554 435978
rect 507622 435922 507678 435978
rect 219878 424294 219934 424350
rect 220002 424294 220058 424350
rect 219878 424170 219934 424226
rect 220002 424170 220058 424226
rect 219878 424046 219934 424102
rect 220002 424046 220058 424102
rect 219878 423922 219934 423978
rect 220002 423922 220058 423978
rect 250598 424294 250654 424350
rect 250722 424294 250778 424350
rect 250598 424170 250654 424226
rect 250722 424170 250778 424226
rect 250598 424046 250654 424102
rect 250722 424046 250778 424102
rect 250598 423922 250654 423978
rect 250722 423922 250778 423978
rect 281318 424294 281374 424350
rect 281442 424294 281498 424350
rect 281318 424170 281374 424226
rect 281442 424170 281498 424226
rect 281318 424046 281374 424102
rect 281442 424046 281498 424102
rect 281318 423922 281374 423978
rect 281442 423922 281498 423978
rect 312038 424294 312094 424350
rect 312162 424294 312218 424350
rect 312038 424170 312094 424226
rect 312162 424170 312218 424226
rect 312038 424046 312094 424102
rect 312162 424046 312218 424102
rect 312038 423922 312094 423978
rect 312162 423922 312218 423978
rect 342758 424294 342814 424350
rect 342882 424294 342938 424350
rect 342758 424170 342814 424226
rect 342882 424170 342938 424226
rect 342758 424046 342814 424102
rect 342882 424046 342938 424102
rect 342758 423922 342814 423978
rect 342882 423922 342938 423978
rect 373478 424294 373534 424350
rect 373602 424294 373658 424350
rect 373478 424170 373534 424226
rect 373602 424170 373658 424226
rect 373478 424046 373534 424102
rect 373602 424046 373658 424102
rect 373478 423922 373534 423978
rect 373602 423922 373658 423978
rect 404198 424294 404254 424350
rect 404322 424294 404378 424350
rect 404198 424170 404254 424226
rect 404322 424170 404378 424226
rect 404198 424046 404254 424102
rect 404322 424046 404378 424102
rect 404198 423922 404254 423978
rect 404322 423922 404378 423978
rect 434918 424294 434974 424350
rect 435042 424294 435098 424350
rect 434918 424170 434974 424226
rect 435042 424170 435098 424226
rect 434918 424046 434974 424102
rect 435042 424046 435098 424102
rect 434918 423922 434974 423978
rect 435042 423922 435098 423978
rect 465638 424294 465694 424350
rect 465762 424294 465818 424350
rect 465638 424170 465694 424226
rect 465762 424170 465818 424226
rect 465638 424046 465694 424102
rect 465762 424046 465818 424102
rect 465638 423922 465694 423978
rect 465762 423922 465818 423978
rect 496358 424294 496414 424350
rect 496482 424294 496538 424350
rect 496358 424170 496414 424226
rect 496482 424170 496538 424226
rect 496358 424046 496414 424102
rect 496482 424046 496538 424102
rect 496358 423922 496414 423978
rect 496482 423922 496538 423978
rect 201250 418294 201306 418350
rect 201374 418294 201430 418350
rect 201498 418294 201554 418350
rect 201622 418294 201678 418350
rect 201250 418170 201306 418226
rect 201374 418170 201430 418226
rect 201498 418170 201554 418226
rect 201622 418170 201678 418226
rect 201250 418046 201306 418102
rect 201374 418046 201430 418102
rect 201498 418046 201554 418102
rect 201622 418046 201678 418102
rect 201250 417922 201306 417978
rect 201374 417922 201430 417978
rect 201498 417922 201554 417978
rect 201622 417922 201678 417978
rect 204518 418294 204574 418350
rect 204642 418294 204698 418350
rect 204518 418170 204574 418226
rect 204642 418170 204698 418226
rect 204518 418046 204574 418102
rect 204642 418046 204698 418102
rect 204518 417922 204574 417978
rect 204642 417922 204698 417978
rect 235238 418294 235294 418350
rect 235362 418294 235418 418350
rect 235238 418170 235294 418226
rect 235362 418170 235418 418226
rect 235238 418046 235294 418102
rect 235362 418046 235418 418102
rect 235238 417922 235294 417978
rect 235362 417922 235418 417978
rect 265958 418294 266014 418350
rect 266082 418294 266138 418350
rect 265958 418170 266014 418226
rect 266082 418170 266138 418226
rect 265958 418046 266014 418102
rect 266082 418046 266138 418102
rect 265958 417922 266014 417978
rect 266082 417922 266138 417978
rect 296678 418294 296734 418350
rect 296802 418294 296858 418350
rect 296678 418170 296734 418226
rect 296802 418170 296858 418226
rect 296678 418046 296734 418102
rect 296802 418046 296858 418102
rect 296678 417922 296734 417978
rect 296802 417922 296858 417978
rect 327398 418294 327454 418350
rect 327522 418294 327578 418350
rect 327398 418170 327454 418226
rect 327522 418170 327578 418226
rect 327398 418046 327454 418102
rect 327522 418046 327578 418102
rect 327398 417922 327454 417978
rect 327522 417922 327578 417978
rect 358118 418294 358174 418350
rect 358242 418294 358298 418350
rect 358118 418170 358174 418226
rect 358242 418170 358298 418226
rect 358118 418046 358174 418102
rect 358242 418046 358298 418102
rect 358118 417922 358174 417978
rect 358242 417922 358298 417978
rect 388838 418294 388894 418350
rect 388962 418294 389018 418350
rect 388838 418170 388894 418226
rect 388962 418170 389018 418226
rect 388838 418046 388894 418102
rect 388962 418046 389018 418102
rect 388838 417922 388894 417978
rect 388962 417922 389018 417978
rect 419558 418294 419614 418350
rect 419682 418294 419738 418350
rect 419558 418170 419614 418226
rect 419682 418170 419738 418226
rect 419558 418046 419614 418102
rect 419682 418046 419738 418102
rect 419558 417922 419614 417978
rect 419682 417922 419738 417978
rect 450278 418294 450334 418350
rect 450402 418294 450458 418350
rect 450278 418170 450334 418226
rect 450402 418170 450458 418226
rect 450278 418046 450334 418102
rect 450402 418046 450458 418102
rect 450278 417922 450334 417978
rect 450402 417922 450458 417978
rect 480998 418294 481054 418350
rect 481122 418294 481178 418350
rect 480998 418170 481054 418226
rect 481122 418170 481178 418226
rect 480998 418046 481054 418102
rect 481122 418046 481178 418102
rect 480998 417922 481054 417978
rect 481122 417922 481178 417978
rect 507250 418294 507306 418350
rect 507374 418294 507430 418350
rect 507498 418294 507554 418350
rect 507622 418294 507678 418350
rect 507250 418170 507306 418226
rect 507374 418170 507430 418226
rect 507498 418170 507554 418226
rect 507622 418170 507678 418226
rect 507250 418046 507306 418102
rect 507374 418046 507430 418102
rect 507498 418046 507554 418102
rect 507622 418046 507678 418102
rect 507250 417922 507306 417978
rect 507374 417922 507430 417978
rect 507498 417922 507554 417978
rect 507622 417922 507678 417978
rect 219878 406294 219934 406350
rect 220002 406294 220058 406350
rect 219878 406170 219934 406226
rect 220002 406170 220058 406226
rect 219878 406046 219934 406102
rect 220002 406046 220058 406102
rect 219878 405922 219934 405978
rect 220002 405922 220058 405978
rect 250598 406294 250654 406350
rect 250722 406294 250778 406350
rect 250598 406170 250654 406226
rect 250722 406170 250778 406226
rect 250598 406046 250654 406102
rect 250722 406046 250778 406102
rect 250598 405922 250654 405978
rect 250722 405922 250778 405978
rect 281318 406294 281374 406350
rect 281442 406294 281498 406350
rect 281318 406170 281374 406226
rect 281442 406170 281498 406226
rect 281318 406046 281374 406102
rect 281442 406046 281498 406102
rect 281318 405922 281374 405978
rect 281442 405922 281498 405978
rect 312038 406294 312094 406350
rect 312162 406294 312218 406350
rect 312038 406170 312094 406226
rect 312162 406170 312218 406226
rect 312038 406046 312094 406102
rect 312162 406046 312218 406102
rect 312038 405922 312094 405978
rect 312162 405922 312218 405978
rect 342758 406294 342814 406350
rect 342882 406294 342938 406350
rect 342758 406170 342814 406226
rect 342882 406170 342938 406226
rect 342758 406046 342814 406102
rect 342882 406046 342938 406102
rect 342758 405922 342814 405978
rect 342882 405922 342938 405978
rect 373478 406294 373534 406350
rect 373602 406294 373658 406350
rect 373478 406170 373534 406226
rect 373602 406170 373658 406226
rect 373478 406046 373534 406102
rect 373602 406046 373658 406102
rect 373478 405922 373534 405978
rect 373602 405922 373658 405978
rect 404198 406294 404254 406350
rect 404322 406294 404378 406350
rect 404198 406170 404254 406226
rect 404322 406170 404378 406226
rect 404198 406046 404254 406102
rect 404322 406046 404378 406102
rect 404198 405922 404254 405978
rect 404322 405922 404378 405978
rect 434918 406294 434974 406350
rect 435042 406294 435098 406350
rect 434918 406170 434974 406226
rect 435042 406170 435098 406226
rect 434918 406046 434974 406102
rect 435042 406046 435098 406102
rect 434918 405922 434974 405978
rect 435042 405922 435098 405978
rect 465638 406294 465694 406350
rect 465762 406294 465818 406350
rect 465638 406170 465694 406226
rect 465762 406170 465818 406226
rect 465638 406046 465694 406102
rect 465762 406046 465818 406102
rect 465638 405922 465694 405978
rect 465762 405922 465818 405978
rect 496358 406294 496414 406350
rect 496482 406294 496538 406350
rect 496358 406170 496414 406226
rect 496482 406170 496538 406226
rect 496358 406046 496414 406102
rect 496482 406046 496538 406102
rect 496358 405922 496414 405978
rect 496482 405922 496538 405978
rect 201250 400294 201306 400350
rect 201374 400294 201430 400350
rect 201498 400294 201554 400350
rect 201622 400294 201678 400350
rect 201250 400170 201306 400226
rect 201374 400170 201430 400226
rect 201498 400170 201554 400226
rect 201622 400170 201678 400226
rect 201250 400046 201306 400102
rect 201374 400046 201430 400102
rect 201498 400046 201554 400102
rect 201622 400046 201678 400102
rect 201250 399922 201306 399978
rect 201374 399922 201430 399978
rect 201498 399922 201554 399978
rect 201622 399922 201678 399978
rect 204518 400294 204574 400350
rect 204642 400294 204698 400350
rect 204518 400170 204574 400226
rect 204642 400170 204698 400226
rect 204518 400046 204574 400102
rect 204642 400046 204698 400102
rect 204518 399922 204574 399978
rect 204642 399922 204698 399978
rect 235238 400294 235294 400350
rect 235362 400294 235418 400350
rect 235238 400170 235294 400226
rect 235362 400170 235418 400226
rect 235238 400046 235294 400102
rect 235362 400046 235418 400102
rect 235238 399922 235294 399978
rect 235362 399922 235418 399978
rect 265958 400294 266014 400350
rect 266082 400294 266138 400350
rect 265958 400170 266014 400226
rect 266082 400170 266138 400226
rect 265958 400046 266014 400102
rect 266082 400046 266138 400102
rect 265958 399922 266014 399978
rect 266082 399922 266138 399978
rect 296678 400294 296734 400350
rect 296802 400294 296858 400350
rect 296678 400170 296734 400226
rect 296802 400170 296858 400226
rect 296678 400046 296734 400102
rect 296802 400046 296858 400102
rect 296678 399922 296734 399978
rect 296802 399922 296858 399978
rect 327398 400294 327454 400350
rect 327522 400294 327578 400350
rect 327398 400170 327454 400226
rect 327522 400170 327578 400226
rect 327398 400046 327454 400102
rect 327522 400046 327578 400102
rect 327398 399922 327454 399978
rect 327522 399922 327578 399978
rect 358118 400294 358174 400350
rect 358242 400294 358298 400350
rect 358118 400170 358174 400226
rect 358242 400170 358298 400226
rect 358118 400046 358174 400102
rect 358242 400046 358298 400102
rect 358118 399922 358174 399978
rect 358242 399922 358298 399978
rect 388838 400294 388894 400350
rect 388962 400294 389018 400350
rect 388838 400170 388894 400226
rect 388962 400170 389018 400226
rect 388838 400046 388894 400102
rect 388962 400046 389018 400102
rect 388838 399922 388894 399978
rect 388962 399922 389018 399978
rect 419558 400294 419614 400350
rect 419682 400294 419738 400350
rect 419558 400170 419614 400226
rect 419682 400170 419738 400226
rect 419558 400046 419614 400102
rect 419682 400046 419738 400102
rect 419558 399922 419614 399978
rect 419682 399922 419738 399978
rect 450278 400294 450334 400350
rect 450402 400294 450458 400350
rect 450278 400170 450334 400226
rect 450402 400170 450458 400226
rect 450278 400046 450334 400102
rect 450402 400046 450458 400102
rect 450278 399922 450334 399978
rect 450402 399922 450458 399978
rect 480998 400294 481054 400350
rect 481122 400294 481178 400350
rect 480998 400170 481054 400226
rect 481122 400170 481178 400226
rect 480998 400046 481054 400102
rect 481122 400046 481178 400102
rect 480998 399922 481054 399978
rect 481122 399922 481178 399978
rect 507250 400294 507306 400350
rect 507374 400294 507430 400350
rect 507498 400294 507554 400350
rect 507622 400294 507678 400350
rect 507250 400170 507306 400226
rect 507374 400170 507430 400226
rect 507498 400170 507554 400226
rect 507622 400170 507678 400226
rect 507250 400046 507306 400102
rect 507374 400046 507430 400102
rect 507498 400046 507554 400102
rect 507622 400046 507678 400102
rect 507250 399922 507306 399978
rect 507374 399922 507430 399978
rect 507498 399922 507554 399978
rect 507622 399922 507678 399978
rect 219878 388294 219934 388350
rect 220002 388294 220058 388350
rect 219878 388170 219934 388226
rect 220002 388170 220058 388226
rect 219878 388046 219934 388102
rect 220002 388046 220058 388102
rect 219878 387922 219934 387978
rect 220002 387922 220058 387978
rect 250598 388294 250654 388350
rect 250722 388294 250778 388350
rect 250598 388170 250654 388226
rect 250722 388170 250778 388226
rect 250598 388046 250654 388102
rect 250722 388046 250778 388102
rect 250598 387922 250654 387978
rect 250722 387922 250778 387978
rect 281318 388294 281374 388350
rect 281442 388294 281498 388350
rect 281318 388170 281374 388226
rect 281442 388170 281498 388226
rect 281318 388046 281374 388102
rect 281442 388046 281498 388102
rect 281318 387922 281374 387978
rect 281442 387922 281498 387978
rect 312038 388294 312094 388350
rect 312162 388294 312218 388350
rect 312038 388170 312094 388226
rect 312162 388170 312218 388226
rect 312038 388046 312094 388102
rect 312162 388046 312218 388102
rect 312038 387922 312094 387978
rect 312162 387922 312218 387978
rect 342758 388294 342814 388350
rect 342882 388294 342938 388350
rect 342758 388170 342814 388226
rect 342882 388170 342938 388226
rect 342758 388046 342814 388102
rect 342882 388046 342938 388102
rect 342758 387922 342814 387978
rect 342882 387922 342938 387978
rect 373478 388294 373534 388350
rect 373602 388294 373658 388350
rect 373478 388170 373534 388226
rect 373602 388170 373658 388226
rect 373478 388046 373534 388102
rect 373602 388046 373658 388102
rect 373478 387922 373534 387978
rect 373602 387922 373658 387978
rect 404198 388294 404254 388350
rect 404322 388294 404378 388350
rect 404198 388170 404254 388226
rect 404322 388170 404378 388226
rect 404198 388046 404254 388102
rect 404322 388046 404378 388102
rect 404198 387922 404254 387978
rect 404322 387922 404378 387978
rect 434918 388294 434974 388350
rect 435042 388294 435098 388350
rect 434918 388170 434974 388226
rect 435042 388170 435098 388226
rect 434918 388046 434974 388102
rect 435042 388046 435098 388102
rect 434918 387922 434974 387978
rect 435042 387922 435098 387978
rect 465638 388294 465694 388350
rect 465762 388294 465818 388350
rect 465638 388170 465694 388226
rect 465762 388170 465818 388226
rect 465638 388046 465694 388102
rect 465762 388046 465818 388102
rect 465638 387922 465694 387978
rect 465762 387922 465818 387978
rect 496358 388294 496414 388350
rect 496482 388294 496538 388350
rect 496358 388170 496414 388226
rect 496482 388170 496538 388226
rect 496358 388046 496414 388102
rect 496482 388046 496538 388102
rect 496358 387922 496414 387978
rect 496482 387922 496538 387978
rect 201250 382294 201306 382350
rect 201374 382294 201430 382350
rect 201498 382294 201554 382350
rect 201622 382294 201678 382350
rect 201250 382170 201306 382226
rect 201374 382170 201430 382226
rect 201498 382170 201554 382226
rect 201622 382170 201678 382226
rect 201250 382046 201306 382102
rect 201374 382046 201430 382102
rect 201498 382046 201554 382102
rect 201622 382046 201678 382102
rect 201250 381922 201306 381978
rect 201374 381922 201430 381978
rect 201498 381922 201554 381978
rect 201622 381922 201678 381978
rect 204518 382294 204574 382350
rect 204642 382294 204698 382350
rect 204518 382170 204574 382226
rect 204642 382170 204698 382226
rect 204518 382046 204574 382102
rect 204642 382046 204698 382102
rect 204518 381922 204574 381978
rect 204642 381922 204698 381978
rect 235238 382294 235294 382350
rect 235362 382294 235418 382350
rect 235238 382170 235294 382226
rect 235362 382170 235418 382226
rect 235238 382046 235294 382102
rect 235362 382046 235418 382102
rect 235238 381922 235294 381978
rect 235362 381922 235418 381978
rect 265958 382294 266014 382350
rect 266082 382294 266138 382350
rect 265958 382170 266014 382226
rect 266082 382170 266138 382226
rect 265958 382046 266014 382102
rect 266082 382046 266138 382102
rect 265958 381922 266014 381978
rect 266082 381922 266138 381978
rect 296678 382294 296734 382350
rect 296802 382294 296858 382350
rect 296678 382170 296734 382226
rect 296802 382170 296858 382226
rect 296678 382046 296734 382102
rect 296802 382046 296858 382102
rect 296678 381922 296734 381978
rect 296802 381922 296858 381978
rect 327398 382294 327454 382350
rect 327522 382294 327578 382350
rect 327398 382170 327454 382226
rect 327522 382170 327578 382226
rect 327398 382046 327454 382102
rect 327522 382046 327578 382102
rect 327398 381922 327454 381978
rect 327522 381922 327578 381978
rect 358118 382294 358174 382350
rect 358242 382294 358298 382350
rect 358118 382170 358174 382226
rect 358242 382170 358298 382226
rect 358118 382046 358174 382102
rect 358242 382046 358298 382102
rect 358118 381922 358174 381978
rect 358242 381922 358298 381978
rect 388838 382294 388894 382350
rect 388962 382294 389018 382350
rect 388838 382170 388894 382226
rect 388962 382170 389018 382226
rect 388838 382046 388894 382102
rect 388962 382046 389018 382102
rect 388838 381922 388894 381978
rect 388962 381922 389018 381978
rect 419558 382294 419614 382350
rect 419682 382294 419738 382350
rect 419558 382170 419614 382226
rect 419682 382170 419738 382226
rect 419558 382046 419614 382102
rect 419682 382046 419738 382102
rect 419558 381922 419614 381978
rect 419682 381922 419738 381978
rect 450278 382294 450334 382350
rect 450402 382294 450458 382350
rect 450278 382170 450334 382226
rect 450402 382170 450458 382226
rect 450278 382046 450334 382102
rect 450402 382046 450458 382102
rect 450278 381922 450334 381978
rect 450402 381922 450458 381978
rect 480998 382294 481054 382350
rect 481122 382294 481178 382350
rect 480998 382170 481054 382226
rect 481122 382170 481178 382226
rect 480998 382046 481054 382102
rect 481122 382046 481178 382102
rect 480998 381922 481054 381978
rect 481122 381922 481178 381978
rect 507250 382294 507306 382350
rect 507374 382294 507430 382350
rect 507498 382294 507554 382350
rect 507622 382294 507678 382350
rect 507250 382170 507306 382226
rect 507374 382170 507430 382226
rect 507498 382170 507554 382226
rect 507622 382170 507678 382226
rect 507250 382046 507306 382102
rect 507374 382046 507430 382102
rect 507498 382046 507554 382102
rect 507622 382046 507678 382102
rect 507250 381922 507306 381978
rect 507374 381922 507430 381978
rect 507498 381922 507554 381978
rect 507622 381922 507678 381978
rect 219878 370294 219934 370350
rect 220002 370294 220058 370350
rect 219878 370170 219934 370226
rect 220002 370170 220058 370226
rect 219878 370046 219934 370102
rect 220002 370046 220058 370102
rect 219878 369922 219934 369978
rect 220002 369922 220058 369978
rect 250598 370294 250654 370350
rect 250722 370294 250778 370350
rect 250598 370170 250654 370226
rect 250722 370170 250778 370226
rect 250598 370046 250654 370102
rect 250722 370046 250778 370102
rect 250598 369922 250654 369978
rect 250722 369922 250778 369978
rect 281318 370294 281374 370350
rect 281442 370294 281498 370350
rect 281318 370170 281374 370226
rect 281442 370170 281498 370226
rect 281318 370046 281374 370102
rect 281442 370046 281498 370102
rect 281318 369922 281374 369978
rect 281442 369922 281498 369978
rect 312038 370294 312094 370350
rect 312162 370294 312218 370350
rect 312038 370170 312094 370226
rect 312162 370170 312218 370226
rect 312038 370046 312094 370102
rect 312162 370046 312218 370102
rect 312038 369922 312094 369978
rect 312162 369922 312218 369978
rect 342758 370294 342814 370350
rect 342882 370294 342938 370350
rect 342758 370170 342814 370226
rect 342882 370170 342938 370226
rect 342758 370046 342814 370102
rect 342882 370046 342938 370102
rect 342758 369922 342814 369978
rect 342882 369922 342938 369978
rect 373478 370294 373534 370350
rect 373602 370294 373658 370350
rect 373478 370170 373534 370226
rect 373602 370170 373658 370226
rect 373478 370046 373534 370102
rect 373602 370046 373658 370102
rect 373478 369922 373534 369978
rect 373602 369922 373658 369978
rect 404198 370294 404254 370350
rect 404322 370294 404378 370350
rect 404198 370170 404254 370226
rect 404322 370170 404378 370226
rect 404198 370046 404254 370102
rect 404322 370046 404378 370102
rect 404198 369922 404254 369978
rect 404322 369922 404378 369978
rect 434918 370294 434974 370350
rect 435042 370294 435098 370350
rect 434918 370170 434974 370226
rect 435042 370170 435098 370226
rect 434918 370046 434974 370102
rect 435042 370046 435098 370102
rect 434918 369922 434974 369978
rect 435042 369922 435098 369978
rect 465638 370294 465694 370350
rect 465762 370294 465818 370350
rect 465638 370170 465694 370226
rect 465762 370170 465818 370226
rect 465638 370046 465694 370102
rect 465762 370046 465818 370102
rect 465638 369922 465694 369978
rect 465762 369922 465818 369978
rect 496358 370294 496414 370350
rect 496482 370294 496538 370350
rect 496358 370170 496414 370226
rect 496482 370170 496538 370226
rect 496358 370046 496414 370102
rect 496482 370046 496538 370102
rect 496358 369922 496414 369978
rect 496482 369922 496538 369978
rect 201250 364294 201306 364350
rect 201374 364294 201430 364350
rect 201498 364294 201554 364350
rect 201622 364294 201678 364350
rect 201250 364170 201306 364226
rect 201374 364170 201430 364226
rect 201498 364170 201554 364226
rect 201622 364170 201678 364226
rect 201250 364046 201306 364102
rect 201374 364046 201430 364102
rect 201498 364046 201554 364102
rect 201622 364046 201678 364102
rect 201250 363922 201306 363978
rect 201374 363922 201430 363978
rect 201498 363922 201554 363978
rect 201622 363922 201678 363978
rect 204518 364294 204574 364350
rect 204642 364294 204698 364350
rect 204518 364170 204574 364226
rect 204642 364170 204698 364226
rect 204518 364046 204574 364102
rect 204642 364046 204698 364102
rect 204518 363922 204574 363978
rect 204642 363922 204698 363978
rect 235238 364294 235294 364350
rect 235362 364294 235418 364350
rect 235238 364170 235294 364226
rect 235362 364170 235418 364226
rect 235238 364046 235294 364102
rect 235362 364046 235418 364102
rect 235238 363922 235294 363978
rect 235362 363922 235418 363978
rect 265958 364294 266014 364350
rect 266082 364294 266138 364350
rect 265958 364170 266014 364226
rect 266082 364170 266138 364226
rect 265958 364046 266014 364102
rect 266082 364046 266138 364102
rect 265958 363922 266014 363978
rect 266082 363922 266138 363978
rect 296678 364294 296734 364350
rect 296802 364294 296858 364350
rect 296678 364170 296734 364226
rect 296802 364170 296858 364226
rect 296678 364046 296734 364102
rect 296802 364046 296858 364102
rect 296678 363922 296734 363978
rect 296802 363922 296858 363978
rect 327398 364294 327454 364350
rect 327522 364294 327578 364350
rect 327398 364170 327454 364226
rect 327522 364170 327578 364226
rect 327398 364046 327454 364102
rect 327522 364046 327578 364102
rect 327398 363922 327454 363978
rect 327522 363922 327578 363978
rect 358118 364294 358174 364350
rect 358242 364294 358298 364350
rect 358118 364170 358174 364226
rect 358242 364170 358298 364226
rect 358118 364046 358174 364102
rect 358242 364046 358298 364102
rect 358118 363922 358174 363978
rect 358242 363922 358298 363978
rect 388838 364294 388894 364350
rect 388962 364294 389018 364350
rect 388838 364170 388894 364226
rect 388962 364170 389018 364226
rect 388838 364046 388894 364102
rect 388962 364046 389018 364102
rect 388838 363922 388894 363978
rect 388962 363922 389018 363978
rect 419558 364294 419614 364350
rect 419682 364294 419738 364350
rect 419558 364170 419614 364226
rect 419682 364170 419738 364226
rect 419558 364046 419614 364102
rect 419682 364046 419738 364102
rect 419558 363922 419614 363978
rect 419682 363922 419738 363978
rect 450278 364294 450334 364350
rect 450402 364294 450458 364350
rect 450278 364170 450334 364226
rect 450402 364170 450458 364226
rect 450278 364046 450334 364102
rect 450402 364046 450458 364102
rect 450278 363922 450334 363978
rect 450402 363922 450458 363978
rect 480998 364294 481054 364350
rect 481122 364294 481178 364350
rect 480998 364170 481054 364226
rect 481122 364170 481178 364226
rect 480998 364046 481054 364102
rect 481122 364046 481178 364102
rect 480998 363922 481054 363978
rect 481122 363922 481178 363978
rect 507250 364294 507306 364350
rect 507374 364294 507430 364350
rect 507498 364294 507554 364350
rect 507622 364294 507678 364350
rect 507250 364170 507306 364226
rect 507374 364170 507430 364226
rect 507498 364170 507554 364226
rect 507622 364170 507678 364226
rect 507250 364046 507306 364102
rect 507374 364046 507430 364102
rect 507498 364046 507554 364102
rect 507622 364046 507678 364102
rect 507250 363922 507306 363978
rect 507374 363922 507430 363978
rect 507498 363922 507554 363978
rect 507622 363922 507678 363978
rect 219878 352294 219934 352350
rect 220002 352294 220058 352350
rect 219878 352170 219934 352226
rect 220002 352170 220058 352226
rect 219878 352046 219934 352102
rect 220002 352046 220058 352102
rect 219878 351922 219934 351978
rect 220002 351922 220058 351978
rect 250598 352294 250654 352350
rect 250722 352294 250778 352350
rect 250598 352170 250654 352226
rect 250722 352170 250778 352226
rect 250598 352046 250654 352102
rect 250722 352046 250778 352102
rect 250598 351922 250654 351978
rect 250722 351922 250778 351978
rect 281318 352294 281374 352350
rect 281442 352294 281498 352350
rect 281318 352170 281374 352226
rect 281442 352170 281498 352226
rect 281318 352046 281374 352102
rect 281442 352046 281498 352102
rect 281318 351922 281374 351978
rect 281442 351922 281498 351978
rect 312038 352294 312094 352350
rect 312162 352294 312218 352350
rect 312038 352170 312094 352226
rect 312162 352170 312218 352226
rect 312038 352046 312094 352102
rect 312162 352046 312218 352102
rect 312038 351922 312094 351978
rect 312162 351922 312218 351978
rect 342758 352294 342814 352350
rect 342882 352294 342938 352350
rect 342758 352170 342814 352226
rect 342882 352170 342938 352226
rect 342758 352046 342814 352102
rect 342882 352046 342938 352102
rect 342758 351922 342814 351978
rect 342882 351922 342938 351978
rect 373478 352294 373534 352350
rect 373602 352294 373658 352350
rect 373478 352170 373534 352226
rect 373602 352170 373658 352226
rect 373478 352046 373534 352102
rect 373602 352046 373658 352102
rect 373478 351922 373534 351978
rect 373602 351922 373658 351978
rect 404198 352294 404254 352350
rect 404322 352294 404378 352350
rect 404198 352170 404254 352226
rect 404322 352170 404378 352226
rect 404198 352046 404254 352102
rect 404322 352046 404378 352102
rect 404198 351922 404254 351978
rect 404322 351922 404378 351978
rect 434918 352294 434974 352350
rect 435042 352294 435098 352350
rect 434918 352170 434974 352226
rect 435042 352170 435098 352226
rect 434918 352046 434974 352102
rect 435042 352046 435098 352102
rect 434918 351922 434974 351978
rect 435042 351922 435098 351978
rect 465638 352294 465694 352350
rect 465762 352294 465818 352350
rect 465638 352170 465694 352226
rect 465762 352170 465818 352226
rect 465638 352046 465694 352102
rect 465762 352046 465818 352102
rect 465638 351922 465694 351978
rect 465762 351922 465818 351978
rect 496358 352294 496414 352350
rect 496482 352294 496538 352350
rect 496358 352170 496414 352226
rect 496482 352170 496538 352226
rect 496358 352046 496414 352102
rect 496482 352046 496538 352102
rect 496358 351922 496414 351978
rect 496482 351922 496538 351978
rect 201250 346294 201306 346350
rect 201374 346294 201430 346350
rect 201498 346294 201554 346350
rect 201622 346294 201678 346350
rect 201250 346170 201306 346226
rect 201374 346170 201430 346226
rect 201498 346170 201554 346226
rect 201622 346170 201678 346226
rect 201250 346046 201306 346102
rect 201374 346046 201430 346102
rect 201498 346046 201554 346102
rect 201622 346046 201678 346102
rect 201250 345922 201306 345978
rect 201374 345922 201430 345978
rect 201498 345922 201554 345978
rect 201622 345922 201678 345978
rect 204518 346294 204574 346350
rect 204642 346294 204698 346350
rect 204518 346170 204574 346226
rect 204642 346170 204698 346226
rect 204518 346046 204574 346102
rect 204642 346046 204698 346102
rect 204518 345922 204574 345978
rect 204642 345922 204698 345978
rect 235238 346294 235294 346350
rect 235362 346294 235418 346350
rect 235238 346170 235294 346226
rect 235362 346170 235418 346226
rect 235238 346046 235294 346102
rect 235362 346046 235418 346102
rect 235238 345922 235294 345978
rect 235362 345922 235418 345978
rect 265958 346294 266014 346350
rect 266082 346294 266138 346350
rect 265958 346170 266014 346226
rect 266082 346170 266138 346226
rect 265958 346046 266014 346102
rect 266082 346046 266138 346102
rect 265958 345922 266014 345978
rect 266082 345922 266138 345978
rect 296678 346294 296734 346350
rect 296802 346294 296858 346350
rect 296678 346170 296734 346226
rect 296802 346170 296858 346226
rect 296678 346046 296734 346102
rect 296802 346046 296858 346102
rect 296678 345922 296734 345978
rect 296802 345922 296858 345978
rect 327398 346294 327454 346350
rect 327522 346294 327578 346350
rect 327398 346170 327454 346226
rect 327522 346170 327578 346226
rect 327398 346046 327454 346102
rect 327522 346046 327578 346102
rect 327398 345922 327454 345978
rect 327522 345922 327578 345978
rect 358118 346294 358174 346350
rect 358242 346294 358298 346350
rect 358118 346170 358174 346226
rect 358242 346170 358298 346226
rect 358118 346046 358174 346102
rect 358242 346046 358298 346102
rect 358118 345922 358174 345978
rect 358242 345922 358298 345978
rect 388838 346294 388894 346350
rect 388962 346294 389018 346350
rect 388838 346170 388894 346226
rect 388962 346170 389018 346226
rect 388838 346046 388894 346102
rect 388962 346046 389018 346102
rect 388838 345922 388894 345978
rect 388962 345922 389018 345978
rect 419558 346294 419614 346350
rect 419682 346294 419738 346350
rect 419558 346170 419614 346226
rect 419682 346170 419738 346226
rect 419558 346046 419614 346102
rect 419682 346046 419738 346102
rect 419558 345922 419614 345978
rect 419682 345922 419738 345978
rect 450278 346294 450334 346350
rect 450402 346294 450458 346350
rect 450278 346170 450334 346226
rect 450402 346170 450458 346226
rect 450278 346046 450334 346102
rect 450402 346046 450458 346102
rect 450278 345922 450334 345978
rect 450402 345922 450458 345978
rect 480998 346294 481054 346350
rect 481122 346294 481178 346350
rect 480998 346170 481054 346226
rect 481122 346170 481178 346226
rect 480998 346046 481054 346102
rect 481122 346046 481178 346102
rect 480998 345922 481054 345978
rect 481122 345922 481178 345978
rect 507250 346294 507306 346350
rect 507374 346294 507430 346350
rect 507498 346294 507554 346350
rect 507622 346294 507678 346350
rect 507250 346170 507306 346226
rect 507374 346170 507430 346226
rect 507498 346170 507554 346226
rect 507622 346170 507678 346226
rect 507250 346046 507306 346102
rect 507374 346046 507430 346102
rect 507498 346046 507554 346102
rect 507622 346046 507678 346102
rect 507250 345922 507306 345978
rect 507374 345922 507430 345978
rect 507498 345922 507554 345978
rect 507622 345922 507678 345978
rect 219878 334294 219934 334350
rect 220002 334294 220058 334350
rect 219878 334170 219934 334226
rect 220002 334170 220058 334226
rect 219878 334046 219934 334102
rect 220002 334046 220058 334102
rect 219878 333922 219934 333978
rect 220002 333922 220058 333978
rect 250598 334294 250654 334350
rect 250722 334294 250778 334350
rect 250598 334170 250654 334226
rect 250722 334170 250778 334226
rect 250598 334046 250654 334102
rect 250722 334046 250778 334102
rect 250598 333922 250654 333978
rect 250722 333922 250778 333978
rect 281318 334294 281374 334350
rect 281442 334294 281498 334350
rect 281318 334170 281374 334226
rect 281442 334170 281498 334226
rect 281318 334046 281374 334102
rect 281442 334046 281498 334102
rect 281318 333922 281374 333978
rect 281442 333922 281498 333978
rect 312038 334294 312094 334350
rect 312162 334294 312218 334350
rect 312038 334170 312094 334226
rect 312162 334170 312218 334226
rect 312038 334046 312094 334102
rect 312162 334046 312218 334102
rect 312038 333922 312094 333978
rect 312162 333922 312218 333978
rect 342758 334294 342814 334350
rect 342882 334294 342938 334350
rect 342758 334170 342814 334226
rect 342882 334170 342938 334226
rect 342758 334046 342814 334102
rect 342882 334046 342938 334102
rect 342758 333922 342814 333978
rect 342882 333922 342938 333978
rect 373478 334294 373534 334350
rect 373602 334294 373658 334350
rect 373478 334170 373534 334226
rect 373602 334170 373658 334226
rect 373478 334046 373534 334102
rect 373602 334046 373658 334102
rect 373478 333922 373534 333978
rect 373602 333922 373658 333978
rect 404198 334294 404254 334350
rect 404322 334294 404378 334350
rect 404198 334170 404254 334226
rect 404322 334170 404378 334226
rect 404198 334046 404254 334102
rect 404322 334046 404378 334102
rect 404198 333922 404254 333978
rect 404322 333922 404378 333978
rect 434918 334294 434974 334350
rect 435042 334294 435098 334350
rect 434918 334170 434974 334226
rect 435042 334170 435098 334226
rect 434918 334046 434974 334102
rect 435042 334046 435098 334102
rect 434918 333922 434974 333978
rect 435042 333922 435098 333978
rect 465638 334294 465694 334350
rect 465762 334294 465818 334350
rect 465638 334170 465694 334226
rect 465762 334170 465818 334226
rect 465638 334046 465694 334102
rect 465762 334046 465818 334102
rect 465638 333922 465694 333978
rect 465762 333922 465818 333978
rect 496358 334294 496414 334350
rect 496482 334294 496538 334350
rect 496358 334170 496414 334226
rect 496482 334170 496538 334226
rect 496358 334046 496414 334102
rect 496482 334046 496538 334102
rect 496358 333922 496414 333978
rect 496482 333922 496538 333978
rect 201250 328294 201306 328350
rect 201374 328294 201430 328350
rect 201498 328294 201554 328350
rect 201622 328294 201678 328350
rect 201250 328170 201306 328226
rect 201374 328170 201430 328226
rect 201498 328170 201554 328226
rect 201622 328170 201678 328226
rect 201250 328046 201306 328102
rect 201374 328046 201430 328102
rect 201498 328046 201554 328102
rect 201622 328046 201678 328102
rect 201250 327922 201306 327978
rect 201374 327922 201430 327978
rect 201498 327922 201554 327978
rect 201622 327922 201678 327978
rect 204518 328294 204574 328350
rect 204642 328294 204698 328350
rect 204518 328170 204574 328226
rect 204642 328170 204698 328226
rect 204518 328046 204574 328102
rect 204642 328046 204698 328102
rect 204518 327922 204574 327978
rect 204642 327922 204698 327978
rect 235238 328294 235294 328350
rect 235362 328294 235418 328350
rect 235238 328170 235294 328226
rect 235362 328170 235418 328226
rect 235238 328046 235294 328102
rect 235362 328046 235418 328102
rect 235238 327922 235294 327978
rect 235362 327922 235418 327978
rect 265958 328294 266014 328350
rect 266082 328294 266138 328350
rect 265958 328170 266014 328226
rect 266082 328170 266138 328226
rect 265958 328046 266014 328102
rect 266082 328046 266138 328102
rect 265958 327922 266014 327978
rect 266082 327922 266138 327978
rect 296678 328294 296734 328350
rect 296802 328294 296858 328350
rect 296678 328170 296734 328226
rect 296802 328170 296858 328226
rect 296678 328046 296734 328102
rect 296802 328046 296858 328102
rect 296678 327922 296734 327978
rect 296802 327922 296858 327978
rect 327398 328294 327454 328350
rect 327522 328294 327578 328350
rect 327398 328170 327454 328226
rect 327522 328170 327578 328226
rect 327398 328046 327454 328102
rect 327522 328046 327578 328102
rect 327398 327922 327454 327978
rect 327522 327922 327578 327978
rect 358118 328294 358174 328350
rect 358242 328294 358298 328350
rect 358118 328170 358174 328226
rect 358242 328170 358298 328226
rect 358118 328046 358174 328102
rect 358242 328046 358298 328102
rect 358118 327922 358174 327978
rect 358242 327922 358298 327978
rect 388838 328294 388894 328350
rect 388962 328294 389018 328350
rect 388838 328170 388894 328226
rect 388962 328170 389018 328226
rect 388838 328046 388894 328102
rect 388962 328046 389018 328102
rect 388838 327922 388894 327978
rect 388962 327922 389018 327978
rect 419558 328294 419614 328350
rect 419682 328294 419738 328350
rect 419558 328170 419614 328226
rect 419682 328170 419738 328226
rect 419558 328046 419614 328102
rect 419682 328046 419738 328102
rect 419558 327922 419614 327978
rect 419682 327922 419738 327978
rect 450278 328294 450334 328350
rect 450402 328294 450458 328350
rect 450278 328170 450334 328226
rect 450402 328170 450458 328226
rect 450278 328046 450334 328102
rect 450402 328046 450458 328102
rect 450278 327922 450334 327978
rect 450402 327922 450458 327978
rect 480998 328294 481054 328350
rect 481122 328294 481178 328350
rect 480998 328170 481054 328226
rect 481122 328170 481178 328226
rect 480998 328046 481054 328102
rect 481122 328046 481178 328102
rect 480998 327922 481054 327978
rect 481122 327922 481178 327978
rect 507250 328294 507306 328350
rect 507374 328294 507430 328350
rect 507498 328294 507554 328350
rect 507622 328294 507678 328350
rect 507250 328170 507306 328226
rect 507374 328170 507430 328226
rect 507498 328170 507554 328226
rect 507622 328170 507678 328226
rect 507250 328046 507306 328102
rect 507374 328046 507430 328102
rect 507498 328046 507554 328102
rect 507622 328046 507678 328102
rect 507250 327922 507306 327978
rect 507374 327922 507430 327978
rect 507498 327922 507554 327978
rect 507622 327922 507678 327978
rect 219878 316294 219934 316350
rect 220002 316294 220058 316350
rect 219878 316170 219934 316226
rect 220002 316170 220058 316226
rect 219878 316046 219934 316102
rect 220002 316046 220058 316102
rect 219878 315922 219934 315978
rect 220002 315922 220058 315978
rect 250598 316294 250654 316350
rect 250722 316294 250778 316350
rect 250598 316170 250654 316226
rect 250722 316170 250778 316226
rect 250598 316046 250654 316102
rect 250722 316046 250778 316102
rect 250598 315922 250654 315978
rect 250722 315922 250778 315978
rect 281318 316294 281374 316350
rect 281442 316294 281498 316350
rect 281318 316170 281374 316226
rect 281442 316170 281498 316226
rect 281318 316046 281374 316102
rect 281442 316046 281498 316102
rect 281318 315922 281374 315978
rect 281442 315922 281498 315978
rect 312038 316294 312094 316350
rect 312162 316294 312218 316350
rect 312038 316170 312094 316226
rect 312162 316170 312218 316226
rect 312038 316046 312094 316102
rect 312162 316046 312218 316102
rect 312038 315922 312094 315978
rect 312162 315922 312218 315978
rect 342758 316294 342814 316350
rect 342882 316294 342938 316350
rect 342758 316170 342814 316226
rect 342882 316170 342938 316226
rect 342758 316046 342814 316102
rect 342882 316046 342938 316102
rect 342758 315922 342814 315978
rect 342882 315922 342938 315978
rect 373478 316294 373534 316350
rect 373602 316294 373658 316350
rect 373478 316170 373534 316226
rect 373602 316170 373658 316226
rect 373478 316046 373534 316102
rect 373602 316046 373658 316102
rect 373478 315922 373534 315978
rect 373602 315922 373658 315978
rect 404198 316294 404254 316350
rect 404322 316294 404378 316350
rect 404198 316170 404254 316226
rect 404322 316170 404378 316226
rect 404198 316046 404254 316102
rect 404322 316046 404378 316102
rect 404198 315922 404254 315978
rect 404322 315922 404378 315978
rect 434918 316294 434974 316350
rect 435042 316294 435098 316350
rect 434918 316170 434974 316226
rect 435042 316170 435098 316226
rect 434918 316046 434974 316102
rect 435042 316046 435098 316102
rect 434918 315922 434974 315978
rect 435042 315922 435098 315978
rect 465638 316294 465694 316350
rect 465762 316294 465818 316350
rect 465638 316170 465694 316226
rect 465762 316170 465818 316226
rect 465638 316046 465694 316102
rect 465762 316046 465818 316102
rect 465638 315922 465694 315978
rect 465762 315922 465818 315978
rect 496358 316294 496414 316350
rect 496482 316294 496538 316350
rect 496358 316170 496414 316226
rect 496482 316170 496538 316226
rect 496358 316046 496414 316102
rect 496482 316046 496538 316102
rect 496358 315922 496414 315978
rect 496482 315922 496538 315978
rect 201250 310294 201306 310350
rect 201374 310294 201430 310350
rect 201498 310294 201554 310350
rect 201622 310294 201678 310350
rect 201250 310170 201306 310226
rect 201374 310170 201430 310226
rect 201498 310170 201554 310226
rect 201622 310170 201678 310226
rect 201250 310046 201306 310102
rect 201374 310046 201430 310102
rect 201498 310046 201554 310102
rect 201622 310046 201678 310102
rect 201250 309922 201306 309978
rect 201374 309922 201430 309978
rect 201498 309922 201554 309978
rect 201622 309922 201678 309978
rect 204518 310294 204574 310350
rect 204642 310294 204698 310350
rect 204518 310170 204574 310226
rect 204642 310170 204698 310226
rect 204518 310046 204574 310102
rect 204642 310046 204698 310102
rect 204518 309922 204574 309978
rect 204642 309922 204698 309978
rect 235238 310294 235294 310350
rect 235362 310294 235418 310350
rect 235238 310170 235294 310226
rect 235362 310170 235418 310226
rect 235238 310046 235294 310102
rect 235362 310046 235418 310102
rect 235238 309922 235294 309978
rect 235362 309922 235418 309978
rect 265958 310294 266014 310350
rect 266082 310294 266138 310350
rect 265958 310170 266014 310226
rect 266082 310170 266138 310226
rect 265958 310046 266014 310102
rect 266082 310046 266138 310102
rect 265958 309922 266014 309978
rect 266082 309922 266138 309978
rect 296678 310294 296734 310350
rect 296802 310294 296858 310350
rect 296678 310170 296734 310226
rect 296802 310170 296858 310226
rect 296678 310046 296734 310102
rect 296802 310046 296858 310102
rect 296678 309922 296734 309978
rect 296802 309922 296858 309978
rect 327398 310294 327454 310350
rect 327522 310294 327578 310350
rect 327398 310170 327454 310226
rect 327522 310170 327578 310226
rect 327398 310046 327454 310102
rect 327522 310046 327578 310102
rect 327398 309922 327454 309978
rect 327522 309922 327578 309978
rect 358118 310294 358174 310350
rect 358242 310294 358298 310350
rect 358118 310170 358174 310226
rect 358242 310170 358298 310226
rect 358118 310046 358174 310102
rect 358242 310046 358298 310102
rect 358118 309922 358174 309978
rect 358242 309922 358298 309978
rect 388838 310294 388894 310350
rect 388962 310294 389018 310350
rect 388838 310170 388894 310226
rect 388962 310170 389018 310226
rect 388838 310046 388894 310102
rect 388962 310046 389018 310102
rect 388838 309922 388894 309978
rect 388962 309922 389018 309978
rect 419558 310294 419614 310350
rect 419682 310294 419738 310350
rect 419558 310170 419614 310226
rect 419682 310170 419738 310226
rect 419558 310046 419614 310102
rect 419682 310046 419738 310102
rect 419558 309922 419614 309978
rect 419682 309922 419738 309978
rect 450278 310294 450334 310350
rect 450402 310294 450458 310350
rect 450278 310170 450334 310226
rect 450402 310170 450458 310226
rect 450278 310046 450334 310102
rect 450402 310046 450458 310102
rect 450278 309922 450334 309978
rect 450402 309922 450458 309978
rect 480998 310294 481054 310350
rect 481122 310294 481178 310350
rect 480998 310170 481054 310226
rect 481122 310170 481178 310226
rect 480998 310046 481054 310102
rect 481122 310046 481178 310102
rect 480998 309922 481054 309978
rect 481122 309922 481178 309978
rect 507250 310294 507306 310350
rect 507374 310294 507430 310350
rect 507498 310294 507554 310350
rect 507622 310294 507678 310350
rect 507250 310170 507306 310226
rect 507374 310170 507430 310226
rect 507498 310170 507554 310226
rect 507622 310170 507678 310226
rect 507250 310046 507306 310102
rect 507374 310046 507430 310102
rect 507498 310046 507554 310102
rect 507622 310046 507678 310102
rect 507250 309922 507306 309978
rect 507374 309922 507430 309978
rect 507498 309922 507554 309978
rect 507622 309922 507678 309978
rect 219878 298294 219934 298350
rect 220002 298294 220058 298350
rect 219878 298170 219934 298226
rect 220002 298170 220058 298226
rect 219878 298046 219934 298102
rect 220002 298046 220058 298102
rect 219878 297922 219934 297978
rect 220002 297922 220058 297978
rect 250598 298294 250654 298350
rect 250722 298294 250778 298350
rect 250598 298170 250654 298226
rect 250722 298170 250778 298226
rect 250598 298046 250654 298102
rect 250722 298046 250778 298102
rect 250598 297922 250654 297978
rect 250722 297922 250778 297978
rect 281318 298294 281374 298350
rect 281442 298294 281498 298350
rect 281318 298170 281374 298226
rect 281442 298170 281498 298226
rect 281318 298046 281374 298102
rect 281442 298046 281498 298102
rect 281318 297922 281374 297978
rect 281442 297922 281498 297978
rect 312038 298294 312094 298350
rect 312162 298294 312218 298350
rect 312038 298170 312094 298226
rect 312162 298170 312218 298226
rect 312038 298046 312094 298102
rect 312162 298046 312218 298102
rect 312038 297922 312094 297978
rect 312162 297922 312218 297978
rect 342758 298294 342814 298350
rect 342882 298294 342938 298350
rect 342758 298170 342814 298226
rect 342882 298170 342938 298226
rect 342758 298046 342814 298102
rect 342882 298046 342938 298102
rect 342758 297922 342814 297978
rect 342882 297922 342938 297978
rect 373478 298294 373534 298350
rect 373602 298294 373658 298350
rect 373478 298170 373534 298226
rect 373602 298170 373658 298226
rect 373478 298046 373534 298102
rect 373602 298046 373658 298102
rect 373478 297922 373534 297978
rect 373602 297922 373658 297978
rect 404198 298294 404254 298350
rect 404322 298294 404378 298350
rect 404198 298170 404254 298226
rect 404322 298170 404378 298226
rect 404198 298046 404254 298102
rect 404322 298046 404378 298102
rect 404198 297922 404254 297978
rect 404322 297922 404378 297978
rect 434918 298294 434974 298350
rect 435042 298294 435098 298350
rect 434918 298170 434974 298226
rect 435042 298170 435098 298226
rect 434918 298046 434974 298102
rect 435042 298046 435098 298102
rect 434918 297922 434974 297978
rect 435042 297922 435098 297978
rect 465638 298294 465694 298350
rect 465762 298294 465818 298350
rect 465638 298170 465694 298226
rect 465762 298170 465818 298226
rect 465638 298046 465694 298102
rect 465762 298046 465818 298102
rect 465638 297922 465694 297978
rect 465762 297922 465818 297978
rect 496358 298294 496414 298350
rect 496482 298294 496538 298350
rect 496358 298170 496414 298226
rect 496482 298170 496538 298226
rect 496358 298046 496414 298102
rect 496482 298046 496538 298102
rect 496358 297922 496414 297978
rect 496482 297922 496538 297978
rect 201250 292294 201306 292350
rect 201374 292294 201430 292350
rect 201498 292294 201554 292350
rect 201622 292294 201678 292350
rect 201250 292170 201306 292226
rect 201374 292170 201430 292226
rect 201498 292170 201554 292226
rect 201622 292170 201678 292226
rect 201250 292046 201306 292102
rect 201374 292046 201430 292102
rect 201498 292046 201554 292102
rect 201622 292046 201678 292102
rect 201250 291922 201306 291978
rect 201374 291922 201430 291978
rect 201498 291922 201554 291978
rect 201622 291922 201678 291978
rect 204518 292294 204574 292350
rect 204642 292294 204698 292350
rect 204518 292170 204574 292226
rect 204642 292170 204698 292226
rect 204518 292046 204574 292102
rect 204642 292046 204698 292102
rect 204518 291922 204574 291978
rect 204642 291922 204698 291978
rect 235238 292294 235294 292350
rect 235362 292294 235418 292350
rect 235238 292170 235294 292226
rect 235362 292170 235418 292226
rect 235238 292046 235294 292102
rect 235362 292046 235418 292102
rect 235238 291922 235294 291978
rect 235362 291922 235418 291978
rect 265958 292294 266014 292350
rect 266082 292294 266138 292350
rect 265958 292170 266014 292226
rect 266082 292170 266138 292226
rect 265958 292046 266014 292102
rect 266082 292046 266138 292102
rect 265958 291922 266014 291978
rect 266082 291922 266138 291978
rect 296678 292294 296734 292350
rect 296802 292294 296858 292350
rect 296678 292170 296734 292226
rect 296802 292170 296858 292226
rect 296678 292046 296734 292102
rect 296802 292046 296858 292102
rect 296678 291922 296734 291978
rect 296802 291922 296858 291978
rect 327398 292294 327454 292350
rect 327522 292294 327578 292350
rect 327398 292170 327454 292226
rect 327522 292170 327578 292226
rect 327398 292046 327454 292102
rect 327522 292046 327578 292102
rect 327398 291922 327454 291978
rect 327522 291922 327578 291978
rect 358118 292294 358174 292350
rect 358242 292294 358298 292350
rect 358118 292170 358174 292226
rect 358242 292170 358298 292226
rect 358118 292046 358174 292102
rect 358242 292046 358298 292102
rect 358118 291922 358174 291978
rect 358242 291922 358298 291978
rect 388838 292294 388894 292350
rect 388962 292294 389018 292350
rect 388838 292170 388894 292226
rect 388962 292170 389018 292226
rect 388838 292046 388894 292102
rect 388962 292046 389018 292102
rect 388838 291922 388894 291978
rect 388962 291922 389018 291978
rect 419558 292294 419614 292350
rect 419682 292294 419738 292350
rect 419558 292170 419614 292226
rect 419682 292170 419738 292226
rect 419558 292046 419614 292102
rect 419682 292046 419738 292102
rect 419558 291922 419614 291978
rect 419682 291922 419738 291978
rect 450278 292294 450334 292350
rect 450402 292294 450458 292350
rect 450278 292170 450334 292226
rect 450402 292170 450458 292226
rect 450278 292046 450334 292102
rect 450402 292046 450458 292102
rect 450278 291922 450334 291978
rect 450402 291922 450458 291978
rect 480998 292294 481054 292350
rect 481122 292294 481178 292350
rect 480998 292170 481054 292226
rect 481122 292170 481178 292226
rect 480998 292046 481054 292102
rect 481122 292046 481178 292102
rect 480998 291922 481054 291978
rect 481122 291922 481178 291978
rect 507250 292294 507306 292350
rect 507374 292294 507430 292350
rect 507498 292294 507554 292350
rect 507622 292294 507678 292350
rect 507250 292170 507306 292226
rect 507374 292170 507430 292226
rect 507498 292170 507554 292226
rect 507622 292170 507678 292226
rect 507250 292046 507306 292102
rect 507374 292046 507430 292102
rect 507498 292046 507554 292102
rect 507622 292046 507678 292102
rect 507250 291922 507306 291978
rect 507374 291922 507430 291978
rect 507498 291922 507554 291978
rect 507622 291922 507678 291978
rect 219878 280294 219934 280350
rect 220002 280294 220058 280350
rect 219878 280170 219934 280226
rect 220002 280170 220058 280226
rect 219878 280046 219934 280102
rect 220002 280046 220058 280102
rect 219878 279922 219934 279978
rect 220002 279922 220058 279978
rect 250598 280294 250654 280350
rect 250722 280294 250778 280350
rect 250598 280170 250654 280226
rect 250722 280170 250778 280226
rect 250598 280046 250654 280102
rect 250722 280046 250778 280102
rect 250598 279922 250654 279978
rect 250722 279922 250778 279978
rect 281318 280294 281374 280350
rect 281442 280294 281498 280350
rect 281318 280170 281374 280226
rect 281442 280170 281498 280226
rect 281318 280046 281374 280102
rect 281442 280046 281498 280102
rect 281318 279922 281374 279978
rect 281442 279922 281498 279978
rect 312038 280294 312094 280350
rect 312162 280294 312218 280350
rect 312038 280170 312094 280226
rect 312162 280170 312218 280226
rect 312038 280046 312094 280102
rect 312162 280046 312218 280102
rect 312038 279922 312094 279978
rect 312162 279922 312218 279978
rect 342758 280294 342814 280350
rect 342882 280294 342938 280350
rect 342758 280170 342814 280226
rect 342882 280170 342938 280226
rect 342758 280046 342814 280102
rect 342882 280046 342938 280102
rect 342758 279922 342814 279978
rect 342882 279922 342938 279978
rect 373478 280294 373534 280350
rect 373602 280294 373658 280350
rect 373478 280170 373534 280226
rect 373602 280170 373658 280226
rect 373478 280046 373534 280102
rect 373602 280046 373658 280102
rect 373478 279922 373534 279978
rect 373602 279922 373658 279978
rect 404198 280294 404254 280350
rect 404322 280294 404378 280350
rect 404198 280170 404254 280226
rect 404322 280170 404378 280226
rect 404198 280046 404254 280102
rect 404322 280046 404378 280102
rect 404198 279922 404254 279978
rect 404322 279922 404378 279978
rect 434918 280294 434974 280350
rect 435042 280294 435098 280350
rect 434918 280170 434974 280226
rect 435042 280170 435098 280226
rect 434918 280046 434974 280102
rect 435042 280046 435098 280102
rect 434918 279922 434974 279978
rect 435042 279922 435098 279978
rect 465638 280294 465694 280350
rect 465762 280294 465818 280350
rect 465638 280170 465694 280226
rect 465762 280170 465818 280226
rect 465638 280046 465694 280102
rect 465762 280046 465818 280102
rect 465638 279922 465694 279978
rect 465762 279922 465818 279978
rect 496358 280294 496414 280350
rect 496482 280294 496538 280350
rect 496358 280170 496414 280226
rect 496482 280170 496538 280226
rect 496358 280046 496414 280102
rect 496482 280046 496538 280102
rect 496358 279922 496414 279978
rect 496482 279922 496538 279978
rect 201250 274294 201306 274350
rect 201374 274294 201430 274350
rect 201498 274294 201554 274350
rect 201622 274294 201678 274350
rect 201250 274170 201306 274226
rect 201374 274170 201430 274226
rect 201498 274170 201554 274226
rect 201622 274170 201678 274226
rect 201250 274046 201306 274102
rect 201374 274046 201430 274102
rect 201498 274046 201554 274102
rect 201622 274046 201678 274102
rect 201250 273922 201306 273978
rect 201374 273922 201430 273978
rect 201498 273922 201554 273978
rect 201622 273922 201678 273978
rect 204518 274294 204574 274350
rect 204642 274294 204698 274350
rect 204518 274170 204574 274226
rect 204642 274170 204698 274226
rect 204518 274046 204574 274102
rect 204642 274046 204698 274102
rect 204518 273922 204574 273978
rect 204642 273922 204698 273978
rect 235238 274294 235294 274350
rect 235362 274294 235418 274350
rect 235238 274170 235294 274226
rect 235362 274170 235418 274226
rect 235238 274046 235294 274102
rect 235362 274046 235418 274102
rect 235238 273922 235294 273978
rect 235362 273922 235418 273978
rect 265958 274294 266014 274350
rect 266082 274294 266138 274350
rect 265958 274170 266014 274226
rect 266082 274170 266138 274226
rect 265958 274046 266014 274102
rect 266082 274046 266138 274102
rect 265958 273922 266014 273978
rect 266082 273922 266138 273978
rect 296678 274294 296734 274350
rect 296802 274294 296858 274350
rect 296678 274170 296734 274226
rect 296802 274170 296858 274226
rect 296678 274046 296734 274102
rect 296802 274046 296858 274102
rect 296678 273922 296734 273978
rect 296802 273922 296858 273978
rect 327398 274294 327454 274350
rect 327522 274294 327578 274350
rect 327398 274170 327454 274226
rect 327522 274170 327578 274226
rect 327398 274046 327454 274102
rect 327522 274046 327578 274102
rect 327398 273922 327454 273978
rect 327522 273922 327578 273978
rect 358118 274294 358174 274350
rect 358242 274294 358298 274350
rect 358118 274170 358174 274226
rect 358242 274170 358298 274226
rect 358118 274046 358174 274102
rect 358242 274046 358298 274102
rect 358118 273922 358174 273978
rect 358242 273922 358298 273978
rect 388838 274294 388894 274350
rect 388962 274294 389018 274350
rect 388838 274170 388894 274226
rect 388962 274170 389018 274226
rect 388838 274046 388894 274102
rect 388962 274046 389018 274102
rect 388838 273922 388894 273978
rect 388962 273922 389018 273978
rect 419558 274294 419614 274350
rect 419682 274294 419738 274350
rect 419558 274170 419614 274226
rect 419682 274170 419738 274226
rect 419558 274046 419614 274102
rect 419682 274046 419738 274102
rect 419558 273922 419614 273978
rect 419682 273922 419738 273978
rect 450278 274294 450334 274350
rect 450402 274294 450458 274350
rect 450278 274170 450334 274226
rect 450402 274170 450458 274226
rect 450278 274046 450334 274102
rect 450402 274046 450458 274102
rect 450278 273922 450334 273978
rect 450402 273922 450458 273978
rect 480998 274294 481054 274350
rect 481122 274294 481178 274350
rect 480998 274170 481054 274226
rect 481122 274170 481178 274226
rect 480998 274046 481054 274102
rect 481122 274046 481178 274102
rect 480998 273922 481054 273978
rect 481122 273922 481178 273978
rect 507250 274294 507306 274350
rect 507374 274294 507430 274350
rect 507498 274294 507554 274350
rect 507622 274294 507678 274350
rect 507250 274170 507306 274226
rect 507374 274170 507430 274226
rect 507498 274170 507554 274226
rect 507622 274170 507678 274226
rect 507250 274046 507306 274102
rect 507374 274046 507430 274102
rect 507498 274046 507554 274102
rect 507622 274046 507678 274102
rect 507250 273922 507306 273978
rect 507374 273922 507430 273978
rect 507498 273922 507554 273978
rect 507622 273922 507678 273978
rect 219878 262294 219934 262350
rect 220002 262294 220058 262350
rect 219878 262170 219934 262226
rect 220002 262170 220058 262226
rect 219878 262046 219934 262102
rect 220002 262046 220058 262102
rect 219878 261922 219934 261978
rect 220002 261922 220058 261978
rect 250598 262294 250654 262350
rect 250722 262294 250778 262350
rect 250598 262170 250654 262226
rect 250722 262170 250778 262226
rect 250598 262046 250654 262102
rect 250722 262046 250778 262102
rect 250598 261922 250654 261978
rect 250722 261922 250778 261978
rect 281318 262294 281374 262350
rect 281442 262294 281498 262350
rect 281318 262170 281374 262226
rect 281442 262170 281498 262226
rect 281318 262046 281374 262102
rect 281442 262046 281498 262102
rect 281318 261922 281374 261978
rect 281442 261922 281498 261978
rect 312038 262294 312094 262350
rect 312162 262294 312218 262350
rect 312038 262170 312094 262226
rect 312162 262170 312218 262226
rect 312038 262046 312094 262102
rect 312162 262046 312218 262102
rect 312038 261922 312094 261978
rect 312162 261922 312218 261978
rect 342758 262294 342814 262350
rect 342882 262294 342938 262350
rect 342758 262170 342814 262226
rect 342882 262170 342938 262226
rect 342758 262046 342814 262102
rect 342882 262046 342938 262102
rect 342758 261922 342814 261978
rect 342882 261922 342938 261978
rect 373478 262294 373534 262350
rect 373602 262294 373658 262350
rect 373478 262170 373534 262226
rect 373602 262170 373658 262226
rect 373478 262046 373534 262102
rect 373602 262046 373658 262102
rect 373478 261922 373534 261978
rect 373602 261922 373658 261978
rect 404198 262294 404254 262350
rect 404322 262294 404378 262350
rect 404198 262170 404254 262226
rect 404322 262170 404378 262226
rect 404198 262046 404254 262102
rect 404322 262046 404378 262102
rect 404198 261922 404254 261978
rect 404322 261922 404378 261978
rect 434918 262294 434974 262350
rect 435042 262294 435098 262350
rect 434918 262170 434974 262226
rect 435042 262170 435098 262226
rect 434918 262046 434974 262102
rect 435042 262046 435098 262102
rect 434918 261922 434974 261978
rect 435042 261922 435098 261978
rect 465638 262294 465694 262350
rect 465762 262294 465818 262350
rect 465638 262170 465694 262226
rect 465762 262170 465818 262226
rect 465638 262046 465694 262102
rect 465762 262046 465818 262102
rect 465638 261922 465694 261978
rect 465762 261922 465818 261978
rect 496358 262294 496414 262350
rect 496482 262294 496538 262350
rect 496358 262170 496414 262226
rect 496482 262170 496538 262226
rect 496358 262046 496414 262102
rect 496482 262046 496538 262102
rect 496358 261922 496414 261978
rect 496482 261922 496538 261978
rect 201250 256294 201306 256350
rect 201374 256294 201430 256350
rect 201498 256294 201554 256350
rect 201622 256294 201678 256350
rect 201250 256170 201306 256226
rect 201374 256170 201430 256226
rect 201498 256170 201554 256226
rect 201622 256170 201678 256226
rect 201250 256046 201306 256102
rect 201374 256046 201430 256102
rect 201498 256046 201554 256102
rect 201622 256046 201678 256102
rect 201250 255922 201306 255978
rect 201374 255922 201430 255978
rect 201498 255922 201554 255978
rect 201622 255922 201678 255978
rect 204518 256294 204574 256350
rect 204642 256294 204698 256350
rect 204518 256170 204574 256226
rect 204642 256170 204698 256226
rect 204518 256046 204574 256102
rect 204642 256046 204698 256102
rect 204518 255922 204574 255978
rect 204642 255922 204698 255978
rect 235238 256294 235294 256350
rect 235362 256294 235418 256350
rect 235238 256170 235294 256226
rect 235362 256170 235418 256226
rect 235238 256046 235294 256102
rect 235362 256046 235418 256102
rect 235238 255922 235294 255978
rect 235362 255922 235418 255978
rect 265958 256294 266014 256350
rect 266082 256294 266138 256350
rect 265958 256170 266014 256226
rect 266082 256170 266138 256226
rect 265958 256046 266014 256102
rect 266082 256046 266138 256102
rect 265958 255922 266014 255978
rect 266082 255922 266138 255978
rect 296678 256294 296734 256350
rect 296802 256294 296858 256350
rect 296678 256170 296734 256226
rect 296802 256170 296858 256226
rect 296678 256046 296734 256102
rect 296802 256046 296858 256102
rect 296678 255922 296734 255978
rect 296802 255922 296858 255978
rect 327398 256294 327454 256350
rect 327522 256294 327578 256350
rect 327398 256170 327454 256226
rect 327522 256170 327578 256226
rect 327398 256046 327454 256102
rect 327522 256046 327578 256102
rect 327398 255922 327454 255978
rect 327522 255922 327578 255978
rect 358118 256294 358174 256350
rect 358242 256294 358298 256350
rect 358118 256170 358174 256226
rect 358242 256170 358298 256226
rect 358118 256046 358174 256102
rect 358242 256046 358298 256102
rect 358118 255922 358174 255978
rect 358242 255922 358298 255978
rect 388838 256294 388894 256350
rect 388962 256294 389018 256350
rect 388838 256170 388894 256226
rect 388962 256170 389018 256226
rect 388838 256046 388894 256102
rect 388962 256046 389018 256102
rect 388838 255922 388894 255978
rect 388962 255922 389018 255978
rect 419558 256294 419614 256350
rect 419682 256294 419738 256350
rect 419558 256170 419614 256226
rect 419682 256170 419738 256226
rect 419558 256046 419614 256102
rect 419682 256046 419738 256102
rect 419558 255922 419614 255978
rect 419682 255922 419738 255978
rect 450278 256294 450334 256350
rect 450402 256294 450458 256350
rect 450278 256170 450334 256226
rect 450402 256170 450458 256226
rect 450278 256046 450334 256102
rect 450402 256046 450458 256102
rect 450278 255922 450334 255978
rect 450402 255922 450458 255978
rect 480998 256294 481054 256350
rect 481122 256294 481178 256350
rect 480998 256170 481054 256226
rect 481122 256170 481178 256226
rect 480998 256046 481054 256102
rect 481122 256046 481178 256102
rect 480998 255922 481054 255978
rect 481122 255922 481178 255978
rect 507250 256294 507306 256350
rect 507374 256294 507430 256350
rect 507498 256294 507554 256350
rect 507622 256294 507678 256350
rect 507250 256170 507306 256226
rect 507374 256170 507430 256226
rect 507498 256170 507554 256226
rect 507622 256170 507678 256226
rect 507250 256046 507306 256102
rect 507374 256046 507430 256102
rect 507498 256046 507554 256102
rect 507622 256046 507678 256102
rect 507250 255922 507306 255978
rect 507374 255922 507430 255978
rect 507498 255922 507554 255978
rect 507622 255922 507678 255978
rect 219878 244294 219934 244350
rect 220002 244294 220058 244350
rect 219878 244170 219934 244226
rect 220002 244170 220058 244226
rect 219878 244046 219934 244102
rect 220002 244046 220058 244102
rect 219878 243922 219934 243978
rect 220002 243922 220058 243978
rect 250598 244294 250654 244350
rect 250722 244294 250778 244350
rect 250598 244170 250654 244226
rect 250722 244170 250778 244226
rect 250598 244046 250654 244102
rect 250722 244046 250778 244102
rect 250598 243922 250654 243978
rect 250722 243922 250778 243978
rect 281318 244294 281374 244350
rect 281442 244294 281498 244350
rect 281318 244170 281374 244226
rect 281442 244170 281498 244226
rect 281318 244046 281374 244102
rect 281442 244046 281498 244102
rect 281318 243922 281374 243978
rect 281442 243922 281498 243978
rect 312038 244294 312094 244350
rect 312162 244294 312218 244350
rect 312038 244170 312094 244226
rect 312162 244170 312218 244226
rect 312038 244046 312094 244102
rect 312162 244046 312218 244102
rect 312038 243922 312094 243978
rect 312162 243922 312218 243978
rect 342758 244294 342814 244350
rect 342882 244294 342938 244350
rect 342758 244170 342814 244226
rect 342882 244170 342938 244226
rect 342758 244046 342814 244102
rect 342882 244046 342938 244102
rect 342758 243922 342814 243978
rect 342882 243922 342938 243978
rect 373478 244294 373534 244350
rect 373602 244294 373658 244350
rect 373478 244170 373534 244226
rect 373602 244170 373658 244226
rect 373478 244046 373534 244102
rect 373602 244046 373658 244102
rect 373478 243922 373534 243978
rect 373602 243922 373658 243978
rect 404198 244294 404254 244350
rect 404322 244294 404378 244350
rect 404198 244170 404254 244226
rect 404322 244170 404378 244226
rect 404198 244046 404254 244102
rect 404322 244046 404378 244102
rect 404198 243922 404254 243978
rect 404322 243922 404378 243978
rect 434918 244294 434974 244350
rect 435042 244294 435098 244350
rect 434918 244170 434974 244226
rect 435042 244170 435098 244226
rect 434918 244046 434974 244102
rect 435042 244046 435098 244102
rect 434918 243922 434974 243978
rect 435042 243922 435098 243978
rect 465638 244294 465694 244350
rect 465762 244294 465818 244350
rect 465638 244170 465694 244226
rect 465762 244170 465818 244226
rect 465638 244046 465694 244102
rect 465762 244046 465818 244102
rect 465638 243922 465694 243978
rect 465762 243922 465818 243978
rect 496358 244294 496414 244350
rect 496482 244294 496538 244350
rect 496358 244170 496414 244226
rect 496482 244170 496538 244226
rect 496358 244046 496414 244102
rect 496482 244046 496538 244102
rect 496358 243922 496414 243978
rect 496482 243922 496538 243978
rect 201250 238294 201306 238350
rect 201374 238294 201430 238350
rect 201498 238294 201554 238350
rect 201622 238294 201678 238350
rect 201250 238170 201306 238226
rect 201374 238170 201430 238226
rect 201498 238170 201554 238226
rect 201622 238170 201678 238226
rect 201250 238046 201306 238102
rect 201374 238046 201430 238102
rect 201498 238046 201554 238102
rect 201622 238046 201678 238102
rect 201250 237922 201306 237978
rect 201374 237922 201430 237978
rect 201498 237922 201554 237978
rect 201622 237922 201678 237978
rect 204518 238294 204574 238350
rect 204642 238294 204698 238350
rect 204518 238170 204574 238226
rect 204642 238170 204698 238226
rect 204518 238046 204574 238102
rect 204642 238046 204698 238102
rect 204518 237922 204574 237978
rect 204642 237922 204698 237978
rect 235238 238294 235294 238350
rect 235362 238294 235418 238350
rect 235238 238170 235294 238226
rect 235362 238170 235418 238226
rect 235238 238046 235294 238102
rect 235362 238046 235418 238102
rect 235238 237922 235294 237978
rect 235362 237922 235418 237978
rect 265958 238294 266014 238350
rect 266082 238294 266138 238350
rect 265958 238170 266014 238226
rect 266082 238170 266138 238226
rect 265958 238046 266014 238102
rect 266082 238046 266138 238102
rect 265958 237922 266014 237978
rect 266082 237922 266138 237978
rect 296678 238294 296734 238350
rect 296802 238294 296858 238350
rect 296678 238170 296734 238226
rect 296802 238170 296858 238226
rect 296678 238046 296734 238102
rect 296802 238046 296858 238102
rect 296678 237922 296734 237978
rect 296802 237922 296858 237978
rect 327398 238294 327454 238350
rect 327522 238294 327578 238350
rect 327398 238170 327454 238226
rect 327522 238170 327578 238226
rect 327398 238046 327454 238102
rect 327522 238046 327578 238102
rect 327398 237922 327454 237978
rect 327522 237922 327578 237978
rect 358118 238294 358174 238350
rect 358242 238294 358298 238350
rect 358118 238170 358174 238226
rect 358242 238170 358298 238226
rect 358118 238046 358174 238102
rect 358242 238046 358298 238102
rect 358118 237922 358174 237978
rect 358242 237922 358298 237978
rect 388838 238294 388894 238350
rect 388962 238294 389018 238350
rect 388838 238170 388894 238226
rect 388962 238170 389018 238226
rect 388838 238046 388894 238102
rect 388962 238046 389018 238102
rect 388838 237922 388894 237978
rect 388962 237922 389018 237978
rect 419558 238294 419614 238350
rect 419682 238294 419738 238350
rect 419558 238170 419614 238226
rect 419682 238170 419738 238226
rect 419558 238046 419614 238102
rect 419682 238046 419738 238102
rect 419558 237922 419614 237978
rect 419682 237922 419738 237978
rect 450278 238294 450334 238350
rect 450402 238294 450458 238350
rect 450278 238170 450334 238226
rect 450402 238170 450458 238226
rect 450278 238046 450334 238102
rect 450402 238046 450458 238102
rect 450278 237922 450334 237978
rect 450402 237922 450458 237978
rect 480998 238294 481054 238350
rect 481122 238294 481178 238350
rect 480998 238170 481054 238226
rect 481122 238170 481178 238226
rect 480998 238046 481054 238102
rect 481122 238046 481178 238102
rect 480998 237922 481054 237978
rect 481122 237922 481178 237978
rect 507250 238294 507306 238350
rect 507374 238294 507430 238350
rect 507498 238294 507554 238350
rect 507622 238294 507678 238350
rect 507250 238170 507306 238226
rect 507374 238170 507430 238226
rect 507498 238170 507554 238226
rect 507622 238170 507678 238226
rect 507250 238046 507306 238102
rect 507374 238046 507430 238102
rect 507498 238046 507554 238102
rect 507622 238046 507678 238102
rect 507250 237922 507306 237978
rect 507374 237922 507430 237978
rect 507498 237922 507554 237978
rect 507622 237922 507678 237978
rect 219878 226294 219934 226350
rect 220002 226294 220058 226350
rect 219878 226170 219934 226226
rect 220002 226170 220058 226226
rect 219878 226046 219934 226102
rect 220002 226046 220058 226102
rect 219878 225922 219934 225978
rect 220002 225922 220058 225978
rect 250598 226294 250654 226350
rect 250722 226294 250778 226350
rect 250598 226170 250654 226226
rect 250722 226170 250778 226226
rect 250598 226046 250654 226102
rect 250722 226046 250778 226102
rect 250598 225922 250654 225978
rect 250722 225922 250778 225978
rect 281318 226294 281374 226350
rect 281442 226294 281498 226350
rect 281318 226170 281374 226226
rect 281442 226170 281498 226226
rect 281318 226046 281374 226102
rect 281442 226046 281498 226102
rect 281318 225922 281374 225978
rect 281442 225922 281498 225978
rect 312038 226294 312094 226350
rect 312162 226294 312218 226350
rect 312038 226170 312094 226226
rect 312162 226170 312218 226226
rect 312038 226046 312094 226102
rect 312162 226046 312218 226102
rect 312038 225922 312094 225978
rect 312162 225922 312218 225978
rect 342758 226294 342814 226350
rect 342882 226294 342938 226350
rect 342758 226170 342814 226226
rect 342882 226170 342938 226226
rect 342758 226046 342814 226102
rect 342882 226046 342938 226102
rect 342758 225922 342814 225978
rect 342882 225922 342938 225978
rect 373478 226294 373534 226350
rect 373602 226294 373658 226350
rect 373478 226170 373534 226226
rect 373602 226170 373658 226226
rect 373478 226046 373534 226102
rect 373602 226046 373658 226102
rect 373478 225922 373534 225978
rect 373602 225922 373658 225978
rect 404198 226294 404254 226350
rect 404322 226294 404378 226350
rect 404198 226170 404254 226226
rect 404322 226170 404378 226226
rect 404198 226046 404254 226102
rect 404322 226046 404378 226102
rect 404198 225922 404254 225978
rect 404322 225922 404378 225978
rect 434918 226294 434974 226350
rect 435042 226294 435098 226350
rect 434918 226170 434974 226226
rect 435042 226170 435098 226226
rect 434918 226046 434974 226102
rect 435042 226046 435098 226102
rect 434918 225922 434974 225978
rect 435042 225922 435098 225978
rect 465638 226294 465694 226350
rect 465762 226294 465818 226350
rect 465638 226170 465694 226226
rect 465762 226170 465818 226226
rect 465638 226046 465694 226102
rect 465762 226046 465818 226102
rect 465638 225922 465694 225978
rect 465762 225922 465818 225978
rect 496358 226294 496414 226350
rect 496482 226294 496538 226350
rect 496358 226170 496414 226226
rect 496482 226170 496538 226226
rect 496358 226046 496414 226102
rect 496482 226046 496538 226102
rect 496358 225922 496414 225978
rect 496482 225922 496538 225978
rect 201250 220294 201306 220350
rect 201374 220294 201430 220350
rect 201498 220294 201554 220350
rect 201622 220294 201678 220350
rect 201250 220170 201306 220226
rect 201374 220170 201430 220226
rect 201498 220170 201554 220226
rect 201622 220170 201678 220226
rect 201250 220046 201306 220102
rect 201374 220046 201430 220102
rect 201498 220046 201554 220102
rect 201622 220046 201678 220102
rect 201250 219922 201306 219978
rect 201374 219922 201430 219978
rect 201498 219922 201554 219978
rect 201622 219922 201678 219978
rect 204518 220294 204574 220350
rect 204642 220294 204698 220350
rect 204518 220170 204574 220226
rect 204642 220170 204698 220226
rect 204518 220046 204574 220102
rect 204642 220046 204698 220102
rect 204518 219922 204574 219978
rect 204642 219922 204698 219978
rect 235238 220294 235294 220350
rect 235362 220294 235418 220350
rect 235238 220170 235294 220226
rect 235362 220170 235418 220226
rect 235238 220046 235294 220102
rect 235362 220046 235418 220102
rect 235238 219922 235294 219978
rect 235362 219922 235418 219978
rect 265958 220294 266014 220350
rect 266082 220294 266138 220350
rect 265958 220170 266014 220226
rect 266082 220170 266138 220226
rect 265958 220046 266014 220102
rect 266082 220046 266138 220102
rect 265958 219922 266014 219978
rect 266082 219922 266138 219978
rect 296678 220294 296734 220350
rect 296802 220294 296858 220350
rect 296678 220170 296734 220226
rect 296802 220170 296858 220226
rect 296678 220046 296734 220102
rect 296802 220046 296858 220102
rect 296678 219922 296734 219978
rect 296802 219922 296858 219978
rect 327398 220294 327454 220350
rect 327522 220294 327578 220350
rect 327398 220170 327454 220226
rect 327522 220170 327578 220226
rect 327398 220046 327454 220102
rect 327522 220046 327578 220102
rect 327398 219922 327454 219978
rect 327522 219922 327578 219978
rect 358118 220294 358174 220350
rect 358242 220294 358298 220350
rect 358118 220170 358174 220226
rect 358242 220170 358298 220226
rect 358118 220046 358174 220102
rect 358242 220046 358298 220102
rect 358118 219922 358174 219978
rect 358242 219922 358298 219978
rect 388838 220294 388894 220350
rect 388962 220294 389018 220350
rect 388838 220170 388894 220226
rect 388962 220170 389018 220226
rect 388838 220046 388894 220102
rect 388962 220046 389018 220102
rect 388838 219922 388894 219978
rect 388962 219922 389018 219978
rect 419558 220294 419614 220350
rect 419682 220294 419738 220350
rect 419558 220170 419614 220226
rect 419682 220170 419738 220226
rect 419558 220046 419614 220102
rect 419682 220046 419738 220102
rect 419558 219922 419614 219978
rect 419682 219922 419738 219978
rect 450278 220294 450334 220350
rect 450402 220294 450458 220350
rect 450278 220170 450334 220226
rect 450402 220170 450458 220226
rect 450278 220046 450334 220102
rect 450402 220046 450458 220102
rect 450278 219922 450334 219978
rect 450402 219922 450458 219978
rect 480998 220294 481054 220350
rect 481122 220294 481178 220350
rect 480998 220170 481054 220226
rect 481122 220170 481178 220226
rect 480998 220046 481054 220102
rect 481122 220046 481178 220102
rect 480998 219922 481054 219978
rect 481122 219922 481178 219978
rect 507250 220294 507306 220350
rect 507374 220294 507430 220350
rect 507498 220294 507554 220350
rect 507622 220294 507678 220350
rect 507250 220170 507306 220226
rect 507374 220170 507430 220226
rect 507498 220170 507554 220226
rect 507622 220170 507678 220226
rect 507250 220046 507306 220102
rect 507374 220046 507430 220102
rect 507498 220046 507554 220102
rect 507622 220046 507678 220102
rect 507250 219922 507306 219978
rect 507374 219922 507430 219978
rect 507498 219922 507554 219978
rect 507622 219922 507678 219978
rect 201250 202294 201306 202350
rect 201374 202294 201430 202350
rect 201498 202294 201554 202350
rect 201622 202294 201678 202350
rect 201250 202170 201306 202226
rect 201374 202170 201430 202226
rect 201498 202170 201554 202226
rect 201622 202170 201678 202226
rect 201250 202046 201306 202102
rect 201374 202046 201430 202102
rect 201498 202046 201554 202102
rect 201622 202046 201678 202102
rect 201250 201922 201306 201978
rect 201374 201922 201430 201978
rect 201498 201922 201554 201978
rect 201622 201922 201678 201978
rect 201250 184294 201306 184350
rect 201374 184294 201430 184350
rect 201498 184294 201554 184350
rect 201622 184294 201678 184350
rect 201250 184170 201306 184226
rect 201374 184170 201430 184226
rect 201498 184170 201554 184226
rect 201622 184170 201678 184226
rect 201250 184046 201306 184102
rect 201374 184046 201430 184102
rect 201498 184046 201554 184102
rect 201622 184046 201678 184102
rect 201250 183922 201306 183978
rect 201374 183922 201430 183978
rect 201498 183922 201554 183978
rect 201622 183922 201678 183978
rect 201250 166294 201306 166350
rect 201374 166294 201430 166350
rect 201498 166294 201554 166350
rect 201622 166294 201678 166350
rect 201250 166170 201306 166226
rect 201374 166170 201430 166226
rect 201498 166170 201554 166226
rect 201622 166170 201678 166226
rect 201250 166046 201306 166102
rect 201374 166046 201430 166102
rect 201498 166046 201554 166102
rect 201622 166046 201678 166102
rect 201250 165922 201306 165978
rect 201374 165922 201430 165978
rect 201498 165922 201554 165978
rect 201622 165922 201678 165978
rect 201250 148294 201306 148350
rect 201374 148294 201430 148350
rect 201498 148294 201554 148350
rect 201622 148294 201678 148350
rect 201250 148170 201306 148226
rect 201374 148170 201430 148226
rect 201498 148170 201554 148226
rect 201622 148170 201678 148226
rect 201250 148046 201306 148102
rect 201374 148046 201430 148102
rect 201498 148046 201554 148102
rect 201622 148046 201678 148102
rect 201250 147922 201306 147978
rect 201374 147922 201430 147978
rect 201498 147922 201554 147978
rect 201622 147922 201678 147978
rect 201250 130294 201306 130350
rect 201374 130294 201430 130350
rect 201498 130294 201554 130350
rect 201622 130294 201678 130350
rect 201250 130170 201306 130226
rect 201374 130170 201430 130226
rect 201498 130170 201554 130226
rect 201622 130170 201678 130226
rect 201250 130046 201306 130102
rect 201374 130046 201430 130102
rect 201498 130046 201554 130102
rect 201622 130046 201678 130102
rect 201250 129922 201306 129978
rect 201374 129922 201430 129978
rect 201498 129922 201554 129978
rect 201622 129922 201678 129978
rect 201250 112294 201306 112350
rect 201374 112294 201430 112350
rect 201498 112294 201554 112350
rect 201622 112294 201678 112350
rect 201250 112170 201306 112226
rect 201374 112170 201430 112226
rect 201498 112170 201554 112226
rect 201622 112170 201678 112226
rect 201250 112046 201306 112102
rect 201374 112046 201430 112102
rect 201498 112046 201554 112102
rect 201622 112046 201678 112102
rect 201250 111922 201306 111978
rect 201374 111922 201430 111978
rect 201498 111922 201554 111978
rect 201622 111922 201678 111978
rect 201250 94294 201306 94350
rect 201374 94294 201430 94350
rect 201498 94294 201554 94350
rect 201622 94294 201678 94350
rect 201250 94170 201306 94226
rect 201374 94170 201430 94226
rect 201498 94170 201554 94226
rect 201622 94170 201678 94226
rect 201250 94046 201306 94102
rect 201374 94046 201430 94102
rect 201498 94046 201554 94102
rect 201622 94046 201678 94102
rect 201250 93922 201306 93978
rect 201374 93922 201430 93978
rect 201498 93922 201554 93978
rect 201622 93922 201678 93978
rect 201250 76294 201306 76350
rect 201374 76294 201430 76350
rect 201498 76294 201554 76350
rect 201622 76294 201678 76350
rect 201250 76170 201306 76226
rect 201374 76170 201430 76226
rect 201498 76170 201554 76226
rect 201622 76170 201678 76226
rect 201250 76046 201306 76102
rect 201374 76046 201430 76102
rect 201498 76046 201554 76102
rect 201622 76046 201678 76102
rect 201250 75922 201306 75978
rect 201374 75922 201430 75978
rect 201498 75922 201554 75978
rect 201622 75922 201678 75978
rect 201250 58294 201306 58350
rect 201374 58294 201430 58350
rect 201498 58294 201554 58350
rect 201622 58294 201678 58350
rect 201250 58170 201306 58226
rect 201374 58170 201430 58226
rect 201498 58170 201554 58226
rect 201622 58170 201678 58226
rect 201250 58046 201306 58102
rect 201374 58046 201430 58102
rect 201498 58046 201554 58102
rect 201622 58046 201678 58102
rect 201250 57922 201306 57978
rect 201374 57922 201430 57978
rect 201498 57922 201554 57978
rect 201622 57922 201678 57978
rect 201250 40294 201306 40350
rect 201374 40294 201430 40350
rect 201498 40294 201554 40350
rect 201622 40294 201678 40350
rect 201250 40170 201306 40226
rect 201374 40170 201430 40226
rect 201498 40170 201554 40226
rect 201622 40170 201678 40226
rect 201250 40046 201306 40102
rect 201374 40046 201430 40102
rect 201498 40046 201554 40102
rect 201622 40046 201678 40102
rect 201250 39922 201306 39978
rect 201374 39922 201430 39978
rect 201498 39922 201554 39978
rect 201622 39922 201678 39978
rect 201250 22294 201306 22350
rect 201374 22294 201430 22350
rect 201498 22294 201554 22350
rect 201622 22294 201678 22350
rect 201250 22170 201306 22226
rect 201374 22170 201430 22226
rect 201498 22170 201554 22226
rect 201622 22170 201678 22226
rect 201250 22046 201306 22102
rect 201374 22046 201430 22102
rect 201498 22046 201554 22102
rect 201622 22046 201678 22102
rect 201250 21922 201306 21978
rect 201374 21922 201430 21978
rect 201498 21922 201554 21978
rect 201622 21922 201678 21978
rect 201250 4294 201306 4350
rect 201374 4294 201430 4350
rect 201498 4294 201554 4350
rect 201622 4294 201678 4350
rect 201250 4170 201306 4226
rect 201374 4170 201430 4226
rect 201498 4170 201554 4226
rect 201622 4170 201678 4226
rect 201250 4046 201306 4102
rect 201374 4046 201430 4102
rect 201498 4046 201554 4102
rect 201622 4046 201678 4102
rect 201250 3922 201306 3978
rect 201374 3922 201430 3978
rect 201498 3922 201554 3978
rect 201622 3922 201678 3978
rect 201250 -216 201306 -160
rect 201374 -216 201430 -160
rect 201498 -216 201554 -160
rect 201622 -216 201678 -160
rect 201250 -340 201306 -284
rect 201374 -340 201430 -284
rect 201498 -340 201554 -284
rect 201622 -340 201678 -284
rect 201250 -464 201306 -408
rect 201374 -464 201430 -408
rect 201498 -464 201554 -408
rect 201622 -464 201678 -408
rect 201250 -588 201306 -532
rect 201374 -588 201430 -532
rect 201498 -588 201554 -532
rect 201622 -588 201678 -532
rect 204970 208294 205026 208350
rect 205094 208294 205150 208350
rect 205218 208294 205274 208350
rect 205342 208294 205398 208350
rect 204970 208170 205026 208226
rect 205094 208170 205150 208226
rect 205218 208170 205274 208226
rect 205342 208170 205398 208226
rect 204970 208046 205026 208102
rect 205094 208046 205150 208102
rect 205218 208046 205274 208102
rect 205342 208046 205398 208102
rect 204970 207922 205026 207978
rect 205094 207922 205150 207978
rect 205218 207922 205274 207978
rect 205342 207922 205398 207978
rect 219878 208294 219934 208350
rect 220002 208294 220058 208350
rect 219878 208170 219934 208226
rect 220002 208170 220058 208226
rect 219878 208046 219934 208102
rect 220002 208046 220058 208102
rect 219878 207922 219934 207978
rect 220002 207922 220058 207978
rect 222970 208294 223026 208350
rect 223094 208294 223150 208350
rect 223218 208294 223274 208350
rect 223342 208294 223398 208350
rect 222970 208170 223026 208226
rect 223094 208170 223150 208226
rect 223218 208170 223274 208226
rect 223342 208170 223398 208226
rect 222970 208046 223026 208102
rect 223094 208046 223150 208102
rect 223218 208046 223274 208102
rect 223342 208046 223398 208102
rect 222970 207922 223026 207978
rect 223094 207922 223150 207978
rect 223218 207922 223274 207978
rect 223342 207922 223398 207978
rect 204970 190294 205026 190350
rect 205094 190294 205150 190350
rect 205218 190294 205274 190350
rect 205342 190294 205398 190350
rect 204970 190170 205026 190226
rect 205094 190170 205150 190226
rect 205218 190170 205274 190226
rect 205342 190170 205398 190226
rect 204970 190046 205026 190102
rect 205094 190046 205150 190102
rect 205218 190046 205274 190102
rect 205342 190046 205398 190102
rect 204970 189922 205026 189978
rect 205094 189922 205150 189978
rect 205218 189922 205274 189978
rect 205342 189922 205398 189978
rect 204970 172294 205026 172350
rect 205094 172294 205150 172350
rect 205218 172294 205274 172350
rect 205342 172294 205398 172350
rect 204970 172170 205026 172226
rect 205094 172170 205150 172226
rect 205218 172170 205274 172226
rect 205342 172170 205398 172226
rect 204970 172046 205026 172102
rect 205094 172046 205150 172102
rect 205218 172046 205274 172102
rect 205342 172046 205398 172102
rect 204970 171922 205026 171978
rect 205094 171922 205150 171978
rect 205218 171922 205274 171978
rect 205342 171922 205398 171978
rect 204970 154294 205026 154350
rect 205094 154294 205150 154350
rect 205218 154294 205274 154350
rect 205342 154294 205398 154350
rect 204970 154170 205026 154226
rect 205094 154170 205150 154226
rect 205218 154170 205274 154226
rect 205342 154170 205398 154226
rect 204970 154046 205026 154102
rect 205094 154046 205150 154102
rect 205218 154046 205274 154102
rect 205342 154046 205398 154102
rect 204970 153922 205026 153978
rect 205094 153922 205150 153978
rect 205218 153922 205274 153978
rect 205342 153922 205398 153978
rect 204970 136294 205026 136350
rect 205094 136294 205150 136350
rect 205218 136294 205274 136350
rect 205342 136294 205398 136350
rect 204970 136170 205026 136226
rect 205094 136170 205150 136226
rect 205218 136170 205274 136226
rect 205342 136170 205398 136226
rect 204970 136046 205026 136102
rect 205094 136046 205150 136102
rect 205218 136046 205274 136102
rect 205342 136046 205398 136102
rect 204970 135922 205026 135978
rect 205094 135922 205150 135978
rect 205218 135922 205274 135978
rect 205342 135922 205398 135978
rect 204970 118294 205026 118350
rect 205094 118294 205150 118350
rect 205218 118294 205274 118350
rect 205342 118294 205398 118350
rect 204970 118170 205026 118226
rect 205094 118170 205150 118226
rect 205218 118170 205274 118226
rect 205342 118170 205398 118226
rect 204970 118046 205026 118102
rect 205094 118046 205150 118102
rect 205218 118046 205274 118102
rect 205342 118046 205398 118102
rect 204970 117922 205026 117978
rect 205094 117922 205150 117978
rect 205218 117922 205274 117978
rect 205342 117922 205398 117978
rect 204970 100294 205026 100350
rect 205094 100294 205150 100350
rect 205218 100294 205274 100350
rect 205342 100294 205398 100350
rect 204970 100170 205026 100226
rect 205094 100170 205150 100226
rect 205218 100170 205274 100226
rect 205342 100170 205398 100226
rect 204970 100046 205026 100102
rect 205094 100046 205150 100102
rect 205218 100046 205274 100102
rect 205342 100046 205398 100102
rect 204970 99922 205026 99978
rect 205094 99922 205150 99978
rect 205218 99922 205274 99978
rect 205342 99922 205398 99978
rect 204970 82294 205026 82350
rect 205094 82294 205150 82350
rect 205218 82294 205274 82350
rect 205342 82294 205398 82350
rect 204970 82170 205026 82226
rect 205094 82170 205150 82226
rect 205218 82170 205274 82226
rect 205342 82170 205398 82226
rect 204970 82046 205026 82102
rect 205094 82046 205150 82102
rect 205218 82046 205274 82102
rect 205342 82046 205398 82102
rect 204970 81922 205026 81978
rect 205094 81922 205150 81978
rect 205218 81922 205274 81978
rect 205342 81922 205398 81978
rect 204970 64294 205026 64350
rect 205094 64294 205150 64350
rect 205218 64294 205274 64350
rect 205342 64294 205398 64350
rect 204970 64170 205026 64226
rect 205094 64170 205150 64226
rect 205218 64170 205274 64226
rect 205342 64170 205398 64226
rect 204970 64046 205026 64102
rect 205094 64046 205150 64102
rect 205218 64046 205274 64102
rect 205342 64046 205398 64102
rect 204970 63922 205026 63978
rect 205094 63922 205150 63978
rect 205218 63922 205274 63978
rect 205342 63922 205398 63978
rect 204970 46294 205026 46350
rect 205094 46294 205150 46350
rect 205218 46294 205274 46350
rect 205342 46294 205398 46350
rect 204970 46170 205026 46226
rect 205094 46170 205150 46226
rect 205218 46170 205274 46226
rect 205342 46170 205398 46226
rect 204970 46046 205026 46102
rect 205094 46046 205150 46102
rect 205218 46046 205274 46102
rect 205342 46046 205398 46102
rect 204970 45922 205026 45978
rect 205094 45922 205150 45978
rect 205218 45922 205274 45978
rect 205342 45922 205398 45978
rect 204970 28294 205026 28350
rect 205094 28294 205150 28350
rect 205218 28294 205274 28350
rect 205342 28294 205398 28350
rect 204970 28170 205026 28226
rect 205094 28170 205150 28226
rect 205218 28170 205274 28226
rect 205342 28170 205398 28226
rect 204970 28046 205026 28102
rect 205094 28046 205150 28102
rect 205218 28046 205274 28102
rect 205342 28046 205398 28102
rect 204970 27922 205026 27978
rect 205094 27922 205150 27978
rect 205218 27922 205274 27978
rect 205342 27922 205398 27978
rect 204970 10294 205026 10350
rect 205094 10294 205150 10350
rect 205218 10294 205274 10350
rect 205342 10294 205398 10350
rect 204970 10170 205026 10226
rect 205094 10170 205150 10226
rect 205218 10170 205274 10226
rect 205342 10170 205398 10226
rect 204970 10046 205026 10102
rect 205094 10046 205150 10102
rect 205218 10046 205274 10102
rect 205342 10046 205398 10102
rect 204970 9922 205026 9978
rect 205094 9922 205150 9978
rect 205218 9922 205274 9978
rect 205342 9922 205398 9978
rect 204970 -1176 205026 -1120
rect 205094 -1176 205150 -1120
rect 205218 -1176 205274 -1120
rect 205342 -1176 205398 -1120
rect 204970 -1300 205026 -1244
rect 205094 -1300 205150 -1244
rect 205218 -1300 205274 -1244
rect 205342 -1300 205398 -1244
rect 204970 -1424 205026 -1368
rect 205094 -1424 205150 -1368
rect 205218 -1424 205274 -1368
rect 205342 -1424 205398 -1368
rect 204970 -1548 205026 -1492
rect 205094 -1548 205150 -1492
rect 205218 -1548 205274 -1492
rect 205342 -1548 205398 -1492
rect 219250 184294 219306 184350
rect 219374 184294 219430 184350
rect 219498 184294 219554 184350
rect 219622 184294 219678 184350
rect 219250 184170 219306 184226
rect 219374 184170 219430 184226
rect 219498 184170 219554 184226
rect 219622 184170 219678 184226
rect 219250 184046 219306 184102
rect 219374 184046 219430 184102
rect 219498 184046 219554 184102
rect 219622 184046 219678 184102
rect 219250 183922 219306 183978
rect 219374 183922 219430 183978
rect 219498 183922 219554 183978
rect 219622 183922 219678 183978
rect 219250 166294 219306 166350
rect 219374 166294 219430 166350
rect 219498 166294 219554 166350
rect 219622 166294 219678 166350
rect 219250 166170 219306 166226
rect 219374 166170 219430 166226
rect 219498 166170 219554 166226
rect 219622 166170 219678 166226
rect 219250 166046 219306 166102
rect 219374 166046 219430 166102
rect 219498 166046 219554 166102
rect 219622 166046 219678 166102
rect 219250 165922 219306 165978
rect 219374 165922 219430 165978
rect 219498 165922 219554 165978
rect 219622 165922 219678 165978
rect 219250 148294 219306 148350
rect 219374 148294 219430 148350
rect 219498 148294 219554 148350
rect 219622 148294 219678 148350
rect 219250 148170 219306 148226
rect 219374 148170 219430 148226
rect 219498 148170 219554 148226
rect 219622 148170 219678 148226
rect 219250 148046 219306 148102
rect 219374 148046 219430 148102
rect 219498 148046 219554 148102
rect 219622 148046 219678 148102
rect 219250 147922 219306 147978
rect 219374 147922 219430 147978
rect 219498 147922 219554 147978
rect 219622 147922 219678 147978
rect 219250 130294 219306 130350
rect 219374 130294 219430 130350
rect 219498 130294 219554 130350
rect 219622 130294 219678 130350
rect 219250 130170 219306 130226
rect 219374 130170 219430 130226
rect 219498 130170 219554 130226
rect 219622 130170 219678 130226
rect 219250 130046 219306 130102
rect 219374 130046 219430 130102
rect 219498 130046 219554 130102
rect 219622 130046 219678 130102
rect 219250 129922 219306 129978
rect 219374 129922 219430 129978
rect 219498 129922 219554 129978
rect 219622 129922 219678 129978
rect 219250 112294 219306 112350
rect 219374 112294 219430 112350
rect 219498 112294 219554 112350
rect 219622 112294 219678 112350
rect 219250 112170 219306 112226
rect 219374 112170 219430 112226
rect 219498 112170 219554 112226
rect 219622 112170 219678 112226
rect 219250 112046 219306 112102
rect 219374 112046 219430 112102
rect 219498 112046 219554 112102
rect 219622 112046 219678 112102
rect 219250 111922 219306 111978
rect 219374 111922 219430 111978
rect 219498 111922 219554 111978
rect 219622 111922 219678 111978
rect 219250 94294 219306 94350
rect 219374 94294 219430 94350
rect 219498 94294 219554 94350
rect 219622 94294 219678 94350
rect 219250 94170 219306 94226
rect 219374 94170 219430 94226
rect 219498 94170 219554 94226
rect 219622 94170 219678 94226
rect 219250 94046 219306 94102
rect 219374 94046 219430 94102
rect 219498 94046 219554 94102
rect 219622 94046 219678 94102
rect 219250 93922 219306 93978
rect 219374 93922 219430 93978
rect 219498 93922 219554 93978
rect 219622 93922 219678 93978
rect 219250 76294 219306 76350
rect 219374 76294 219430 76350
rect 219498 76294 219554 76350
rect 219622 76294 219678 76350
rect 219250 76170 219306 76226
rect 219374 76170 219430 76226
rect 219498 76170 219554 76226
rect 219622 76170 219678 76226
rect 219250 76046 219306 76102
rect 219374 76046 219430 76102
rect 219498 76046 219554 76102
rect 219622 76046 219678 76102
rect 219250 75922 219306 75978
rect 219374 75922 219430 75978
rect 219498 75922 219554 75978
rect 219622 75922 219678 75978
rect 219250 58294 219306 58350
rect 219374 58294 219430 58350
rect 219498 58294 219554 58350
rect 219622 58294 219678 58350
rect 219250 58170 219306 58226
rect 219374 58170 219430 58226
rect 219498 58170 219554 58226
rect 219622 58170 219678 58226
rect 219250 58046 219306 58102
rect 219374 58046 219430 58102
rect 219498 58046 219554 58102
rect 219622 58046 219678 58102
rect 219250 57922 219306 57978
rect 219374 57922 219430 57978
rect 219498 57922 219554 57978
rect 219622 57922 219678 57978
rect 219250 40294 219306 40350
rect 219374 40294 219430 40350
rect 219498 40294 219554 40350
rect 219622 40294 219678 40350
rect 219250 40170 219306 40226
rect 219374 40170 219430 40226
rect 219498 40170 219554 40226
rect 219622 40170 219678 40226
rect 219250 40046 219306 40102
rect 219374 40046 219430 40102
rect 219498 40046 219554 40102
rect 219622 40046 219678 40102
rect 219250 39922 219306 39978
rect 219374 39922 219430 39978
rect 219498 39922 219554 39978
rect 219622 39922 219678 39978
rect 219250 22294 219306 22350
rect 219374 22294 219430 22350
rect 219498 22294 219554 22350
rect 219622 22294 219678 22350
rect 219250 22170 219306 22226
rect 219374 22170 219430 22226
rect 219498 22170 219554 22226
rect 219622 22170 219678 22226
rect 219250 22046 219306 22102
rect 219374 22046 219430 22102
rect 219498 22046 219554 22102
rect 219622 22046 219678 22102
rect 219250 21922 219306 21978
rect 219374 21922 219430 21978
rect 219498 21922 219554 21978
rect 219622 21922 219678 21978
rect 219250 4294 219306 4350
rect 219374 4294 219430 4350
rect 219498 4294 219554 4350
rect 219622 4294 219678 4350
rect 219250 4170 219306 4226
rect 219374 4170 219430 4226
rect 219498 4170 219554 4226
rect 219622 4170 219678 4226
rect 219250 4046 219306 4102
rect 219374 4046 219430 4102
rect 219498 4046 219554 4102
rect 219622 4046 219678 4102
rect 219250 3922 219306 3978
rect 219374 3922 219430 3978
rect 219498 3922 219554 3978
rect 219622 3922 219678 3978
rect 219250 -216 219306 -160
rect 219374 -216 219430 -160
rect 219498 -216 219554 -160
rect 219622 -216 219678 -160
rect 219250 -340 219306 -284
rect 219374 -340 219430 -284
rect 219498 -340 219554 -284
rect 219622 -340 219678 -284
rect 219250 -464 219306 -408
rect 219374 -464 219430 -408
rect 219498 -464 219554 -408
rect 219622 -464 219678 -408
rect 219250 -588 219306 -532
rect 219374 -588 219430 -532
rect 219498 -588 219554 -532
rect 219622 -588 219678 -532
rect 222970 190294 223026 190350
rect 223094 190294 223150 190350
rect 223218 190294 223274 190350
rect 223342 190294 223398 190350
rect 222970 190170 223026 190226
rect 223094 190170 223150 190226
rect 223218 190170 223274 190226
rect 223342 190170 223398 190226
rect 222970 190046 223026 190102
rect 223094 190046 223150 190102
rect 223218 190046 223274 190102
rect 223342 190046 223398 190102
rect 222970 189922 223026 189978
rect 223094 189922 223150 189978
rect 223218 189922 223274 189978
rect 223342 189922 223398 189978
rect 222970 172294 223026 172350
rect 223094 172294 223150 172350
rect 223218 172294 223274 172350
rect 223342 172294 223398 172350
rect 222970 172170 223026 172226
rect 223094 172170 223150 172226
rect 223218 172170 223274 172226
rect 223342 172170 223398 172226
rect 222970 172046 223026 172102
rect 223094 172046 223150 172102
rect 223218 172046 223274 172102
rect 223342 172046 223398 172102
rect 222970 171922 223026 171978
rect 223094 171922 223150 171978
rect 223218 171922 223274 171978
rect 223342 171922 223398 171978
rect 222970 154294 223026 154350
rect 223094 154294 223150 154350
rect 223218 154294 223274 154350
rect 223342 154294 223398 154350
rect 222970 154170 223026 154226
rect 223094 154170 223150 154226
rect 223218 154170 223274 154226
rect 223342 154170 223398 154226
rect 222970 154046 223026 154102
rect 223094 154046 223150 154102
rect 223218 154046 223274 154102
rect 223342 154046 223398 154102
rect 222970 153922 223026 153978
rect 223094 153922 223150 153978
rect 223218 153922 223274 153978
rect 223342 153922 223398 153978
rect 222970 136294 223026 136350
rect 223094 136294 223150 136350
rect 223218 136294 223274 136350
rect 223342 136294 223398 136350
rect 222970 136170 223026 136226
rect 223094 136170 223150 136226
rect 223218 136170 223274 136226
rect 223342 136170 223398 136226
rect 222970 136046 223026 136102
rect 223094 136046 223150 136102
rect 223218 136046 223274 136102
rect 223342 136046 223398 136102
rect 222970 135922 223026 135978
rect 223094 135922 223150 135978
rect 223218 135922 223274 135978
rect 223342 135922 223398 135978
rect 222970 118294 223026 118350
rect 223094 118294 223150 118350
rect 223218 118294 223274 118350
rect 223342 118294 223398 118350
rect 222970 118170 223026 118226
rect 223094 118170 223150 118226
rect 223218 118170 223274 118226
rect 223342 118170 223398 118226
rect 222970 118046 223026 118102
rect 223094 118046 223150 118102
rect 223218 118046 223274 118102
rect 223342 118046 223398 118102
rect 222970 117922 223026 117978
rect 223094 117922 223150 117978
rect 223218 117922 223274 117978
rect 223342 117922 223398 117978
rect 222970 100294 223026 100350
rect 223094 100294 223150 100350
rect 223218 100294 223274 100350
rect 223342 100294 223398 100350
rect 222970 100170 223026 100226
rect 223094 100170 223150 100226
rect 223218 100170 223274 100226
rect 223342 100170 223398 100226
rect 222970 100046 223026 100102
rect 223094 100046 223150 100102
rect 223218 100046 223274 100102
rect 223342 100046 223398 100102
rect 222970 99922 223026 99978
rect 223094 99922 223150 99978
rect 223218 99922 223274 99978
rect 223342 99922 223398 99978
rect 222970 82294 223026 82350
rect 223094 82294 223150 82350
rect 223218 82294 223274 82350
rect 223342 82294 223398 82350
rect 222970 82170 223026 82226
rect 223094 82170 223150 82226
rect 223218 82170 223274 82226
rect 223342 82170 223398 82226
rect 222970 82046 223026 82102
rect 223094 82046 223150 82102
rect 223218 82046 223274 82102
rect 223342 82046 223398 82102
rect 222970 81922 223026 81978
rect 223094 81922 223150 81978
rect 223218 81922 223274 81978
rect 223342 81922 223398 81978
rect 222970 64294 223026 64350
rect 223094 64294 223150 64350
rect 223218 64294 223274 64350
rect 223342 64294 223398 64350
rect 222970 64170 223026 64226
rect 223094 64170 223150 64226
rect 223218 64170 223274 64226
rect 223342 64170 223398 64226
rect 222970 64046 223026 64102
rect 223094 64046 223150 64102
rect 223218 64046 223274 64102
rect 223342 64046 223398 64102
rect 222970 63922 223026 63978
rect 223094 63922 223150 63978
rect 223218 63922 223274 63978
rect 223342 63922 223398 63978
rect 222970 46294 223026 46350
rect 223094 46294 223150 46350
rect 223218 46294 223274 46350
rect 223342 46294 223398 46350
rect 222970 46170 223026 46226
rect 223094 46170 223150 46226
rect 223218 46170 223274 46226
rect 223342 46170 223398 46226
rect 222970 46046 223026 46102
rect 223094 46046 223150 46102
rect 223218 46046 223274 46102
rect 223342 46046 223398 46102
rect 222970 45922 223026 45978
rect 223094 45922 223150 45978
rect 223218 45922 223274 45978
rect 223342 45922 223398 45978
rect 222970 28294 223026 28350
rect 223094 28294 223150 28350
rect 223218 28294 223274 28350
rect 223342 28294 223398 28350
rect 222970 28170 223026 28226
rect 223094 28170 223150 28226
rect 223218 28170 223274 28226
rect 223342 28170 223398 28226
rect 222970 28046 223026 28102
rect 223094 28046 223150 28102
rect 223218 28046 223274 28102
rect 223342 28046 223398 28102
rect 222970 27922 223026 27978
rect 223094 27922 223150 27978
rect 223218 27922 223274 27978
rect 223342 27922 223398 27978
rect 222970 10294 223026 10350
rect 223094 10294 223150 10350
rect 223218 10294 223274 10350
rect 223342 10294 223398 10350
rect 222970 10170 223026 10226
rect 223094 10170 223150 10226
rect 223218 10170 223274 10226
rect 223342 10170 223398 10226
rect 222970 10046 223026 10102
rect 223094 10046 223150 10102
rect 223218 10046 223274 10102
rect 223342 10046 223398 10102
rect 222970 9922 223026 9978
rect 223094 9922 223150 9978
rect 223218 9922 223274 9978
rect 223342 9922 223398 9978
rect 222970 -1176 223026 -1120
rect 223094 -1176 223150 -1120
rect 223218 -1176 223274 -1120
rect 223342 -1176 223398 -1120
rect 222970 -1300 223026 -1244
rect 223094 -1300 223150 -1244
rect 223218 -1300 223274 -1244
rect 223342 -1300 223398 -1244
rect 222970 -1424 223026 -1368
rect 223094 -1424 223150 -1368
rect 223218 -1424 223274 -1368
rect 223342 -1424 223398 -1368
rect 222970 -1548 223026 -1492
rect 223094 -1548 223150 -1492
rect 223218 -1548 223274 -1492
rect 223342 -1548 223398 -1492
rect 237250 202294 237306 202350
rect 237374 202294 237430 202350
rect 237498 202294 237554 202350
rect 237622 202294 237678 202350
rect 237250 202170 237306 202226
rect 237374 202170 237430 202226
rect 237498 202170 237554 202226
rect 237622 202170 237678 202226
rect 237250 202046 237306 202102
rect 237374 202046 237430 202102
rect 237498 202046 237554 202102
rect 237622 202046 237678 202102
rect 237250 201922 237306 201978
rect 237374 201922 237430 201978
rect 237498 201922 237554 201978
rect 237622 201922 237678 201978
rect 237250 184294 237306 184350
rect 237374 184294 237430 184350
rect 237498 184294 237554 184350
rect 237622 184294 237678 184350
rect 237250 184170 237306 184226
rect 237374 184170 237430 184226
rect 237498 184170 237554 184226
rect 237622 184170 237678 184226
rect 237250 184046 237306 184102
rect 237374 184046 237430 184102
rect 237498 184046 237554 184102
rect 237622 184046 237678 184102
rect 237250 183922 237306 183978
rect 237374 183922 237430 183978
rect 237498 183922 237554 183978
rect 237622 183922 237678 183978
rect 237250 166294 237306 166350
rect 237374 166294 237430 166350
rect 237498 166294 237554 166350
rect 237622 166294 237678 166350
rect 237250 166170 237306 166226
rect 237374 166170 237430 166226
rect 237498 166170 237554 166226
rect 237622 166170 237678 166226
rect 237250 166046 237306 166102
rect 237374 166046 237430 166102
rect 237498 166046 237554 166102
rect 237622 166046 237678 166102
rect 237250 165922 237306 165978
rect 237374 165922 237430 165978
rect 237498 165922 237554 165978
rect 237622 165922 237678 165978
rect 237250 148294 237306 148350
rect 237374 148294 237430 148350
rect 237498 148294 237554 148350
rect 237622 148294 237678 148350
rect 237250 148170 237306 148226
rect 237374 148170 237430 148226
rect 237498 148170 237554 148226
rect 237622 148170 237678 148226
rect 237250 148046 237306 148102
rect 237374 148046 237430 148102
rect 237498 148046 237554 148102
rect 237622 148046 237678 148102
rect 237250 147922 237306 147978
rect 237374 147922 237430 147978
rect 237498 147922 237554 147978
rect 237622 147922 237678 147978
rect 237250 130294 237306 130350
rect 237374 130294 237430 130350
rect 237498 130294 237554 130350
rect 237622 130294 237678 130350
rect 237250 130170 237306 130226
rect 237374 130170 237430 130226
rect 237498 130170 237554 130226
rect 237622 130170 237678 130226
rect 237250 130046 237306 130102
rect 237374 130046 237430 130102
rect 237498 130046 237554 130102
rect 237622 130046 237678 130102
rect 237250 129922 237306 129978
rect 237374 129922 237430 129978
rect 237498 129922 237554 129978
rect 237622 129922 237678 129978
rect 237250 112294 237306 112350
rect 237374 112294 237430 112350
rect 237498 112294 237554 112350
rect 237622 112294 237678 112350
rect 237250 112170 237306 112226
rect 237374 112170 237430 112226
rect 237498 112170 237554 112226
rect 237622 112170 237678 112226
rect 237250 112046 237306 112102
rect 237374 112046 237430 112102
rect 237498 112046 237554 112102
rect 237622 112046 237678 112102
rect 237250 111922 237306 111978
rect 237374 111922 237430 111978
rect 237498 111922 237554 111978
rect 237622 111922 237678 111978
rect 237250 94294 237306 94350
rect 237374 94294 237430 94350
rect 237498 94294 237554 94350
rect 237622 94294 237678 94350
rect 237250 94170 237306 94226
rect 237374 94170 237430 94226
rect 237498 94170 237554 94226
rect 237622 94170 237678 94226
rect 237250 94046 237306 94102
rect 237374 94046 237430 94102
rect 237498 94046 237554 94102
rect 237622 94046 237678 94102
rect 237250 93922 237306 93978
rect 237374 93922 237430 93978
rect 237498 93922 237554 93978
rect 237622 93922 237678 93978
rect 237250 76294 237306 76350
rect 237374 76294 237430 76350
rect 237498 76294 237554 76350
rect 237622 76294 237678 76350
rect 237250 76170 237306 76226
rect 237374 76170 237430 76226
rect 237498 76170 237554 76226
rect 237622 76170 237678 76226
rect 237250 76046 237306 76102
rect 237374 76046 237430 76102
rect 237498 76046 237554 76102
rect 237622 76046 237678 76102
rect 237250 75922 237306 75978
rect 237374 75922 237430 75978
rect 237498 75922 237554 75978
rect 237622 75922 237678 75978
rect 237250 58294 237306 58350
rect 237374 58294 237430 58350
rect 237498 58294 237554 58350
rect 237622 58294 237678 58350
rect 237250 58170 237306 58226
rect 237374 58170 237430 58226
rect 237498 58170 237554 58226
rect 237622 58170 237678 58226
rect 237250 58046 237306 58102
rect 237374 58046 237430 58102
rect 237498 58046 237554 58102
rect 237622 58046 237678 58102
rect 237250 57922 237306 57978
rect 237374 57922 237430 57978
rect 237498 57922 237554 57978
rect 237622 57922 237678 57978
rect 237250 40294 237306 40350
rect 237374 40294 237430 40350
rect 237498 40294 237554 40350
rect 237622 40294 237678 40350
rect 237250 40170 237306 40226
rect 237374 40170 237430 40226
rect 237498 40170 237554 40226
rect 237622 40170 237678 40226
rect 237250 40046 237306 40102
rect 237374 40046 237430 40102
rect 237498 40046 237554 40102
rect 237622 40046 237678 40102
rect 237250 39922 237306 39978
rect 237374 39922 237430 39978
rect 237498 39922 237554 39978
rect 237622 39922 237678 39978
rect 237250 22294 237306 22350
rect 237374 22294 237430 22350
rect 237498 22294 237554 22350
rect 237622 22294 237678 22350
rect 237250 22170 237306 22226
rect 237374 22170 237430 22226
rect 237498 22170 237554 22226
rect 237622 22170 237678 22226
rect 237250 22046 237306 22102
rect 237374 22046 237430 22102
rect 237498 22046 237554 22102
rect 237622 22046 237678 22102
rect 237250 21922 237306 21978
rect 237374 21922 237430 21978
rect 237498 21922 237554 21978
rect 237622 21922 237678 21978
rect 237250 4294 237306 4350
rect 237374 4294 237430 4350
rect 237498 4294 237554 4350
rect 237622 4294 237678 4350
rect 237250 4170 237306 4226
rect 237374 4170 237430 4226
rect 237498 4170 237554 4226
rect 237622 4170 237678 4226
rect 237250 4046 237306 4102
rect 237374 4046 237430 4102
rect 237498 4046 237554 4102
rect 237622 4046 237678 4102
rect 237250 3922 237306 3978
rect 237374 3922 237430 3978
rect 237498 3922 237554 3978
rect 237622 3922 237678 3978
rect 237250 -216 237306 -160
rect 237374 -216 237430 -160
rect 237498 -216 237554 -160
rect 237622 -216 237678 -160
rect 237250 -340 237306 -284
rect 237374 -340 237430 -284
rect 237498 -340 237554 -284
rect 237622 -340 237678 -284
rect 237250 -464 237306 -408
rect 237374 -464 237430 -408
rect 237498 -464 237554 -408
rect 237622 -464 237678 -408
rect 237250 -588 237306 -532
rect 237374 -588 237430 -532
rect 237498 -588 237554 -532
rect 237622 -588 237678 -532
rect 240970 208294 241026 208350
rect 241094 208294 241150 208350
rect 241218 208294 241274 208350
rect 241342 208294 241398 208350
rect 240970 208170 241026 208226
rect 241094 208170 241150 208226
rect 241218 208170 241274 208226
rect 241342 208170 241398 208226
rect 240970 208046 241026 208102
rect 241094 208046 241150 208102
rect 241218 208046 241274 208102
rect 241342 208046 241398 208102
rect 240970 207922 241026 207978
rect 241094 207922 241150 207978
rect 241218 207922 241274 207978
rect 241342 207922 241398 207978
rect 250598 208294 250654 208350
rect 250722 208294 250778 208350
rect 250598 208170 250654 208226
rect 250722 208170 250778 208226
rect 250598 208046 250654 208102
rect 250722 208046 250778 208102
rect 250598 207922 250654 207978
rect 250722 207922 250778 207978
rect 240970 190294 241026 190350
rect 241094 190294 241150 190350
rect 241218 190294 241274 190350
rect 241342 190294 241398 190350
rect 240970 190170 241026 190226
rect 241094 190170 241150 190226
rect 241218 190170 241274 190226
rect 241342 190170 241398 190226
rect 240970 190046 241026 190102
rect 241094 190046 241150 190102
rect 241218 190046 241274 190102
rect 241342 190046 241398 190102
rect 240970 189922 241026 189978
rect 241094 189922 241150 189978
rect 241218 189922 241274 189978
rect 241342 189922 241398 189978
rect 240970 172294 241026 172350
rect 241094 172294 241150 172350
rect 241218 172294 241274 172350
rect 241342 172294 241398 172350
rect 240970 172170 241026 172226
rect 241094 172170 241150 172226
rect 241218 172170 241274 172226
rect 241342 172170 241398 172226
rect 240970 172046 241026 172102
rect 241094 172046 241150 172102
rect 241218 172046 241274 172102
rect 241342 172046 241398 172102
rect 240970 171922 241026 171978
rect 241094 171922 241150 171978
rect 241218 171922 241274 171978
rect 241342 171922 241398 171978
rect 240970 154294 241026 154350
rect 241094 154294 241150 154350
rect 241218 154294 241274 154350
rect 241342 154294 241398 154350
rect 240970 154170 241026 154226
rect 241094 154170 241150 154226
rect 241218 154170 241274 154226
rect 241342 154170 241398 154226
rect 240970 154046 241026 154102
rect 241094 154046 241150 154102
rect 241218 154046 241274 154102
rect 241342 154046 241398 154102
rect 240970 153922 241026 153978
rect 241094 153922 241150 153978
rect 241218 153922 241274 153978
rect 241342 153922 241398 153978
rect 240970 136294 241026 136350
rect 241094 136294 241150 136350
rect 241218 136294 241274 136350
rect 241342 136294 241398 136350
rect 240970 136170 241026 136226
rect 241094 136170 241150 136226
rect 241218 136170 241274 136226
rect 241342 136170 241398 136226
rect 240970 136046 241026 136102
rect 241094 136046 241150 136102
rect 241218 136046 241274 136102
rect 241342 136046 241398 136102
rect 240970 135922 241026 135978
rect 241094 135922 241150 135978
rect 241218 135922 241274 135978
rect 241342 135922 241398 135978
rect 240970 118294 241026 118350
rect 241094 118294 241150 118350
rect 241218 118294 241274 118350
rect 241342 118294 241398 118350
rect 240970 118170 241026 118226
rect 241094 118170 241150 118226
rect 241218 118170 241274 118226
rect 241342 118170 241398 118226
rect 240970 118046 241026 118102
rect 241094 118046 241150 118102
rect 241218 118046 241274 118102
rect 241342 118046 241398 118102
rect 240970 117922 241026 117978
rect 241094 117922 241150 117978
rect 241218 117922 241274 117978
rect 241342 117922 241398 117978
rect 240970 100294 241026 100350
rect 241094 100294 241150 100350
rect 241218 100294 241274 100350
rect 241342 100294 241398 100350
rect 240970 100170 241026 100226
rect 241094 100170 241150 100226
rect 241218 100170 241274 100226
rect 241342 100170 241398 100226
rect 240970 100046 241026 100102
rect 241094 100046 241150 100102
rect 241218 100046 241274 100102
rect 241342 100046 241398 100102
rect 240970 99922 241026 99978
rect 241094 99922 241150 99978
rect 241218 99922 241274 99978
rect 241342 99922 241398 99978
rect 240970 82294 241026 82350
rect 241094 82294 241150 82350
rect 241218 82294 241274 82350
rect 241342 82294 241398 82350
rect 240970 82170 241026 82226
rect 241094 82170 241150 82226
rect 241218 82170 241274 82226
rect 241342 82170 241398 82226
rect 240970 82046 241026 82102
rect 241094 82046 241150 82102
rect 241218 82046 241274 82102
rect 241342 82046 241398 82102
rect 240970 81922 241026 81978
rect 241094 81922 241150 81978
rect 241218 81922 241274 81978
rect 241342 81922 241398 81978
rect 240970 64294 241026 64350
rect 241094 64294 241150 64350
rect 241218 64294 241274 64350
rect 241342 64294 241398 64350
rect 240970 64170 241026 64226
rect 241094 64170 241150 64226
rect 241218 64170 241274 64226
rect 241342 64170 241398 64226
rect 240970 64046 241026 64102
rect 241094 64046 241150 64102
rect 241218 64046 241274 64102
rect 241342 64046 241398 64102
rect 240970 63922 241026 63978
rect 241094 63922 241150 63978
rect 241218 63922 241274 63978
rect 241342 63922 241398 63978
rect 240970 46294 241026 46350
rect 241094 46294 241150 46350
rect 241218 46294 241274 46350
rect 241342 46294 241398 46350
rect 240970 46170 241026 46226
rect 241094 46170 241150 46226
rect 241218 46170 241274 46226
rect 241342 46170 241398 46226
rect 240970 46046 241026 46102
rect 241094 46046 241150 46102
rect 241218 46046 241274 46102
rect 241342 46046 241398 46102
rect 240970 45922 241026 45978
rect 241094 45922 241150 45978
rect 241218 45922 241274 45978
rect 241342 45922 241398 45978
rect 240970 28294 241026 28350
rect 241094 28294 241150 28350
rect 241218 28294 241274 28350
rect 241342 28294 241398 28350
rect 240970 28170 241026 28226
rect 241094 28170 241150 28226
rect 241218 28170 241274 28226
rect 241342 28170 241398 28226
rect 240970 28046 241026 28102
rect 241094 28046 241150 28102
rect 241218 28046 241274 28102
rect 241342 28046 241398 28102
rect 240970 27922 241026 27978
rect 241094 27922 241150 27978
rect 241218 27922 241274 27978
rect 241342 27922 241398 27978
rect 240970 10294 241026 10350
rect 241094 10294 241150 10350
rect 241218 10294 241274 10350
rect 241342 10294 241398 10350
rect 240970 10170 241026 10226
rect 241094 10170 241150 10226
rect 241218 10170 241274 10226
rect 241342 10170 241398 10226
rect 240970 10046 241026 10102
rect 241094 10046 241150 10102
rect 241218 10046 241274 10102
rect 241342 10046 241398 10102
rect 240970 9922 241026 9978
rect 241094 9922 241150 9978
rect 241218 9922 241274 9978
rect 241342 9922 241398 9978
rect 240970 -1176 241026 -1120
rect 241094 -1176 241150 -1120
rect 241218 -1176 241274 -1120
rect 241342 -1176 241398 -1120
rect 240970 -1300 241026 -1244
rect 241094 -1300 241150 -1244
rect 241218 -1300 241274 -1244
rect 241342 -1300 241398 -1244
rect 240970 -1424 241026 -1368
rect 241094 -1424 241150 -1368
rect 241218 -1424 241274 -1368
rect 241342 -1424 241398 -1368
rect 240970 -1548 241026 -1492
rect 241094 -1548 241150 -1492
rect 241218 -1548 241274 -1492
rect 241342 -1548 241398 -1492
rect 255250 202294 255306 202350
rect 255374 202294 255430 202350
rect 255498 202294 255554 202350
rect 255622 202294 255678 202350
rect 255250 202170 255306 202226
rect 255374 202170 255430 202226
rect 255498 202170 255554 202226
rect 255622 202170 255678 202226
rect 255250 202046 255306 202102
rect 255374 202046 255430 202102
rect 255498 202046 255554 202102
rect 255622 202046 255678 202102
rect 255250 201922 255306 201978
rect 255374 201922 255430 201978
rect 255498 201922 255554 201978
rect 255622 201922 255678 201978
rect 255250 184294 255306 184350
rect 255374 184294 255430 184350
rect 255498 184294 255554 184350
rect 255622 184294 255678 184350
rect 255250 184170 255306 184226
rect 255374 184170 255430 184226
rect 255498 184170 255554 184226
rect 255622 184170 255678 184226
rect 255250 184046 255306 184102
rect 255374 184046 255430 184102
rect 255498 184046 255554 184102
rect 255622 184046 255678 184102
rect 255250 183922 255306 183978
rect 255374 183922 255430 183978
rect 255498 183922 255554 183978
rect 255622 183922 255678 183978
rect 255250 166294 255306 166350
rect 255374 166294 255430 166350
rect 255498 166294 255554 166350
rect 255622 166294 255678 166350
rect 255250 166170 255306 166226
rect 255374 166170 255430 166226
rect 255498 166170 255554 166226
rect 255622 166170 255678 166226
rect 255250 166046 255306 166102
rect 255374 166046 255430 166102
rect 255498 166046 255554 166102
rect 255622 166046 255678 166102
rect 255250 165922 255306 165978
rect 255374 165922 255430 165978
rect 255498 165922 255554 165978
rect 255622 165922 255678 165978
rect 255250 148294 255306 148350
rect 255374 148294 255430 148350
rect 255498 148294 255554 148350
rect 255622 148294 255678 148350
rect 255250 148170 255306 148226
rect 255374 148170 255430 148226
rect 255498 148170 255554 148226
rect 255622 148170 255678 148226
rect 255250 148046 255306 148102
rect 255374 148046 255430 148102
rect 255498 148046 255554 148102
rect 255622 148046 255678 148102
rect 255250 147922 255306 147978
rect 255374 147922 255430 147978
rect 255498 147922 255554 147978
rect 255622 147922 255678 147978
rect 255250 130294 255306 130350
rect 255374 130294 255430 130350
rect 255498 130294 255554 130350
rect 255622 130294 255678 130350
rect 255250 130170 255306 130226
rect 255374 130170 255430 130226
rect 255498 130170 255554 130226
rect 255622 130170 255678 130226
rect 255250 130046 255306 130102
rect 255374 130046 255430 130102
rect 255498 130046 255554 130102
rect 255622 130046 255678 130102
rect 255250 129922 255306 129978
rect 255374 129922 255430 129978
rect 255498 129922 255554 129978
rect 255622 129922 255678 129978
rect 255250 112294 255306 112350
rect 255374 112294 255430 112350
rect 255498 112294 255554 112350
rect 255622 112294 255678 112350
rect 255250 112170 255306 112226
rect 255374 112170 255430 112226
rect 255498 112170 255554 112226
rect 255622 112170 255678 112226
rect 255250 112046 255306 112102
rect 255374 112046 255430 112102
rect 255498 112046 255554 112102
rect 255622 112046 255678 112102
rect 255250 111922 255306 111978
rect 255374 111922 255430 111978
rect 255498 111922 255554 111978
rect 255622 111922 255678 111978
rect 255250 94294 255306 94350
rect 255374 94294 255430 94350
rect 255498 94294 255554 94350
rect 255622 94294 255678 94350
rect 255250 94170 255306 94226
rect 255374 94170 255430 94226
rect 255498 94170 255554 94226
rect 255622 94170 255678 94226
rect 255250 94046 255306 94102
rect 255374 94046 255430 94102
rect 255498 94046 255554 94102
rect 255622 94046 255678 94102
rect 255250 93922 255306 93978
rect 255374 93922 255430 93978
rect 255498 93922 255554 93978
rect 255622 93922 255678 93978
rect 255250 76294 255306 76350
rect 255374 76294 255430 76350
rect 255498 76294 255554 76350
rect 255622 76294 255678 76350
rect 255250 76170 255306 76226
rect 255374 76170 255430 76226
rect 255498 76170 255554 76226
rect 255622 76170 255678 76226
rect 255250 76046 255306 76102
rect 255374 76046 255430 76102
rect 255498 76046 255554 76102
rect 255622 76046 255678 76102
rect 255250 75922 255306 75978
rect 255374 75922 255430 75978
rect 255498 75922 255554 75978
rect 255622 75922 255678 75978
rect 255250 58294 255306 58350
rect 255374 58294 255430 58350
rect 255498 58294 255554 58350
rect 255622 58294 255678 58350
rect 255250 58170 255306 58226
rect 255374 58170 255430 58226
rect 255498 58170 255554 58226
rect 255622 58170 255678 58226
rect 255250 58046 255306 58102
rect 255374 58046 255430 58102
rect 255498 58046 255554 58102
rect 255622 58046 255678 58102
rect 255250 57922 255306 57978
rect 255374 57922 255430 57978
rect 255498 57922 255554 57978
rect 255622 57922 255678 57978
rect 255250 40294 255306 40350
rect 255374 40294 255430 40350
rect 255498 40294 255554 40350
rect 255622 40294 255678 40350
rect 255250 40170 255306 40226
rect 255374 40170 255430 40226
rect 255498 40170 255554 40226
rect 255622 40170 255678 40226
rect 255250 40046 255306 40102
rect 255374 40046 255430 40102
rect 255498 40046 255554 40102
rect 255622 40046 255678 40102
rect 255250 39922 255306 39978
rect 255374 39922 255430 39978
rect 255498 39922 255554 39978
rect 255622 39922 255678 39978
rect 255250 22294 255306 22350
rect 255374 22294 255430 22350
rect 255498 22294 255554 22350
rect 255622 22294 255678 22350
rect 255250 22170 255306 22226
rect 255374 22170 255430 22226
rect 255498 22170 255554 22226
rect 255622 22170 255678 22226
rect 255250 22046 255306 22102
rect 255374 22046 255430 22102
rect 255498 22046 255554 22102
rect 255622 22046 255678 22102
rect 255250 21922 255306 21978
rect 255374 21922 255430 21978
rect 255498 21922 255554 21978
rect 255622 21922 255678 21978
rect 255250 4294 255306 4350
rect 255374 4294 255430 4350
rect 255498 4294 255554 4350
rect 255622 4294 255678 4350
rect 255250 4170 255306 4226
rect 255374 4170 255430 4226
rect 255498 4170 255554 4226
rect 255622 4170 255678 4226
rect 255250 4046 255306 4102
rect 255374 4046 255430 4102
rect 255498 4046 255554 4102
rect 255622 4046 255678 4102
rect 255250 3922 255306 3978
rect 255374 3922 255430 3978
rect 255498 3922 255554 3978
rect 255622 3922 255678 3978
rect 255250 -216 255306 -160
rect 255374 -216 255430 -160
rect 255498 -216 255554 -160
rect 255622 -216 255678 -160
rect 255250 -340 255306 -284
rect 255374 -340 255430 -284
rect 255498 -340 255554 -284
rect 255622 -340 255678 -284
rect 255250 -464 255306 -408
rect 255374 -464 255430 -408
rect 255498 -464 255554 -408
rect 255622 -464 255678 -408
rect 255250 -588 255306 -532
rect 255374 -588 255430 -532
rect 255498 -588 255554 -532
rect 255622 -588 255678 -532
rect 258970 208294 259026 208350
rect 259094 208294 259150 208350
rect 259218 208294 259274 208350
rect 259342 208294 259398 208350
rect 258970 208170 259026 208226
rect 259094 208170 259150 208226
rect 259218 208170 259274 208226
rect 259342 208170 259398 208226
rect 258970 208046 259026 208102
rect 259094 208046 259150 208102
rect 259218 208046 259274 208102
rect 259342 208046 259398 208102
rect 258970 207922 259026 207978
rect 259094 207922 259150 207978
rect 259218 207922 259274 207978
rect 259342 207922 259398 207978
rect 258970 190294 259026 190350
rect 259094 190294 259150 190350
rect 259218 190294 259274 190350
rect 259342 190294 259398 190350
rect 258970 190170 259026 190226
rect 259094 190170 259150 190226
rect 259218 190170 259274 190226
rect 259342 190170 259398 190226
rect 258970 190046 259026 190102
rect 259094 190046 259150 190102
rect 259218 190046 259274 190102
rect 259342 190046 259398 190102
rect 258970 189922 259026 189978
rect 259094 189922 259150 189978
rect 259218 189922 259274 189978
rect 259342 189922 259398 189978
rect 258970 172294 259026 172350
rect 259094 172294 259150 172350
rect 259218 172294 259274 172350
rect 259342 172294 259398 172350
rect 258970 172170 259026 172226
rect 259094 172170 259150 172226
rect 259218 172170 259274 172226
rect 259342 172170 259398 172226
rect 258970 172046 259026 172102
rect 259094 172046 259150 172102
rect 259218 172046 259274 172102
rect 259342 172046 259398 172102
rect 258970 171922 259026 171978
rect 259094 171922 259150 171978
rect 259218 171922 259274 171978
rect 259342 171922 259398 171978
rect 258970 154294 259026 154350
rect 259094 154294 259150 154350
rect 259218 154294 259274 154350
rect 259342 154294 259398 154350
rect 258970 154170 259026 154226
rect 259094 154170 259150 154226
rect 259218 154170 259274 154226
rect 259342 154170 259398 154226
rect 258970 154046 259026 154102
rect 259094 154046 259150 154102
rect 259218 154046 259274 154102
rect 259342 154046 259398 154102
rect 258970 153922 259026 153978
rect 259094 153922 259150 153978
rect 259218 153922 259274 153978
rect 259342 153922 259398 153978
rect 258970 136294 259026 136350
rect 259094 136294 259150 136350
rect 259218 136294 259274 136350
rect 259342 136294 259398 136350
rect 258970 136170 259026 136226
rect 259094 136170 259150 136226
rect 259218 136170 259274 136226
rect 259342 136170 259398 136226
rect 258970 136046 259026 136102
rect 259094 136046 259150 136102
rect 259218 136046 259274 136102
rect 259342 136046 259398 136102
rect 258970 135922 259026 135978
rect 259094 135922 259150 135978
rect 259218 135922 259274 135978
rect 259342 135922 259398 135978
rect 258970 118294 259026 118350
rect 259094 118294 259150 118350
rect 259218 118294 259274 118350
rect 259342 118294 259398 118350
rect 258970 118170 259026 118226
rect 259094 118170 259150 118226
rect 259218 118170 259274 118226
rect 259342 118170 259398 118226
rect 258970 118046 259026 118102
rect 259094 118046 259150 118102
rect 259218 118046 259274 118102
rect 259342 118046 259398 118102
rect 258970 117922 259026 117978
rect 259094 117922 259150 117978
rect 259218 117922 259274 117978
rect 259342 117922 259398 117978
rect 258970 100294 259026 100350
rect 259094 100294 259150 100350
rect 259218 100294 259274 100350
rect 259342 100294 259398 100350
rect 258970 100170 259026 100226
rect 259094 100170 259150 100226
rect 259218 100170 259274 100226
rect 259342 100170 259398 100226
rect 258970 100046 259026 100102
rect 259094 100046 259150 100102
rect 259218 100046 259274 100102
rect 259342 100046 259398 100102
rect 258970 99922 259026 99978
rect 259094 99922 259150 99978
rect 259218 99922 259274 99978
rect 259342 99922 259398 99978
rect 258970 82294 259026 82350
rect 259094 82294 259150 82350
rect 259218 82294 259274 82350
rect 259342 82294 259398 82350
rect 258970 82170 259026 82226
rect 259094 82170 259150 82226
rect 259218 82170 259274 82226
rect 259342 82170 259398 82226
rect 258970 82046 259026 82102
rect 259094 82046 259150 82102
rect 259218 82046 259274 82102
rect 259342 82046 259398 82102
rect 258970 81922 259026 81978
rect 259094 81922 259150 81978
rect 259218 81922 259274 81978
rect 259342 81922 259398 81978
rect 258970 64294 259026 64350
rect 259094 64294 259150 64350
rect 259218 64294 259274 64350
rect 259342 64294 259398 64350
rect 258970 64170 259026 64226
rect 259094 64170 259150 64226
rect 259218 64170 259274 64226
rect 259342 64170 259398 64226
rect 258970 64046 259026 64102
rect 259094 64046 259150 64102
rect 259218 64046 259274 64102
rect 259342 64046 259398 64102
rect 258970 63922 259026 63978
rect 259094 63922 259150 63978
rect 259218 63922 259274 63978
rect 259342 63922 259398 63978
rect 258970 46294 259026 46350
rect 259094 46294 259150 46350
rect 259218 46294 259274 46350
rect 259342 46294 259398 46350
rect 258970 46170 259026 46226
rect 259094 46170 259150 46226
rect 259218 46170 259274 46226
rect 259342 46170 259398 46226
rect 258970 46046 259026 46102
rect 259094 46046 259150 46102
rect 259218 46046 259274 46102
rect 259342 46046 259398 46102
rect 258970 45922 259026 45978
rect 259094 45922 259150 45978
rect 259218 45922 259274 45978
rect 259342 45922 259398 45978
rect 258970 28294 259026 28350
rect 259094 28294 259150 28350
rect 259218 28294 259274 28350
rect 259342 28294 259398 28350
rect 258970 28170 259026 28226
rect 259094 28170 259150 28226
rect 259218 28170 259274 28226
rect 259342 28170 259398 28226
rect 258970 28046 259026 28102
rect 259094 28046 259150 28102
rect 259218 28046 259274 28102
rect 259342 28046 259398 28102
rect 258970 27922 259026 27978
rect 259094 27922 259150 27978
rect 259218 27922 259274 27978
rect 259342 27922 259398 27978
rect 258970 10294 259026 10350
rect 259094 10294 259150 10350
rect 259218 10294 259274 10350
rect 259342 10294 259398 10350
rect 258970 10170 259026 10226
rect 259094 10170 259150 10226
rect 259218 10170 259274 10226
rect 259342 10170 259398 10226
rect 258970 10046 259026 10102
rect 259094 10046 259150 10102
rect 259218 10046 259274 10102
rect 259342 10046 259398 10102
rect 258970 9922 259026 9978
rect 259094 9922 259150 9978
rect 259218 9922 259274 9978
rect 259342 9922 259398 9978
rect 258970 -1176 259026 -1120
rect 259094 -1176 259150 -1120
rect 259218 -1176 259274 -1120
rect 259342 -1176 259398 -1120
rect 258970 -1300 259026 -1244
rect 259094 -1300 259150 -1244
rect 259218 -1300 259274 -1244
rect 259342 -1300 259398 -1244
rect 258970 -1424 259026 -1368
rect 259094 -1424 259150 -1368
rect 259218 -1424 259274 -1368
rect 259342 -1424 259398 -1368
rect 258970 -1548 259026 -1492
rect 259094 -1548 259150 -1492
rect 259218 -1548 259274 -1492
rect 259342 -1548 259398 -1492
rect 273250 202294 273306 202350
rect 273374 202294 273430 202350
rect 273498 202294 273554 202350
rect 273622 202294 273678 202350
rect 273250 202170 273306 202226
rect 273374 202170 273430 202226
rect 273498 202170 273554 202226
rect 273622 202170 273678 202226
rect 273250 202046 273306 202102
rect 273374 202046 273430 202102
rect 273498 202046 273554 202102
rect 273622 202046 273678 202102
rect 273250 201922 273306 201978
rect 273374 201922 273430 201978
rect 273498 201922 273554 201978
rect 273622 201922 273678 201978
rect 273250 184294 273306 184350
rect 273374 184294 273430 184350
rect 273498 184294 273554 184350
rect 273622 184294 273678 184350
rect 273250 184170 273306 184226
rect 273374 184170 273430 184226
rect 273498 184170 273554 184226
rect 273622 184170 273678 184226
rect 273250 184046 273306 184102
rect 273374 184046 273430 184102
rect 273498 184046 273554 184102
rect 273622 184046 273678 184102
rect 273250 183922 273306 183978
rect 273374 183922 273430 183978
rect 273498 183922 273554 183978
rect 273622 183922 273678 183978
rect 273250 166294 273306 166350
rect 273374 166294 273430 166350
rect 273498 166294 273554 166350
rect 273622 166294 273678 166350
rect 273250 166170 273306 166226
rect 273374 166170 273430 166226
rect 273498 166170 273554 166226
rect 273622 166170 273678 166226
rect 273250 166046 273306 166102
rect 273374 166046 273430 166102
rect 273498 166046 273554 166102
rect 273622 166046 273678 166102
rect 273250 165922 273306 165978
rect 273374 165922 273430 165978
rect 273498 165922 273554 165978
rect 273622 165922 273678 165978
rect 273250 148294 273306 148350
rect 273374 148294 273430 148350
rect 273498 148294 273554 148350
rect 273622 148294 273678 148350
rect 273250 148170 273306 148226
rect 273374 148170 273430 148226
rect 273498 148170 273554 148226
rect 273622 148170 273678 148226
rect 273250 148046 273306 148102
rect 273374 148046 273430 148102
rect 273498 148046 273554 148102
rect 273622 148046 273678 148102
rect 273250 147922 273306 147978
rect 273374 147922 273430 147978
rect 273498 147922 273554 147978
rect 273622 147922 273678 147978
rect 273250 130294 273306 130350
rect 273374 130294 273430 130350
rect 273498 130294 273554 130350
rect 273622 130294 273678 130350
rect 273250 130170 273306 130226
rect 273374 130170 273430 130226
rect 273498 130170 273554 130226
rect 273622 130170 273678 130226
rect 273250 130046 273306 130102
rect 273374 130046 273430 130102
rect 273498 130046 273554 130102
rect 273622 130046 273678 130102
rect 273250 129922 273306 129978
rect 273374 129922 273430 129978
rect 273498 129922 273554 129978
rect 273622 129922 273678 129978
rect 273250 112294 273306 112350
rect 273374 112294 273430 112350
rect 273498 112294 273554 112350
rect 273622 112294 273678 112350
rect 273250 112170 273306 112226
rect 273374 112170 273430 112226
rect 273498 112170 273554 112226
rect 273622 112170 273678 112226
rect 273250 112046 273306 112102
rect 273374 112046 273430 112102
rect 273498 112046 273554 112102
rect 273622 112046 273678 112102
rect 273250 111922 273306 111978
rect 273374 111922 273430 111978
rect 273498 111922 273554 111978
rect 273622 111922 273678 111978
rect 273250 94294 273306 94350
rect 273374 94294 273430 94350
rect 273498 94294 273554 94350
rect 273622 94294 273678 94350
rect 273250 94170 273306 94226
rect 273374 94170 273430 94226
rect 273498 94170 273554 94226
rect 273622 94170 273678 94226
rect 273250 94046 273306 94102
rect 273374 94046 273430 94102
rect 273498 94046 273554 94102
rect 273622 94046 273678 94102
rect 273250 93922 273306 93978
rect 273374 93922 273430 93978
rect 273498 93922 273554 93978
rect 273622 93922 273678 93978
rect 273250 76294 273306 76350
rect 273374 76294 273430 76350
rect 273498 76294 273554 76350
rect 273622 76294 273678 76350
rect 273250 76170 273306 76226
rect 273374 76170 273430 76226
rect 273498 76170 273554 76226
rect 273622 76170 273678 76226
rect 273250 76046 273306 76102
rect 273374 76046 273430 76102
rect 273498 76046 273554 76102
rect 273622 76046 273678 76102
rect 273250 75922 273306 75978
rect 273374 75922 273430 75978
rect 273498 75922 273554 75978
rect 273622 75922 273678 75978
rect 273250 58294 273306 58350
rect 273374 58294 273430 58350
rect 273498 58294 273554 58350
rect 273622 58294 273678 58350
rect 273250 58170 273306 58226
rect 273374 58170 273430 58226
rect 273498 58170 273554 58226
rect 273622 58170 273678 58226
rect 273250 58046 273306 58102
rect 273374 58046 273430 58102
rect 273498 58046 273554 58102
rect 273622 58046 273678 58102
rect 273250 57922 273306 57978
rect 273374 57922 273430 57978
rect 273498 57922 273554 57978
rect 273622 57922 273678 57978
rect 273250 40294 273306 40350
rect 273374 40294 273430 40350
rect 273498 40294 273554 40350
rect 273622 40294 273678 40350
rect 273250 40170 273306 40226
rect 273374 40170 273430 40226
rect 273498 40170 273554 40226
rect 273622 40170 273678 40226
rect 273250 40046 273306 40102
rect 273374 40046 273430 40102
rect 273498 40046 273554 40102
rect 273622 40046 273678 40102
rect 273250 39922 273306 39978
rect 273374 39922 273430 39978
rect 273498 39922 273554 39978
rect 273622 39922 273678 39978
rect 273250 22294 273306 22350
rect 273374 22294 273430 22350
rect 273498 22294 273554 22350
rect 273622 22294 273678 22350
rect 273250 22170 273306 22226
rect 273374 22170 273430 22226
rect 273498 22170 273554 22226
rect 273622 22170 273678 22226
rect 273250 22046 273306 22102
rect 273374 22046 273430 22102
rect 273498 22046 273554 22102
rect 273622 22046 273678 22102
rect 273250 21922 273306 21978
rect 273374 21922 273430 21978
rect 273498 21922 273554 21978
rect 273622 21922 273678 21978
rect 273250 4294 273306 4350
rect 273374 4294 273430 4350
rect 273498 4294 273554 4350
rect 273622 4294 273678 4350
rect 273250 4170 273306 4226
rect 273374 4170 273430 4226
rect 273498 4170 273554 4226
rect 273622 4170 273678 4226
rect 273250 4046 273306 4102
rect 273374 4046 273430 4102
rect 273498 4046 273554 4102
rect 273622 4046 273678 4102
rect 273250 3922 273306 3978
rect 273374 3922 273430 3978
rect 273498 3922 273554 3978
rect 273622 3922 273678 3978
rect 273250 -216 273306 -160
rect 273374 -216 273430 -160
rect 273498 -216 273554 -160
rect 273622 -216 273678 -160
rect 273250 -340 273306 -284
rect 273374 -340 273430 -284
rect 273498 -340 273554 -284
rect 273622 -340 273678 -284
rect 273250 -464 273306 -408
rect 273374 -464 273430 -408
rect 273498 -464 273554 -408
rect 273622 -464 273678 -408
rect 273250 -588 273306 -532
rect 273374 -588 273430 -532
rect 273498 -588 273554 -532
rect 273622 -588 273678 -532
rect 276970 208294 277026 208350
rect 277094 208294 277150 208350
rect 277218 208294 277274 208350
rect 277342 208294 277398 208350
rect 276970 208170 277026 208226
rect 277094 208170 277150 208226
rect 277218 208170 277274 208226
rect 277342 208170 277398 208226
rect 276970 208046 277026 208102
rect 277094 208046 277150 208102
rect 277218 208046 277274 208102
rect 277342 208046 277398 208102
rect 276970 207922 277026 207978
rect 277094 207922 277150 207978
rect 277218 207922 277274 207978
rect 277342 207922 277398 207978
rect 281318 208294 281374 208350
rect 281442 208294 281498 208350
rect 281318 208170 281374 208226
rect 281442 208170 281498 208226
rect 281318 208046 281374 208102
rect 281442 208046 281498 208102
rect 281318 207922 281374 207978
rect 281442 207922 281498 207978
rect 276970 190294 277026 190350
rect 277094 190294 277150 190350
rect 277218 190294 277274 190350
rect 277342 190294 277398 190350
rect 276970 190170 277026 190226
rect 277094 190170 277150 190226
rect 277218 190170 277274 190226
rect 277342 190170 277398 190226
rect 276970 190046 277026 190102
rect 277094 190046 277150 190102
rect 277218 190046 277274 190102
rect 277342 190046 277398 190102
rect 276970 189922 277026 189978
rect 277094 189922 277150 189978
rect 277218 189922 277274 189978
rect 277342 189922 277398 189978
rect 276970 172294 277026 172350
rect 277094 172294 277150 172350
rect 277218 172294 277274 172350
rect 277342 172294 277398 172350
rect 276970 172170 277026 172226
rect 277094 172170 277150 172226
rect 277218 172170 277274 172226
rect 277342 172170 277398 172226
rect 276970 172046 277026 172102
rect 277094 172046 277150 172102
rect 277218 172046 277274 172102
rect 277342 172046 277398 172102
rect 276970 171922 277026 171978
rect 277094 171922 277150 171978
rect 277218 171922 277274 171978
rect 277342 171922 277398 171978
rect 276970 154294 277026 154350
rect 277094 154294 277150 154350
rect 277218 154294 277274 154350
rect 277342 154294 277398 154350
rect 276970 154170 277026 154226
rect 277094 154170 277150 154226
rect 277218 154170 277274 154226
rect 277342 154170 277398 154226
rect 276970 154046 277026 154102
rect 277094 154046 277150 154102
rect 277218 154046 277274 154102
rect 277342 154046 277398 154102
rect 276970 153922 277026 153978
rect 277094 153922 277150 153978
rect 277218 153922 277274 153978
rect 277342 153922 277398 153978
rect 276970 136294 277026 136350
rect 277094 136294 277150 136350
rect 277218 136294 277274 136350
rect 277342 136294 277398 136350
rect 276970 136170 277026 136226
rect 277094 136170 277150 136226
rect 277218 136170 277274 136226
rect 277342 136170 277398 136226
rect 276970 136046 277026 136102
rect 277094 136046 277150 136102
rect 277218 136046 277274 136102
rect 277342 136046 277398 136102
rect 276970 135922 277026 135978
rect 277094 135922 277150 135978
rect 277218 135922 277274 135978
rect 277342 135922 277398 135978
rect 276970 118294 277026 118350
rect 277094 118294 277150 118350
rect 277218 118294 277274 118350
rect 277342 118294 277398 118350
rect 276970 118170 277026 118226
rect 277094 118170 277150 118226
rect 277218 118170 277274 118226
rect 277342 118170 277398 118226
rect 276970 118046 277026 118102
rect 277094 118046 277150 118102
rect 277218 118046 277274 118102
rect 277342 118046 277398 118102
rect 276970 117922 277026 117978
rect 277094 117922 277150 117978
rect 277218 117922 277274 117978
rect 277342 117922 277398 117978
rect 276970 100294 277026 100350
rect 277094 100294 277150 100350
rect 277218 100294 277274 100350
rect 277342 100294 277398 100350
rect 276970 100170 277026 100226
rect 277094 100170 277150 100226
rect 277218 100170 277274 100226
rect 277342 100170 277398 100226
rect 276970 100046 277026 100102
rect 277094 100046 277150 100102
rect 277218 100046 277274 100102
rect 277342 100046 277398 100102
rect 276970 99922 277026 99978
rect 277094 99922 277150 99978
rect 277218 99922 277274 99978
rect 277342 99922 277398 99978
rect 276970 82294 277026 82350
rect 277094 82294 277150 82350
rect 277218 82294 277274 82350
rect 277342 82294 277398 82350
rect 276970 82170 277026 82226
rect 277094 82170 277150 82226
rect 277218 82170 277274 82226
rect 277342 82170 277398 82226
rect 276970 82046 277026 82102
rect 277094 82046 277150 82102
rect 277218 82046 277274 82102
rect 277342 82046 277398 82102
rect 276970 81922 277026 81978
rect 277094 81922 277150 81978
rect 277218 81922 277274 81978
rect 277342 81922 277398 81978
rect 276970 64294 277026 64350
rect 277094 64294 277150 64350
rect 277218 64294 277274 64350
rect 277342 64294 277398 64350
rect 276970 64170 277026 64226
rect 277094 64170 277150 64226
rect 277218 64170 277274 64226
rect 277342 64170 277398 64226
rect 276970 64046 277026 64102
rect 277094 64046 277150 64102
rect 277218 64046 277274 64102
rect 277342 64046 277398 64102
rect 276970 63922 277026 63978
rect 277094 63922 277150 63978
rect 277218 63922 277274 63978
rect 277342 63922 277398 63978
rect 276970 46294 277026 46350
rect 277094 46294 277150 46350
rect 277218 46294 277274 46350
rect 277342 46294 277398 46350
rect 276970 46170 277026 46226
rect 277094 46170 277150 46226
rect 277218 46170 277274 46226
rect 277342 46170 277398 46226
rect 276970 46046 277026 46102
rect 277094 46046 277150 46102
rect 277218 46046 277274 46102
rect 277342 46046 277398 46102
rect 276970 45922 277026 45978
rect 277094 45922 277150 45978
rect 277218 45922 277274 45978
rect 277342 45922 277398 45978
rect 276970 28294 277026 28350
rect 277094 28294 277150 28350
rect 277218 28294 277274 28350
rect 277342 28294 277398 28350
rect 276970 28170 277026 28226
rect 277094 28170 277150 28226
rect 277218 28170 277274 28226
rect 277342 28170 277398 28226
rect 276970 28046 277026 28102
rect 277094 28046 277150 28102
rect 277218 28046 277274 28102
rect 277342 28046 277398 28102
rect 276970 27922 277026 27978
rect 277094 27922 277150 27978
rect 277218 27922 277274 27978
rect 277342 27922 277398 27978
rect 276970 10294 277026 10350
rect 277094 10294 277150 10350
rect 277218 10294 277274 10350
rect 277342 10294 277398 10350
rect 276970 10170 277026 10226
rect 277094 10170 277150 10226
rect 277218 10170 277274 10226
rect 277342 10170 277398 10226
rect 276970 10046 277026 10102
rect 277094 10046 277150 10102
rect 277218 10046 277274 10102
rect 277342 10046 277398 10102
rect 276970 9922 277026 9978
rect 277094 9922 277150 9978
rect 277218 9922 277274 9978
rect 277342 9922 277398 9978
rect 276970 -1176 277026 -1120
rect 277094 -1176 277150 -1120
rect 277218 -1176 277274 -1120
rect 277342 -1176 277398 -1120
rect 276970 -1300 277026 -1244
rect 277094 -1300 277150 -1244
rect 277218 -1300 277274 -1244
rect 277342 -1300 277398 -1244
rect 276970 -1424 277026 -1368
rect 277094 -1424 277150 -1368
rect 277218 -1424 277274 -1368
rect 277342 -1424 277398 -1368
rect 276970 -1548 277026 -1492
rect 277094 -1548 277150 -1492
rect 277218 -1548 277274 -1492
rect 277342 -1548 277398 -1492
rect 291250 202294 291306 202350
rect 291374 202294 291430 202350
rect 291498 202294 291554 202350
rect 291622 202294 291678 202350
rect 291250 202170 291306 202226
rect 291374 202170 291430 202226
rect 291498 202170 291554 202226
rect 291622 202170 291678 202226
rect 291250 202046 291306 202102
rect 291374 202046 291430 202102
rect 291498 202046 291554 202102
rect 291622 202046 291678 202102
rect 291250 201922 291306 201978
rect 291374 201922 291430 201978
rect 291498 201922 291554 201978
rect 291622 201922 291678 201978
rect 291250 184294 291306 184350
rect 291374 184294 291430 184350
rect 291498 184294 291554 184350
rect 291622 184294 291678 184350
rect 291250 184170 291306 184226
rect 291374 184170 291430 184226
rect 291498 184170 291554 184226
rect 291622 184170 291678 184226
rect 291250 184046 291306 184102
rect 291374 184046 291430 184102
rect 291498 184046 291554 184102
rect 291622 184046 291678 184102
rect 291250 183922 291306 183978
rect 291374 183922 291430 183978
rect 291498 183922 291554 183978
rect 291622 183922 291678 183978
rect 291250 166294 291306 166350
rect 291374 166294 291430 166350
rect 291498 166294 291554 166350
rect 291622 166294 291678 166350
rect 291250 166170 291306 166226
rect 291374 166170 291430 166226
rect 291498 166170 291554 166226
rect 291622 166170 291678 166226
rect 291250 166046 291306 166102
rect 291374 166046 291430 166102
rect 291498 166046 291554 166102
rect 291622 166046 291678 166102
rect 291250 165922 291306 165978
rect 291374 165922 291430 165978
rect 291498 165922 291554 165978
rect 291622 165922 291678 165978
rect 291250 148294 291306 148350
rect 291374 148294 291430 148350
rect 291498 148294 291554 148350
rect 291622 148294 291678 148350
rect 291250 148170 291306 148226
rect 291374 148170 291430 148226
rect 291498 148170 291554 148226
rect 291622 148170 291678 148226
rect 291250 148046 291306 148102
rect 291374 148046 291430 148102
rect 291498 148046 291554 148102
rect 291622 148046 291678 148102
rect 291250 147922 291306 147978
rect 291374 147922 291430 147978
rect 291498 147922 291554 147978
rect 291622 147922 291678 147978
rect 291250 130294 291306 130350
rect 291374 130294 291430 130350
rect 291498 130294 291554 130350
rect 291622 130294 291678 130350
rect 291250 130170 291306 130226
rect 291374 130170 291430 130226
rect 291498 130170 291554 130226
rect 291622 130170 291678 130226
rect 291250 130046 291306 130102
rect 291374 130046 291430 130102
rect 291498 130046 291554 130102
rect 291622 130046 291678 130102
rect 291250 129922 291306 129978
rect 291374 129922 291430 129978
rect 291498 129922 291554 129978
rect 291622 129922 291678 129978
rect 291250 112294 291306 112350
rect 291374 112294 291430 112350
rect 291498 112294 291554 112350
rect 291622 112294 291678 112350
rect 291250 112170 291306 112226
rect 291374 112170 291430 112226
rect 291498 112170 291554 112226
rect 291622 112170 291678 112226
rect 291250 112046 291306 112102
rect 291374 112046 291430 112102
rect 291498 112046 291554 112102
rect 291622 112046 291678 112102
rect 291250 111922 291306 111978
rect 291374 111922 291430 111978
rect 291498 111922 291554 111978
rect 291622 111922 291678 111978
rect 291250 94294 291306 94350
rect 291374 94294 291430 94350
rect 291498 94294 291554 94350
rect 291622 94294 291678 94350
rect 291250 94170 291306 94226
rect 291374 94170 291430 94226
rect 291498 94170 291554 94226
rect 291622 94170 291678 94226
rect 291250 94046 291306 94102
rect 291374 94046 291430 94102
rect 291498 94046 291554 94102
rect 291622 94046 291678 94102
rect 291250 93922 291306 93978
rect 291374 93922 291430 93978
rect 291498 93922 291554 93978
rect 291622 93922 291678 93978
rect 291250 76294 291306 76350
rect 291374 76294 291430 76350
rect 291498 76294 291554 76350
rect 291622 76294 291678 76350
rect 291250 76170 291306 76226
rect 291374 76170 291430 76226
rect 291498 76170 291554 76226
rect 291622 76170 291678 76226
rect 291250 76046 291306 76102
rect 291374 76046 291430 76102
rect 291498 76046 291554 76102
rect 291622 76046 291678 76102
rect 291250 75922 291306 75978
rect 291374 75922 291430 75978
rect 291498 75922 291554 75978
rect 291622 75922 291678 75978
rect 291250 58294 291306 58350
rect 291374 58294 291430 58350
rect 291498 58294 291554 58350
rect 291622 58294 291678 58350
rect 291250 58170 291306 58226
rect 291374 58170 291430 58226
rect 291498 58170 291554 58226
rect 291622 58170 291678 58226
rect 291250 58046 291306 58102
rect 291374 58046 291430 58102
rect 291498 58046 291554 58102
rect 291622 58046 291678 58102
rect 291250 57922 291306 57978
rect 291374 57922 291430 57978
rect 291498 57922 291554 57978
rect 291622 57922 291678 57978
rect 291250 40294 291306 40350
rect 291374 40294 291430 40350
rect 291498 40294 291554 40350
rect 291622 40294 291678 40350
rect 291250 40170 291306 40226
rect 291374 40170 291430 40226
rect 291498 40170 291554 40226
rect 291622 40170 291678 40226
rect 291250 40046 291306 40102
rect 291374 40046 291430 40102
rect 291498 40046 291554 40102
rect 291622 40046 291678 40102
rect 291250 39922 291306 39978
rect 291374 39922 291430 39978
rect 291498 39922 291554 39978
rect 291622 39922 291678 39978
rect 291250 22294 291306 22350
rect 291374 22294 291430 22350
rect 291498 22294 291554 22350
rect 291622 22294 291678 22350
rect 291250 22170 291306 22226
rect 291374 22170 291430 22226
rect 291498 22170 291554 22226
rect 291622 22170 291678 22226
rect 291250 22046 291306 22102
rect 291374 22046 291430 22102
rect 291498 22046 291554 22102
rect 291622 22046 291678 22102
rect 291250 21922 291306 21978
rect 291374 21922 291430 21978
rect 291498 21922 291554 21978
rect 291622 21922 291678 21978
rect 291250 4294 291306 4350
rect 291374 4294 291430 4350
rect 291498 4294 291554 4350
rect 291622 4294 291678 4350
rect 291250 4170 291306 4226
rect 291374 4170 291430 4226
rect 291498 4170 291554 4226
rect 291622 4170 291678 4226
rect 291250 4046 291306 4102
rect 291374 4046 291430 4102
rect 291498 4046 291554 4102
rect 291622 4046 291678 4102
rect 291250 3922 291306 3978
rect 291374 3922 291430 3978
rect 291498 3922 291554 3978
rect 291622 3922 291678 3978
rect 291250 -216 291306 -160
rect 291374 -216 291430 -160
rect 291498 -216 291554 -160
rect 291622 -216 291678 -160
rect 291250 -340 291306 -284
rect 291374 -340 291430 -284
rect 291498 -340 291554 -284
rect 291622 -340 291678 -284
rect 291250 -464 291306 -408
rect 291374 -464 291430 -408
rect 291498 -464 291554 -408
rect 291622 -464 291678 -408
rect 291250 -588 291306 -532
rect 291374 -588 291430 -532
rect 291498 -588 291554 -532
rect 291622 -588 291678 -532
rect 294970 208294 295026 208350
rect 295094 208294 295150 208350
rect 295218 208294 295274 208350
rect 295342 208294 295398 208350
rect 294970 208170 295026 208226
rect 295094 208170 295150 208226
rect 295218 208170 295274 208226
rect 295342 208170 295398 208226
rect 294970 208046 295026 208102
rect 295094 208046 295150 208102
rect 295218 208046 295274 208102
rect 295342 208046 295398 208102
rect 294970 207922 295026 207978
rect 295094 207922 295150 207978
rect 295218 207922 295274 207978
rect 295342 207922 295398 207978
rect 294970 190294 295026 190350
rect 295094 190294 295150 190350
rect 295218 190294 295274 190350
rect 295342 190294 295398 190350
rect 294970 190170 295026 190226
rect 295094 190170 295150 190226
rect 295218 190170 295274 190226
rect 295342 190170 295398 190226
rect 294970 190046 295026 190102
rect 295094 190046 295150 190102
rect 295218 190046 295274 190102
rect 295342 190046 295398 190102
rect 294970 189922 295026 189978
rect 295094 189922 295150 189978
rect 295218 189922 295274 189978
rect 295342 189922 295398 189978
rect 294970 172294 295026 172350
rect 295094 172294 295150 172350
rect 295218 172294 295274 172350
rect 295342 172294 295398 172350
rect 294970 172170 295026 172226
rect 295094 172170 295150 172226
rect 295218 172170 295274 172226
rect 295342 172170 295398 172226
rect 294970 172046 295026 172102
rect 295094 172046 295150 172102
rect 295218 172046 295274 172102
rect 295342 172046 295398 172102
rect 294970 171922 295026 171978
rect 295094 171922 295150 171978
rect 295218 171922 295274 171978
rect 295342 171922 295398 171978
rect 294970 154294 295026 154350
rect 295094 154294 295150 154350
rect 295218 154294 295274 154350
rect 295342 154294 295398 154350
rect 294970 154170 295026 154226
rect 295094 154170 295150 154226
rect 295218 154170 295274 154226
rect 295342 154170 295398 154226
rect 294970 154046 295026 154102
rect 295094 154046 295150 154102
rect 295218 154046 295274 154102
rect 295342 154046 295398 154102
rect 294970 153922 295026 153978
rect 295094 153922 295150 153978
rect 295218 153922 295274 153978
rect 295342 153922 295398 153978
rect 294970 136294 295026 136350
rect 295094 136294 295150 136350
rect 295218 136294 295274 136350
rect 295342 136294 295398 136350
rect 294970 136170 295026 136226
rect 295094 136170 295150 136226
rect 295218 136170 295274 136226
rect 295342 136170 295398 136226
rect 294970 136046 295026 136102
rect 295094 136046 295150 136102
rect 295218 136046 295274 136102
rect 295342 136046 295398 136102
rect 294970 135922 295026 135978
rect 295094 135922 295150 135978
rect 295218 135922 295274 135978
rect 295342 135922 295398 135978
rect 294970 118294 295026 118350
rect 295094 118294 295150 118350
rect 295218 118294 295274 118350
rect 295342 118294 295398 118350
rect 294970 118170 295026 118226
rect 295094 118170 295150 118226
rect 295218 118170 295274 118226
rect 295342 118170 295398 118226
rect 294970 118046 295026 118102
rect 295094 118046 295150 118102
rect 295218 118046 295274 118102
rect 295342 118046 295398 118102
rect 294970 117922 295026 117978
rect 295094 117922 295150 117978
rect 295218 117922 295274 117978
rect 295342 117922 295398 117978
rect 294970 100294 295026 100350
rect 295094 100294 295150 100350
rect 295218 100294 295274 100350
rect 295342 100294 295398 100350
rect 294970 100170 295026 100226
rect 295094 100170 295150 100226
rect 295218 100170 295274 100226
rect 295342 100170 295398 100226
rect 294970 100046 295026 100102
rect 295094 100046 295150 100102
rect 295218 100046 295274 100102
rect 295342 100046 295398 100102
rect 294970 99922 295026 99978
rect 295094 99922 295150 99978
rect 295218 99922 295274 99978
rect 295342 99922 295398 99978
rect 294970 82294 295026 82350
rect 295094 82294 295150 82350
rect 295218 82294 295274 82350
rect 295342 82294 295398 82350
rect 294970 82170 295026 82226
rect 295094 82170 295150 82226
rect 295218 82170 295274 82226
rect 295342 82170 295398 82226
rect 294970 82046 295026 82102
rect 295094 82046 295150 82102
rect 295218 82046 295274 82102
rect 295342 82046 295398 82102
rect 294970 81922 295026 81978
rect 295094 81922 295150 81978
rect 295218 81922 295274 81978
rect 295342 81922 295398 81978
rect 294970 64294 295026 64350
rect 295094 64294 295150 64350
rect 295218 64294 295274 64350
rect 295342 64294 295398 64350
rect 294970 64170 295026 64226
rect 295094 64170 295150 64226
rect 295218 64170 295274 64226
rect 295342 64170 295398 64226
rect 294970 64046 295026 64102
rect 295094 64046 295150 64102
rect 295218 64046 295274 64102
rect 295342 64046 295398 64102
rect 294970 63922 295026 63978
rect 295094 63922 295150 63978
rect 295218 63922 295274 63978
rect 295342 63922 295398 63978
rect 294970 46294 295026 46350
rect 295094 46294 295150 46350
rect 295218 46294 295274 46350
rect 295342 46294 295398 46350
rect 294970 46170 295026 46226
rect 295094 46170 295150 46226
rect 295218 46170 295274 46226
rect 295342 46170 295398 46226
rect 294970 46046 295026 46102
rect 295094 46046 295150 46102
rect 295218 46046 295274 46102
rect 295342 46046 295398 46102
rect 294970 45922 295026 45978
rect 295094 45922 295150 45978
rect 295218 45922 295274 45978
rect 295342 45922 295398 45978
rect 294970 28294 295026 28350
rect 295094 28294 295150 28350
rect 295218 28294 295274 28350
rect 295342 28294 295398 28350
rect 294970 28170 295026 28226
rect 295094 28170 295150 28226
rect 295218 28170 295274 28226
rect 295342 28170 295398 28226
rect 294970 28046 295026 28102
rect 295094 28046 295150 28102
rect 295218 28046 295274 28102
rect 295342 28046 295398 28102
rect 294970 27922 295026 27978
rect 295094 27922 295150 27978
rect 295218 27922 295274 27978
rect 295342 27922 295398 27978
rect 294970 10294 295026 10350
rect 295094 10294 295150 10350
rect 295218 10294 295274 10350
rect 295342 10294 295398 10350
rect 294970 10170 295026 10226
rect 295094 10170 295150 10226
rect 295218 10170 295274 10226
rect 295342 10170 295398 10226
rect 294970 10046 295026 10102
rect 295094 10046 295150 10102
rect 295218 10046 295274 10102
rect 295342 10046 295398 10102
rect 294970 9922 295026 9978
rect 295094 9922 295150 9978
rect 295218 9922 295274 9978
rect 295342 9922 295398 9978
rect 294970 -1176 295026 -1120
rect 295094 -1176 295150 -1120
rect 295218 -1176 295274 -1120
rect 295342 -1176 295398 -1120
rect 294970 -1300 295026 -1244
rect 295094 -1300 295150 -1244
rect 295218 -1300 295274 -1244
rect 295342 -1300 295398 -1244
rect 294970 -1424 295026 -1368
rect 295094 -1424 295150 -1368
rect 295218 -1424 295274 -1368
rect 295342 -1424 295398 -1368
rect 294970 -1548 295026 -1492
rect 295094 -1548 295150 -1492
rect 295218 -1548 295274 -1492
rect 295342 -1548 295398 -1492
rect 312038 208294 312094 208350
rect 312162 208294 312218 208350
rect 312038 208170 312094 208226
rect 312162 208170 312218 208226
rect 312038 208046 312094 208102
rect 312162 208046 312218 208102
rect 312038 207922 312094 207978
rect 312162 207922 312218 207978
rect 312970 208294 313026 208350
rect 313094 208294 313150 208350
rect 313218 208294 313274 208350
rect 313342 208294 313398 208350
rect 312970 208170 313026 208226
rect 313094 208170 313150 208226
rect 313218 208170 313274 208226
rect 313342 208170 313398 208226
rect 312970 208046 313026 208102
rect 313094 208046 313150 208102
rect 313218 208046 313274 208102
rect 313342 208046 313398 208102
rect 312970 207922 313026 207978
rect 313094 207922 313150 207978
rect 313218 207922 313274 207978
rect 313342 207922 313398 207978
rect 309250 202294 309306 202350
rect 309374 202294 309430 202350
rect 309498 202294 309554 202350
rect 309622 202294 309678 202350
rect 309250 202170 309306 202226
rect 309374 202170 309430 202226
rect 309498 202170 309554 202226
rect 309622 202170 309678 202226
rect 309250 202046 309306 202102
rect 309374 202046 309430 202102
rect 309498 202046 309554 202102
rect 309622 202046 309678 202102
rect 309250 201922 309306 201978
rect 309374 201922 309430 201978
rect 309498 201922 309554 201978
rect 309622 201922 309678 201978
rect 309250 184294 309306 184350
rect 309374 184294 309430 184350
rect 309498 184294 309554 184350
rect 309622 184294 309678 184350
rect 309250 184170 309306 184226
rect 309374 184170 309430 184226
rect 309498 184170 309554 184226
rect 309622 184170 309678 184226
rect 309250 184046 309306 184102
rect 309374 184046 309430 184102
rect 309498 184046 309554 184102
rect 309622 184046 309678 184102
rect 309250 183922 309306 183978
rect 309374 183922 309430 183978
rect 309498 183922 309554 183978
rect 309622 183922 309678 183978
rect 309250 166294 309306 166350
rect 309374 166294 309430 166350
rect 309498 166294 309554 166350
rect 309622 166294 309678 166350
rect 309250 166170 309306 166226
rect 309374 166170 309430 166226
rect 309498 166170 309554 166226
rect 309622 166170 309678 166226
rect 309250 166046 309306 166102
rect 309374 166046 309430 166102
rect 309498 166046 309554 166102
rect 309622 166046 309678 166102
rect 309250 165922 309306 165978
rect 309374 165922 309430 165978
rect 309498 165922 309554 165978
rect 309622 165922 309678 165978
rect 309250 148294 309306 148350
rect 309374 148294 309430 148350
rect 309498 148294 309554 148350
rect 309622 148294 309678 148350
rect 309250 148170 309306 148226
rect 309374 148170 309430 148226
rect 309498 148170 309554 148226
rect 309622 148170 309678 148226
rect 309250 148046 309306 148102
rect 309374 148046 309430 148102
rect 309498 148046 309554 148102
rect 309622 148046 309678 148102
rect 309250 147922 309306 147978
rect 309374 147922 309430 147978
rect 309498 147922 309554 147978
rect 309622 147922 309678 147978
rect 309250 130294 309306 130350
rect 309374 130294 309430 130350
rect 309498 130294 309554 130350
rect 309622 130294 309678 130350
rect 309250 130170 309306 130226
rect 309374 130170 309430 130226
rect 309498 130170 309554 130226
rect 309622 130170 309678 130226
rect 309250 130046 309306 130102
rect 309374 130046 309430 130102
rect 309498 130046 309554 130102
rect 309622 130046 309678 130102
rect 309250 129922 309306 129978
rect 309374 129922 309430 129978
rect 309498 129922 309554 129978
rect 309622 129922 309678 129978
rect 309250 112294 309306 112350
rect 309374 112294 309430 112350
rect 309498 112294 309554 112350
rect 309622 112294 309678 112350
rect 309250 112170 309306 112226
rect 309374 112170 309430 112226
rect 309498 112170 309554 112226
rect 309622 112170 309678 112226
rect 309250 112046 309306 112102
rect 309374 112046 309430 112102
rect 309498 112046 309554 112102
rect 309622 112046 309678 112102
rect 309250 111922 309306 111978
rect 309374 111922 309430 111978
rect 309498 111922 309554 111978
rect 309622 111922 309678 111978
rect 309250 94294 309306 94350
rect 309374 94294 309430 94350
rect 309498 94294 309554 94350
rect 309622 94294 309678 94350
rect 309250 94170 309306 94226
rect 309374 94170 309430 94226
rect 309498 94170 309554 94226
rect 309622 94170 309678 94226
rect 309250 94046 309306 94102
rect 309374 94046 309430 94102
rect 309498 94046 309554 94102
rect 309622 94046 309678 94102
rect 309250 93922 309306 93978
rect 309374 93922 309430 93978
rect 309498 93922 309554 93978
rect 309622 93922 309678 93978
rect 309250 76294 309306 76350
rect 309374 76294 309430 76350
rect 309498 76294 309554 76350
rect 309622 76294 309678 76350
rect 309250 76170 309306 76226
rect 309374 76170 309430 76226
rect 309498 76170 309554 76226
rect 309622 76170 309678 76226
rect 309250 76046 309306 76102
rect 309374 76046 309430 76102
rect 309498 76046 309554 76102
rect 309622 76046 309678 76102
rect 309250 75922 309306 75978
rect 309374 75922 309430 75978
rect 309498 75922 309554 75978
rect 309622 75922 309678 75978
rect 309250 58294 309306 58350
rect 309374 58294 309430 58350
rect 309498 58294 309554 58350
rect 309622 58294 309678 58350
rect 309250 58170 309306 58226
rect 309374 58170 309430 58226
rect 309498 58170 309554 58226
rect 309622 58170 309678 58226
rect 309250 58046 309306 58102
rect 309374 58046 309430 58102
rect 309498 58046 309554 58102
rect 309622 58046 309678 58102
rect 309250 57922 309306 57978
rect 309374 57922 309430 57978
rect 309498 57922 309554 57978
rect 309622 57922 309678 57978
rect 309250 40294 309306 40350
rect 309374 40294 309430 40350
rect 309498 40294 309554 40350
rect 309622 40294 309678 40350
rect 309250 40170 309306 40226
rect 309374 40170 309430 40226
rect 309498 40170 309554 40226
rect 309622 40170 309678 40226
rect 309250 40046 309306 40102
rect 309374 40046 309430 40102
rect 309498 40046 309554 40102
rect 309622 40046 309678 40102
rect 309250 39922 309306 39978
rect 309374 39922 309430 39978
rect 309498 39922 309554 39978
rect 309622 39922 309678 39978
rect 309250 22294 309306 22350
rect 309374 22294 309430 22350
rect 309498 22294 309554 22350
rect 309622 22294 309678 22350
rect 309250 22170 309306 22226
rect 309374 22170 309430 22226
rect 309498 22170 309554 22226
rect 309622 22170 309678 22226
rect 309250 22046 309306 22102
rect 309374 22046 309430 22102
rect 309498 22046 309554 22102
rect 309622 22046 309678 22102
rect 309250 21922 309306 21978
rect 309374 21922 309430 21978
rect 309498 21922 309554 21978
rect 309622 21922 309678 21978
rect 309250 4294 309306 4350
rect 309374 4294 309430 4350
rect 309498 4294 309554 4350
rect 309622 4294 309678 4350
rect 309250 4170 309306 4226
rect 309374 4170 309430 4226
rect 309498 4170 309554 4226
rect 309622 4170 309678 4226
rect 309250 4046 309306 4102
rect 309374 4046 309430 4102
rect 309498 4046 309554 4102
rect 309622 4046 309678 4102
rect 309250 3922 309306 3978
rect 309374 3922 309430 3978
rect 309498 3922 309554 3978
rect 309622 3922 309678 3978
rect 309250 -216 309306 -160
rect 309374 -216 309430 -160
rect 309498 -216 309554 -160
rect 309622 -216 309678 -160
rect 309250 -340 309306 -284
rect 309374 -340 309430 -284
rect 309498 -340 309554 -284
rect 309622 -340 309678 -284
rect 309250 -464 309306 -408
rect 309374 -464 309430 -408
rect 309498 -464 309554 -408
rect 309622 -464 309678 -408
rect 309250 -588 309306 -532
rect 309374 -588 309430 -532
rect 309498 -588 309554 -532
rect 309622 -588 309678 -532
rect 330970 208294 331026 208350
rect 331094 208294 331150 208350
rect 331218 208294 331274 208350
rect 331342 208294 331398 208350
rect 330970 208170 331026 208226
rect 331094 208170 331150 208226
rect 331218 208170 331274 208226
rect 331342 208170 331398 208226
rect 330970 208046 331026 208102
rect 331094 208046 331150 208102
rect 331218 208046 331274 208102
rect 331342 208046 331398 208102
rect 330970 207922 331026 207978
rect 331094 207922 331150 207978
rect 331218 207922 331274 207978
rect 331342 207922 331398 207978
rect 312970 190294 313026 190350
rect 313094 190294 313150 190350
rect 313218 190294 313274 190350
rect 313342 190294 313398 190350
rect 312970 190170 313026 190226
rect 313094 190170 313150 190226
rect 313218 190170 313274 190226
rect 313342 190170 313398 190226
rect 312970 190046 313026 190102
rect 313094 190046 313150 190102
rect 313218 190046 313274 190102
rect 313342 190046 313398 190102
rect 312970 189922 313026 189978
rect 313094 189922 313150 189978
rect 313218 189922 313274 189978
rect 313342 189922 313398 189978
rect 312970 172294 313026 172350
rect 313094 172294 313150 172350
rect 313218 172294 313274 172350
rect 313342 172294 313398 172350
rect 312970 172170 313026 172226
rect 313094 172170 313150 172226
rect 313218 172170 313274 172226
rect 313342 172170 313398 172226
rect 312970 172046 313026 172102
rect 313094 172046 313150 172102
rect 313218 172046 313274 172102
rect 313342 172046 313398 172102
rect 312970 171922 313026 171978
rect 313094 171922 313150 171978
rect 313218 171922 313274 171978
rect 313342 171922 313398 171978
rect 312970 154294 313026 154350
rect 313094 154294 313150 154350
rect 313218 154294 313274 154350
rect 313342 154294 313398 154350
rect 312970 154170 313026 154226
rect 313094 154170 313150 154226
rect 313218 154170 313274 154226
rect 313342 154170 313398 154226
rect 312970 154046 313026 154102
rect 313094 154046 313150 154102
rect 313218 154046 313274 154102
rect 313342 154046 313398 154102
rect 312970 153922 313026 153978
rect 313094 153922 313150 153978
rect 313218 153922 313274 153978
rect 313342 153922 313398 153978
rect 312970 136294 313026 136350
rect 313094 136294 313150 136350
rect 313218 136294 313274 136350
rect 313342 136294 313398 136350
rect 312970 136170 313026 136226
rect 313094 136170 313150 136226
rect 313218 136170 313274 136226
rect 313342 136170 313398 136226
rect 312970 136046 313026 136102
rect 313094 136046 313150 136102
rect 313218 136046 313274 136102
rect 313342 136046 313398 136102
rect 312970 135922 313026 135978
rect 313094 135922 313150 135978
rect 313218 135922 313274 135978
rect 313342 135922 313398 135978
rect 312970 118294 313026 118350
rect 313094 118294 313150 118350
rect 313218 118294 313274 118350
rect 313342 118294 313398 118350
rect 312970 118170 313026 118226
rect 313094 118170 313150 118226
rect 313218 118170 313274 118226
rect 313342 118170 313398 118226
rect 312970 118046 313026 118102
rect 313094 118046 313150 118102
rect 313218 118046 313274 118102
rect 313342 118046 313398 118102
rect 312970 117922 313026 117978
rect 313094 117922 313150 117978
rect 313218 117922 313274 117978
rect 313342 117922 313398 117978
rect 312970 100294 313026 100350
rect 313094 100294 313150 100350
rect 313218 100294 313274 100350
rect 313342 100294 313398 100350
rect 312970 100170 313026 100226
rect 313094 100170 313150 100226
rect 313218 100170 313274 100226
rect 313342 100170 313398 100226
rect 312970 100046 313026 100102
rect 313094 100046 313150 100102
rect 313218 100046 313274 100102
rect 313342 100046 313398 100102
rect 312970 99922 313026 99978
rect 313094 99922 313150 99978
rect 313218 99922 313274 99978
rect 313342 99922 313398 99978
rect 312970 82294 313026 82350
rect 313094 82294 313150 82350
rect 313218 82294 313274 82350
rect 313342 82294 313398 82350
rect 312970 82170 313026 82226
rect 313094 82170 313150 82226
rect 313218 82170 313274 82226
rect 313342 82170 313398 82226
rect 312970 82046 313026 82102
rect 313094 82046 313150 82102
rect 313218 82046 313274 82102
rect 313342 82046 313398 82102
rect 312970 81922 313026 81978
rect 313094 81922 313150 81978
rect 313218 81922 313274 81978
rect 313342 81922 313398 81978
rect 312970 64294 313026 64350
rect 313094 64294 313150 64350
rect 313218 64294 313274 64350
rect 313342 64294 313398 64350
rect 312970 64170 313026 64226
rect 313094 64170 313150 64226
rect 313218 64170 313274 64226
rect 313342 64170 313398 64226
rect 312970 64046 313026 64102
rect 313094 64046 313150 64102
rect 313218 64046 313274 64102
rect 313342 64046 313398 64102
rect 312970 63922 313026 63978
rect 313094 63922 313150 63978
rect 313218 63922 313274 63978
rect 313342 63922 313398 63978
rect 312970 46294 313026 46350
rect 313094 46294 313150 46350
rect 313218 46294 313274 46350
rect 313342 46294 313398 46350
rect 312970 46170 313026 46226
rect 313094 46170 313150 46226
rect 313218 46170 313274 46226
rect 313342 46170 313398 46226
rect 312970 46046 313026 46102
rect 313094 46046 313150 46102
rect 313218 46046 313274 46102
rect 313342 46046 313398 46102
rect 312970 45922 313026 45978
rect 313094 45922 313150 45978
rect 313218 45922 313274 45978
rect 313342 45922 313398 45978
rect 312970 28294 313026 28350
rect 313094 28294 313150 28350
rect 313218 28294 313274 28350
rect 313342 28294 313398 28350
rect 312970 28170 313026 28226
rect 313094 28170 313150 28226
rect 313218 28170 313274 28226
rect 313342 28170 313398 28226
rect 312970 28046 313026 28102
rect 313094 28046 313150 28102
rect 313218 28046 313274 28102
rect 313342 28046 313398 28102
rect 312970 27922 313026 27978
rect 313094 27922 313150 27978
rect 313218 27922 313274 27978
rect 313342 27922 313398 27978
rect 312970 10294 313026 10350
rect 313094 10294 313150 10350
rect 313218 10294 313274 10350
rect 313342 10294 313398 10350
rect 312970 10170 313026 10226
rect 313094 10170 313150 10226
rect 313218 10170 313274 10226
rect 313342 10170 313398 10226
rect 312970 10046 313026 10102
rect 313094 10046 313150 10102
rect 313218 10046 313274 10102
rect 313342 10046 313398 10102
rect 312970 9922 313026 9978
rect 313094 9922 313150 9978
rect 313218 9922 313274 9978
rect 313342 9922 313398 9978
rect 312970 -1176 313026 -1120
rect 313094 -1176 313150 -1120
rect 313218 -1176 313274 -1120
rect 313342 -1176 313398 -1120
rect 312970 -1300 313026 -1244
rect 313094 -1300 313150 -1244
rect 313218 -1300 313274 -1244
rect 313342 -1300 313398 -1244
rect 312970 -1424 313026 -1368
rect 313094 -1424 313150 -1368
rect 313218 -1424 313274 -1368
rect 313342 -1424 313398 -1368
rect 312970 -1548 313026 -1492
rect 313094 -1548 313150 -1492
rect 313218 -1548 313274 -1492
rect 313342 -1548 313398 -1492
rect 327250 184294 327306 184350
rect 327374 184294 327430 184350
rect 327498 184294 327554 184350
rect 327622 184294 327678 184350
rect 327250 184170 327306 184226
rect 327374 184170 327430 184226
rect 327498 184170 327554 184226
rect 327622 184170 327678 184226
rect 327250 184046 327306 184102
rect 327374 184046 327430 184102
rect 327498 184046 327554 184102
rect 327622 184046 327678 184102
rect 327250 183922 327306 183978
rect 327374 183922 327430 183978
rect 327498 183922 327554 183978
rect 327622 183922 327678 183978
rect 327250 166294 327306 166350
rect 327374 166294 327430 166350
rect 327498 166294 327554 166350
rect 327622 166294 327678 166350
rect 327250 166170 327306 166226
rect 327374 166170 327430 166226
rect 327498 166170 327554 166226
rect 327622 166170 327678 166226
rect 327250 166046 327306 166102
rect 327374 166046 327430 166102
rect 327498 166046 327554 166102
rect 327622 166046 327678 166102
rect 327250 165922 327306 165978
rect 327374 165922 327430 165978
rect 327498 165922 327554 165978
rect 327622 165922 327678 165978
rect 327250 148294 327306 148350
rect 327374 148294 327430 148350
rect 327498 148294 327554 148350
rect 327622 148294 327678 148350
rect 327250 148170 327306 148226
rect 327374 148170 327430 148226
rect 327498 148170 327554 148226
rect 327622 148170 327678 148226
rect 327250 148046 327306 148102
rect 327374 148046 327430 148102
rect 327498 148046 327554 148102
rect 327622 148046 327678 148102
rect 327250 147922 327306 147978
rect 327374 147922 327430 147978
rect 327498 147922 327554 147978
rect 327622 147922 327678 147978
rect 327250 130294 327306 130350
rect 327374 130294 327430 130350
rect 327498 130294 327554 130350
rect 327622 130294 327678 130350
rect 327250 130170 327306 130226
rect 327374 130170 327430 130226
rect 327498 130170 327554 130226
rect 327622 130170 327678 130226
rect 327250 130046 327306 130102
rect 327374 130046 327430 130102
rect 327498 130046 327554 130102
rect 327622 130046 327678 130102
rect 327250 129922 327306 129978
rect 327374 129922 327430 129978
rect 327498 129922 327554 129978
rect 327622 129922 327678 129978
rect 327250 112294 327306 112350
rect 327374 112294 327430 112350
rect 327498 112294 327554 112350
rect 327622 112294 327678 112350
rect 327250 112170 327306 112226
rect 327374 112170 327430 112226
rect 327498 112170 327554 112226
rect 327622 112170 327678 112226
rect 327250 112046 327306 112102
rect 327374 112046 327430 112102
rect 327498 112046 327554 112102
rect 327622 112046 327678 112102
rect 327250 111922 327306 111978
rect 327374 111922 327430 111978
rect 327498 111922 327554 111978
rect 327622 111922 327678 111978
rect 327250 94294 327306 94350
rect 327374 94294 327430 94350
rect 327498 94294 327554 94350
rect 327622 94294 327678 94350
rect 327250 94170 327306 94226
rect 327374 94170 327430 94226
rect 327498 94170 327554 94226
rect 327622 94170 327678 94226
rect 327250 94046 327306 94102
rect 327374 94046 327430 94102
rect 327498 94046 327554 94102
rect 327622 94046 327678 94102
rect 327250 93922 327306 93978
rect 327374 93922 327430 93978
rect 327498 93922 327554 93978
rect 327622 93922 327678 93978
rect 327250 76294 327306 76350
rect 327374 76294 327430 76350
rect 327498 76294 327554 76350
rect 327622 76294 327678 76350
rect 327250 76170 327306 76226
rect 327374 76170 327430 76226
rect 327498 76170 327554 76226
rect 327622 76170 327678 76226
rect 327250 76046 327306 76102
rect 327374 76046 327430 76102
rect 327498 76046 327554 76102
rect 327622 76046 327678 76102
rect 327250 75922 327306 75978
rect 327374 75922 327430 75978
rect 327498 75922 327554 75978
rect 327622 75922 327678 75978
rect 327250 58294 327306 58350
rect 327374 58294 327430 58350
rect 327498 58294 327554 58350
rect 327622 58294 327678 58350
rect 327250 58170 327306 58226
rect 327374 58170 327430 58226
rect 327498 58170 327554 58226
rect 327622 58170 327678 58226
rect 327250 58046 327306 58102
rect 327374 58046 327430 58102
rect 327498 58046 327554 58102
rect 327622 58046 327678 58102
rect 327250 57922 327306 57978
rect 327374 57922 327430 57978
rect 327498 57922 327554 57978
rect 327622 57922 327678 57978
rect 327250 40294 327306 40350
rect 327374 40294 327430 40350
rect 327498 40294 327554 40350
rect 327622 40294 327678 40350
rect 327250 40170 327306 40226
rect 327374 40170 327430 40226
rect 327498 40170 327554 40226
rect 327622 40170 327678 40226
rect 327250 40046 327306 40102
rect 327374 40046 327430 40102
rect 327498 40046 327554 40102
rect 327622 40046 327678 40102
rect 327250 39922 327306 39978
rect 327374 39922 327430 39978
rect 327498 39922 327554 39978
rect 327622 39922 327678 39978
rect 327250 22294 327306 22350
rect 327374 22294 327430 22350
rect 327498 22294 327554 22350
rect 327622 22294 327678 22350
rect 327250 22170 327306 22226
rect 327374 22170 327430 22226
rect 327498 22170 327554 22226
rect 327622 22170 327678 22226
rect 327250 22046 327306 22102
rect 327374 22046 327430 22102
rect 327498 22046 327554 22102
rect 327622 22046 327678 22102
rect 327250 21922 327306 21978
rect 327374 21922 327430 21978
rect 327498 21922 327554 21978
rect 327622 21922 327678 21978
rect 327250 4294 327306 4350
rect 327374 4294 327430 4350
rect 327498 4294 327554 4350
rect 327622 4294 327678 4350
rect 327250 4170 327306 4226
rect 327374 4170 327430 4226
rect 327498 4170 327554 4226
rect 327622 4170 327678 4226
rect 327250 4046 327306 4102
rect 327374 4046 327430 4102
rect 327498 4046 327554 4102
rect 327622 4046 327678 4102
rect 327250 3922 327306 3978
rect 327374 3922 327430 3978
rect 327498 3922 327554 3978
rect 327622 3922 327678 3978
rect 327250 -216 327306 -160
rect 327374 -216 327430 -160
rect 327498 -216 327554 -160
rect 327622 -216 327678 -160
rect 327250 -340 327306 -284
rect 327374 -340 327430 -284
rect 327498 -340 327554 -284
rect 327622 -340 327678 -284
rect 327250 -464 327306 -408
rect 327374 -464 327430 -408
rect 327498 -464 327554 -408
rect 327622 -464 327678 -408
rect 327250 -588 327306 -532
rect 327374 -588 327430 -532
rect 327498 -588 327554 -532
rect 327622 -588 327678 -532
rect 342758 208294 342814 208350
rect 342882 208294 342938 208350
rect 342758 208170 342814 208226
rect 342882 208170 342938 208226
rect 342758 208046 342814 208102
rect 342882 208046 342938 208102
rect 342758 207922 342814 207978
rect 342882 207922 342938 207978
rect 330970 190294 331026 190350
rect 331094 190294 331150 190350
rect 331218 190294 331274 190350
rect 331342 190294 331398 190350
rect 330970 190170 331026 190226
rect 331094 190170 331150 190226
rect 331218 190170 331274 190226
rect 331342 190170 331398 190226
rect 330970 190046 331026 190102
rect 331094 190046 331150 190102
rect 331218 190046 331274 190102
rect 331342 190046 331398 190102
rect 330970 189922 331026 189978
rect 331094 189922 331150 189978
rect 331218 189922 331274 189978
rect 331342 189922 331398 189978
rect 330970 172294 331026 172350
rect 331094 172294 331150 172350
rect 331218 172294 331274 172350
rect 331342 172294 331398 172350
rect 330970 172170 331026 172226
rect 331094 172170 331150 172226
rect 331218 172170 331274 172226
rect 331342 172170 331398 172226
rect 330970 172046 331026 172102
rect 331094 172046 331150 172102
rect 331218 172046 331274 172102
rect 331342 172046 331398 172102
rect 330970 171922 331026 171978
rect 331094 171922 331150 171978
rect 331218 171922 331274 171978
rect 331342 171922 331398 171978
rect 330970 154294 331026 154350
rect 331094 154294 331150 154350
rect 331218 154294 331274 154350
rect 331342 154294 331398 154350
rect 330970 154170 331026 154226
rect 331094 154170 331150 154226
rect 331218 154170 331274 154226
rect 331342 154170 331398 154226
rect 330970 154046 331026 154102
rect 331094 154046 331150 154102
rect 331218 154046 331274 154102
rect 331342 154046 331398 154102
rect 330970 153922 331026 153978
rect 331094 153922 331150 153978
rect 331218 153922 331274 153978
rect 331342 153922 331398 153978
rect 330970 136294 331026 136350
rect 331094 136294 331150 136350
rect 331218 136294 331274 136350
rect 331342 136294 331398 136350
rect 330970 136170 331026 136226
rect 331094 136170 331150 136226
rect 331218 136170 331274 136226
rect 331342 136170 331398 136226
rect 330970 136046 331026 136102
rect 331094 136046 331150 136102
rect 331218 136046 331274 136102
rect 331342 136046 331398 136102
rect 330970 135922 331026 135978
rect 331094 135922 331150 135978
rect 331218 135922 331274 135978
rect 331342 135922 331398 135978
rect 330970 118294 331026 118350
rect 331094 118294 331150 118350
rect 331218 118294 331274 118350
rect 331342 118294 331398 118350
rect 330970 118170 331026 118226
rect 331094 118170 331150 118226
rect 331218 118170 331274 118226
rect 331342 118170 331398 118226
rect 330970 118046 331026 118102
rect 331094 118046 331150 118102
rect 331218 118046 331274 118102
rect 331342 118046 331398 118102
rect 330970 117922 331026 117978
rect 331094 117922 331150 117978
rect 331218 117922 331274 117978
rect 331342 117922 331398 117978
rect 330970 100294 331026 100350
rect 331094 100294 331150 100350
rect 331218 100294 331274 100350
rect 331342 100294 331398 100350
rect 330970 100170 331026 100226
rect 331094 100170 331150 100226
rect 331218 100170 331274 100226
rect 331342 100170 331398 100226
rect 330970 100046 331026 100102
rect 331094 100046 331150 100102
rect 331218 100046 331274 100102
rect 331342 100046 331398 100102
rect 330970 99922 331026 99978
rect 331094 99922 331150 99978
rect 331218 99922 331274 99978
rect 331342 99922 331398 99978
rect 330970 82294 331026 82350
rect 331094 82294 331150 82350
rect 331218 82294 331274 82350
rect 331342 82294 331398 82350
rect 330970 82170 331026 82226
rect 331094 82170 331150 82226
rect 331218 82170 331274 82226
rect 331342 82170 331398 82226
rect 330970 82046 331026 82102
rect 331094 82046 331150 82102
rect 331218 82046 331274 82102
rect 331342 82046 331398 82102
rect 330970 81922 331026 81978
rect 331094 81922 331150 81978
rect 331218 81922 331274 81978
rect 331342 81922 331398 81978
rect 330970 64294 331026 64350
rect 331094 64294 331150 64350
rect 331218 64294 331274 64350
rect 331342 64294 331398 64350
rect 330970 64170 331026 64226
rect 331094 64170 331150 64226
rect 331218 64170 331274 64226
rect 331342 64170 331398 64226
rect 330970 64046 331026 64102
rect 331094 64046 331150 64102
rect 331218 64046 331274 64102
rect 331342 64046 331398 64102
rect 330970 63922 331026 63978
rect 331094 63922 331150 63978
rect 331218 63922 331274 63978
rect 331342 63922 331398 63978
rect 330970 46294 331026 46350
rect 331094 46294 331150 46350
rect 331218 46294 331274 46350
rect 331342 46294 331398 46350
rect 330970 46170 331026 46226
rect 331094 46170 331150 46226
rect 331218 46170 331274 46226
rect 331342 46170 331398 46226
rect 330970 46046 331026 46102
rect 331094 46046 331150 46102
rect 331218 46046 331274 46102
rect 331342 46046 331398 46102
rect 330970 45922 331026 45978
rect 331094 45922 331150 45978
rect 331218 45922 331274 45978
rect 331342 45922 331398 45978
rect 330970 28294 331026 28350
rect 331094 28294 331150 28350
rect 331218 28294 331274 28350
rect 331342 28294 331398 28350
rect 330970 28170 331026 28226
rect 331094 28170 331150 28226
rect 331218 28170 331274 28226
rect 331342 28170 331398 28226
rect 330970 28046 331026 28102
rect 331094 28046 331150 28102
rect 331218 28046 331274 28102
rect 331342 28046 331398 28102
rect 330970 27922 331026 27978
rect 331094 27922 331150 27978
rect 331218 27922 331274 27978
rect 331342 27922 331398 27978
rect 330970 10294 331026 10350
rect 331094 10294 331150 10350
rect 331218 10294 331274 10350
rect 331342 10294 331398 10350
rect 330970 10170 331026 10226
rect 331094 10170 331150 10226
rect 331218 10170 331274 10226
rect 331342 10170 331398 10226
rect 330970 10046 331026 10102
rect 331094 10046 331150 10102
rect 331218 10046 331274 10102
rect 331342 10046 331398 10102
rect 330970 9922 331026 9978
rect 331094 9922 331150 9978
rect 331218 9922 331274 9978
rect 331342 9922 331398 9978
rect 330970 -1176 331026 -1120
rect 331094 -1176 331150 -1120
rect 331218 -1176 331274 -1120
rect 331342 -1176 331398 -1120
rect 330970 -1300 331026 -1244
rect 331094 -1300 331150 -1244
rect 331218 -1300 331274 -1244
rect 331342 -1300 331398 -1244
rect 330970 -1424 331026 -1368
rect 331094 -1424 331150 -1368
rect 331218 -1424 331274 -1368
rect 331342 -1424 331398 -1368
rect 330970 -1548 331026 -1492
rect 331094 -1548 331150 -1492
rect 331218 -1548 331274 -1492
rect 331342 -1548 331398 -1492
rect 345250 202294 345306 202350
rect 345374 202294 345430 202350
rect 345498 202294 345554 202350
rect 345622 202294 345678 202350
rect 345250 202170 345306 202226
rect 345374 202170 345430 202226
rect 345498 202170 345554 202226
rect 345622 202170 345678 202226
rect 345250 202046 345306 202102
rect 345374 202046 345430 202102
rect 345498 202046 345554 202102
rect 345622 202046 345678 202102
rect 345250 201922 345306 201978
rect 345374 201922 345430 201978
rect 345498 201922 345554 201978
rect 345622 201922 345678 201978
rect 345250 184294 345306 184350
rect 345374 184294 345430 184350
rect 345498 184294 345554 184350
rect 345622 184294 345678 184350
rect 345250 184170 345306 184226
rect 345374 184170 345430 184226
rect 345498 184170 345554 184226
rect 345622 184170 345678 184226
rect 345250 184046 345306 184102
rect 345374 184046 345430 184102
rect 345498 184046 345554 184102
rect 345622 184046 345678 184102
rect 345250 183922 345306 183978
rect 345374 183922 345430 183978
rect 345498 183922 345554 183978
rect 345622 183922 345678 183978
rect 345250 166294 345306 166350
rect 345374 166294 345430 166350
rect 345498 166294 345554 166350
rect 345622 166294 345678 166350
rect 345250 166170 345306 166226
rect 345374 166170 345430 166226
rect 345498 166170 345554 166226
rect 345622 166170 345678 166226
rect 345250 166046 345306 166102
rect 345374 166046 345430 166102
rect 345498 166046 345554 166102
rect 345622 166046 345678 166102
rect 345250 165922 345306 165978
rect 345374 165922 345430 165978
rect 345498 165922 345554 165978
rect 345622 165922 345678 165978
rect 345250 148294 345306 148350
rect 345374 148294 345430 148350
rect 345498 148294 345554 148350
rect 345622 148294 345678 148350
rect 345250 148170 345306 148226
rect 345374 148170 345430 148226
rect 345498 148170 345554 148226
rect 345622 148170 345678 148226
rect 345250 148046 345306 148102
rect 345374 148046 345430 148102
rect 345498 148046 345554 148102
rect 345622 148046 345678 148102
rect 345250 147922 345306 147978
rect 345374 147922 345430 147978
rect 345498 147922 345554 147978
rect 345622 147922 345678 147978
rect 345250 130294 345306 130350
rect 345374 130294 345430 130350
rect 345498 130294 345554 130350
rect 345622 130294 345678 130350
rect 345250 130170 345306 130226
rect 345374 130170 345430 130226
rect 345498 130170 345554 130226
rect 345622 130170 345678 130226
rect 345250 130046 345306 130102
rect 345374 130046 345430 130102
rect 345498 130046 345554 130102
rect 345622 130046 345678 130102
rect 345250 129922 345306 129978
rect 345374 129922 345430 129978
rect 345498 129922 345554 129978
rect 345622 129922 345678 129978
rect 345250 112294 345306 112350
rect 345374 112294 345430 112350
rect 345498 112294 345554 112350
rect 345622 112294 345678 112350
rect 345250 112170 345306 112226
rect 345374 112170 345430 112226
rect 345498 112170 345554 112226
rect 345622 112170 345678 112226
rect 345250 112046 345306 112102
rect 345374 112046 345430 112102
rect 345498 112046 345554 112102
rect 345622 112046 345678 112102
rect 345250 111922 345306 111978
rect 345374 111922 345430 111978
rect 345498 111922 345554 111978
rect 345622 111922 345678 111978
rect 345250 94294 345306 94350
rect 345374 94294 345430 94350
rect 345498 94294 345554 94350
rect 345622 94294 345678 94350
rect 345250 94170 345306 94226
rect 345374 94170 345430 94226
rect 345498 94170 345554 94226
rect 345622 94170 345678 94226
rect 345250 94046 345306 94102
rect 345374 94046 345430 94102
rect 345498 94046 345554 94102
rect 345622 94046 345678 94102
rect 345250 93922 345306 93978
rect 345374 93922 345430 93978
rect 345498 93922 345554 93978
rect 345622 93922 345678 93978
rect 345250 76294 345306 76350
rect 345374 76294 345430 76350
rect 345498 76294 345554 76350
rect 345622 76294 345678 76350
rect 345250 76170 345306 76226
rect 345374 76170 345430 76226
rect 345498 76170 345554 76226
rect 345622 76170 345678 76226
rect 345250 76046 345306 76102
rect 345374 76046 345430 76102
rect 345498 76046 345554 76102
rect 345622 76046 345678 76102
rect 345250 75922 345306 75978
rect 345374 75922 345430 75978
rect 345498 75922 345554 75978
rect 345622 75922 345678 75978
rect 345250 58294 345306 58350
rect 345374 58294 345430 58350
rect 345498 58294 345554 58350
rect 345622 58294 345678 58350
rect 345250 58170 345306 58226
rect 345374 58170 345430 58226
rect 345498 58170 345554 58226
rect 345622 58170 345678 58226
rect 345250 58046 345306 58102
rect 345374 58046 345430 58102
rect 345498 58046 345554 58102
rect 345622 58046 345678 58102
rect 345250 57922 345306 57978
rect 345374 57922 345430 57978
rect 345498 57922 345554 57978
rect 345622 57922 345678 57978
rect 345250 40294 345306 40350
rect 345374 40294 345430 40350
rect 345498 40294 345554 40350
rect 345622 40294 345678 40350
rect 345250 40170 345306 40226
rect 345374 40170 345430 40226
rect 345498 40170 345554 40226
rect 345622 40170 345678 40226
rect 345250 40046 345306 40102
rect 345374 40046 345430 40102
rect 345498 40046 345554 40102
rect 345622 40046 345678 40102
rect 345250 39922 345306 39978
rect 345374 39922 345430 39978
rect 345498 39922 345554 39978
rect 345622 39922 345678 39978
rect 345250 22294 345306 22350
rect 345374 22294 345430 22350
rect 345498 22294 345554 22350
rect 345622 22294 345678 22350
rect 345250 22170 345306 22226
rect 345374 22170 345430 22226
rect 345498 22170 345554 22226
rect 345622 22170 345678 22226
rect 345250 22046 345306 22102
rect 345374 22046 345430 22102
rect 345498 22046 345554 22102
rect 345622 22046 345678 22102
rect 345250 21922 345306 21978
rect 345374 21922 345430 21978
rect 345498 21922 345554 21978
rect 345622 21922 345678 21978
rect 345250 4294 345306 4350
rect 345374 4294 345430 4350
rect 345498 4294 345554 4350
rect 345622 4294 345678 4350
rect 345250 4170 345306 4226
rect 345374 4170 345430 4226
rect 345498 4170 345554 4226
rect 345622 4170 345678 4226
rect 345250 4046 345306 4102
rect 345374 4046 345430 4102
rect 345498 4046 345554 4102
rect 345622 4046 345678 4102
rect 345250 3922 345306 3978
rect 345374 3922 345430 3978
rect 345498 3922 345554 3978
rect 345622 3922 345678 3978
rect 345250 -216 345306 -160
rect 345374 -216 345430 -160
rect 345498 -216 345554 -160
rect 345622 -216 345678 -160
rect 345250 -340 345306 -284
rect 345374 -340 345430 -284
rect 345498 -340 345554 -284
rect 345622 -340 345678 -284
rect 345250 -464 345306 -408
rect 345374 -464 345430 -408
rect 345498 -464 345554 -408
rect 345622 -464 345678 -408
rect 345250 -588 345306 -532
rect 345374 -588 345430 -532
rect 345498 -588 345554 -532
rect 345622 -588 345678 -532
rect 348970 208294 349026 208350
rect 349094 208294 349150 208350
rect 349218 208294 349274 208350
rect 349342 208294 349398 208350
rect 348970 208170 349026 208226
rect 349094 208170 349150 208226
rect 349218 208170 349274 208226
rect 349342 208170 349398 208226
rect 348970 208046 349026 208102
rect 349094 208046 349150 208102
rect 349218 208046 349274 208102
rect 349342 208046 349398 208102
rect 348970 207922 349026 207978
rect 349094 207922 349150 207978
rect 349218 207922 349274 207978
rect 349342 207922 349398 207978
rect 348970 190294 349026 190350
rect 349094 190294 349150 190350
rect 349218 190294 349274 190350
rect 349342 190294 349398 190350
rect 348970 190170 349026 190226
rect 349094 190170 349150 190226
rect 349218 190170 349274 190226
rect 349342 190170 349398 190226
rect 348970 190046 349026 190102
rect 349094 190046 349150 190102
rect 349218 190046 349274 190102
rect 349342 190046 349398 190102
rect 348970 189922 349026 189978
rect 349094 189922 349150 189978
rect 349218 189922 349274 189978
rect 349342 189922 349398 189978
rect 348970 172294 349026 172350
rect 349094 172294 349150 172350
rect 349218 172294 349274 172350
rect 349342 172294 349398 172350
rect 348970 172170 349026 172226
rect 349094 172170 349150 172226
rect 349218 172170 349274 172226
rect 349342 172170 349398 172226
rect 348970 172046 349026 172102
rect 349094 172046 349150 172102
rect 349218 172046 349274 172102
rect 349342 172046 349398 172102
rect 348970 171922 349026 171978
rect 349094 171922 349150 171978
rect 349218 171922 349274 171978
rect 349342 171922 349398 171978
rect 348970 154294 349026 154350
rect 349094 154294 349150 154350
rect 349218 154294 349274 154350
rect 349342 154294 349398 154350
rect 348970 154170 349026 154226
rect 349094 154170 349150 154226
rect 349218 154170 349274 154226
rect 349342 154170 349398 154226
rect 348970 154046 349026 154102
rect 349094 154046 349150 154102
rect 349218 154046 349274 154102
rect 349342 154046 349398 154102
rect 348970 153922 349026 153978
rect 349094 153922 349150 153978
rect 349218 153922 349274 153978
rect 349342 153922 349398 153978
rect 348970 136294 349026 136350
rect 349094 136294 349150 136350
rect 349218 136294 349274 136350
rect 349342 136294 349398 136350
rect 348970 136170 349026 136226
rect 349094 136170 349150 136226
rect 349218 136170 349274 136226
rect 349342 136170 349398 136226
rect 348970 136046 349026 136102
rect 349094 136046 349150 136102
rect 349218 136046 349274 136102
rect 349342 136046 349398 136102
rect 348970 135922 349026 135978
rect 349094 135922 349150 135978
rect 349218 135922 349274 135978
rect 349342 135922 349398 135978
rect 348970 118294 349026 118350
rect 349094 118294 349150 118350
rect 349218 118294 349274 118350
rect 349342 118294 349398 118350
rect 348970 118170 349026 118226
rect 349094 118170 349150 118226
rect 349218 118170 349274 118226
rect 349342 118170 349398 118226
rect 348970 118046 349026 118102
rect 349094 118046 349150 118102
rect 349218 118046 349274 118102
rect 349342 118046 349398 118102
rect 348970 117922 349026 117978
rect 349094 117922 349150 117978
rect 349218 117922 349274 117978
rect 349342 117922 349398 117978
rect 348970 100294 349026 100350
rect 349094 100294 349150 100350
rect 349218 100294 349274 100350
rect 349342 100294 349398 100350
rect 348970 100170 349026 100226
rect 349094 100170 349150 100226
rect 349218 100170 349274 100226
rect 349342 100170 349398 100226
rect 348970 100046 349026 100102
rect 349094 100046 349150 100102
rect 349218 100046 349274 100102
rect 349342 100046 349398 100102
rect 348970 99922 349026 99978
rect 349094 99922 349150 99978
rect 349218 99922 349274 99978
rect 349342 99922 349398 99978
rect 348970 82294 349026 82350
rect 349094 82294 349150 82350
rect 349218 82294 349274 82350
rect 349342 82294 349398 82350
rect 348970 82170 349026 82226
rect 349094 82170 349150 82226
rect 349218 82170 349274 82226
rect 349342 82170 349398 82226
rect 348970 82046 349026 82102
rect 349094 82046 349150 82102
rect 349218 82046 349274 82102
rect 349342 82046 349398 82102
rect 348970 81922 349026 81978
rect 349094 81922 349150 81978
rect 349218 81922 349274 81978
rect 349342 81922 349398 81978
rect 348970 64294 349026 64350
rect 349094 64294 349150 64350
rect 349218 64294 349274 64350
rect 349342 64294 349398 64350
rect 348970 64170 349026 64226
rect 349094 64170 349150 64226
rect 349218 64170 349274 64226
rect 349342 64170 349398 64226
rect 348970 64046 349026 64102
rect 349094 64046 349150 64102
rect 349218 64046 349274 64102
rect 349342 64046 349398 64102
rect 348970 63922 349026 63978
rect 349094 63922 349150 63978
rect 349218 63922 349274 63978
rect 349342 63922 349398 63978
rect 348970 46294 349026 46350
rect 349094 46294 349150 46350
rect 349218 46294 349274 46350
rect 349342 46294 349398 46350
rect 348970 46170 349026 46226
rect 349094 46170 349150 46226
rect 349218 46170 349274 46226
rect 349342 46170 349398 46226
rect 348970 46046 349026 46102
rect 349094 46046 349150 46102
rect 349218 46046 349274 46102
rect 349342 46046 349398 46102
rect 348970 45922 349026 45978
rect 349094 45922 349150 45978
rect 349218 45922 349274 45978
rect 349342 45922 349398 45978
rect 348970 28294 349026 28350
rect 349094 28294 349150 28350
rect 349218 28294 349274 28350
rect 349342 28294 349398 28350
rect 348970 28170 349026 28226
rect 349094 28170 349150 28226
rect 349218 28170 349274 28226
rect 349342 28170 349398 28226
rect 348970 28046 349026 28102
rect 349094 28046 349150 28102
rect 349218 28046 349274 28102
rect 349342 28046 349398 28102
rect 348970 27922 349026 27978
rect 349094 27922 349150 27978
rect 349218 27922 349274 27978
rect 349342 27922 349398 27978
rect 348970 10294 349026 10350
rect 349094 10294 349150 10350
rect 349218 10294 349274 10350
rect 349342 10294 349398 10350
rect 348970 10170 349026 10226
rect 349094 10170 349150 10226
rect 349218 10170 349274 10226
rect 349342 10170 349398 10226
rect 348970 10046 349026 10102
rect 349094 10046 349150 10102
rect 349218 10046 349274 10102
rect 349342 10046 349398 10102
rect 348970 9922 349026 9978
rect 349094 9922 349150 9978
rect 349218 9922 349274 9978
rect 349342 9922 349398 9978
rect 348970 -1176 349026 -1120
rect 349094 -1176 349150 -1120
rect 349218 -1176 349274 -1120
rect 349342 -1176 349398 -1120
rect 348970 -1300 349026 -1244
rect 349094 -1300 349150 -1244
rect 349218 -1300 349274 -1244
rect 349342 -1300 349398 -1244
rect 348970 -1424 349026 -1368
rect 349094 -1424 349150 -1368
rect 349218 -1424 349274 -1368
rect 349342 -1424 349398 -1368
rect 348970 -1548 349026 -1492
rect 349094 -1548 349150 -1492
rect 349218 -1548 349274 -1492
rect 349342 -1548 349398 -1492
rect 363250 202294 363306 202350
rect 363374 202294 363430 202350
rect 363498 202294 363554 202350
rect 363622 202294 363678 202350
rect 363250 202170 363306 202226
rect 363374 202170 363430 202226
rect 363498 202170 363554 202226
rect 363622 202170 363678 202226
rect 363250 202046 363306 202102
rect 363374 202046 363430 202102
rect 363498 202046 363554 202102
rect 363622 202046 363678 202102
rect 363250 201922 363306 201978
rect 363374 201922 363430 201978
rect 363498 201922 363554 201978
rect 363622 201922 363678 201978
rect 363250 184294 363306 184350
rect 363374 184294 363430 184350
rect 363498 184294 363554 184350
rect 363622 184294 363678 184350
rect 363250 184170 363306 184226
rect 363374 184170 363430 184226
rect 363498 184170 363554 184226
rect 363622 184170 363678 184226
rect 363250 184046 363306 184102
rect 363374 184046 363430 184102
rect 363498 184046 363554 184102
rect 363622 184046 363678 184102
rect 363250 183922 363306 183978
rect 363374 183922 363430 183978
rect 363498 183922 363554 183978
rect 363622 183922 363678 183978
rect 363250 166294 363306 166350
rect 363374 166294 363430 166350
rect 363498 166294 363554 166350
rect 363622 166294 363678 166350
rect 363250 166170 363306 166226
rect 363374 166170 363430 166226
rect 363498 166170 363554 166226
rect 363622 166170 363678 166226
rect 363250 166046 363306 166102
rect 363374 166046 363430 166102
rect 363498 166046 363554 166102
rect 363622 166046 363678 166102
rect 363250 165922 363306 165978
rect 363374 165922 363430 165978
rect 363498 165922 363554 165978
rect 363622 165922 363678 165978
rect 363250 148294 363306 148350
rect 363374 148294 363430 148350
rect 363498 148294 363554 148350
rect 363622 148294 363678 148350
rect 363250 148170 363306 148226
rect 363374 148170 363430 148226
rect 363498 148170 363554 148226
rect 363622 148170 363678 148226
rect 363250 148046 363306 148102
rect 363374 148046 363430 148102
rect 363498 148046 363554 148102
rect 363622 148046 363678 148102
rect 363250 147922 363306 147978
rect 363374 147922 363430 147978
rect 363498 147922 363554 147978
rect 363622 147922 363678 147978
rect 363250 130294 363306 130350
rect 363374 130294 363430 130350
rect 363498 130294 363554 130350
rect 363622 130294 363678 130350
rect 363250 130170 363306 130226
rect 363374 130170 363430 130226
rect 363498 130170 363554 130226
rect 363622 130170 363678 130226
rect 363250 130046 363306 130102
rect 363374 130046 363430 130102
rect 363498 130046 363554 130102
rect 363622 130046 363678 130102
rect 363250 129922 363306 129978
rect 363374 129922 363430 129978
rect 363498 129922 363554 129978
rect 363622 129922 363678 129978
rect 363250 112294 363306 112350
rect 363374 112294 363430 112350
rect 363498 112294 363554 112350
rect 363622 112294 363678 112350
rect 363250 112170 363306 112226
rect 363374 112170 363430 112226
rect 363498 112170 363554 112226
rect 363622 112170 363678 112226
rect 363250 112046 363306 112102
rect 363374 112046 363430 112102
rect 363498 112046 363554 112102
rect 363622 112046 363678 112102
rect 363250 111922 363306 111978
rect 363374 111922 363430 111978
rect 363498 111922 363554 111978
rect 363622 111922 363678 111978
rect 363250 94294 363306 94350
rect 363374 94294 363430 94350
rect 363498 94294 363554 94350
rect 363622 94294 363678 94350
rect 363250 94170 363306 94226
rect 363374 94170 363430 94226
rect 363498 94170 363554 94226
rect 363622 94170 363678 94226
rect 363250 94046 363306 94102
rect 363374 94046 363430 94102
rect 363498 94046 363554 94102
rect 363622 94046 363678 94102
rect 363250 93922 363306 93978
rect 363374 93922 363430 93978
rect 363498 93922 363554 93978
rect 363622 93922 363678 93978
rect 363250 76294 363306 76350
rect 363374 76294 363430 76350
rect 363498 76294 363554 76350
rect 363622 76294 363678 76350
rect 363250 76170 363306 76226
rect 363374 76170 363430 76226
rect 363498 76170 363554 76226
rect 363622 76170 363678 76226
rect 363250 76046 363306 76102
rect 363374 76046 363430 76102
rect 363498 76046 363554 76102
rect 363622 76046 363678 76102
rect 363250 75922 363306 75978
rect 363374 75922 363430 75978
rect 363498 75922 363554 75978
rect 363622 75922 363678 75978
rect 363250 58294 363306 58350
rect 363374 58294 363430 58350
rect 363498 58294 363554 58350
rect 363622 58294 363678 58350
rect 363250 58170 363306 58226
rect 363374 58170 363430 58226
rect 363498 58170 363554 58226
rect 363622 58170 363678 58226
rect 363250 58046 363306 58102
rect 363374 58046 363430 58102
rect 363498 58046 363554 58102
rect 363622 58046 363678 58102
rect 363250 57922 363306 57978
rect 363374 57922 363430 57978
rect 363498 57922 363554 57978
rect 363622 57922 363678 57978
rect 363250 40294 363306 40350
rect 363374 40294 363430 40350
rect 363498 40294 363554 40350
rect 363622 40294 363678 40350
rect 363250 40170 363306 40226
rect 363374 40170 363430 40226
rect 363498 40170 363554 40226
rect 363622 40170 363678 40226
rect 363250 40046 363306 40102
rect 363374 40046 363430 40102
rect 363498 40046 363554 40102
rect 363622 40046 363678 40102
rect 363250 39922 363306 39978
rect 363374 39922 363430 39978
rect 363498 39922 363554 39978
rect 363622 39922 363678 39978
rect 363250 22294 363306 22350
rect 363374 22294 363430 22350
rect 363498 22294 363554 22350
rect 363622 22294 363678 22350
rect 363250 22170 363306 22226
rect 363374 22170 363430 22226
rect 363498 22170 363554 22226
rect 363622 22170 363678 22226
rect 363250 22046 363306 22102
rect 363374 22046 363430 22102
rect 363498 22046 363554 22102
rect 363622 22046 363678 22102
rect 363250 21922 363306 21978
rect 363374 21922 363430 21978
rect 363498 21922 363554 21978
rect 363622 21922 363678 21978
rect 363250 4294 363306 4350
rect 363374 4294 363430 4350
rect 363498 4294 363554 4350
rect 363622 4294 363678 4350
rect 363250 4170 363306 4226
rect 363374 4170 363430 4226
rect 363498 4170 363554 4226
rect 363622 4170 363678 4226
rect 363250 4046 363306 4102
rect 363374 4046 363430 4102
rect 363498 4046 363554 4102
rect 363622 4046 363678 4102
rect 363250 3922 363306 3978
rect 363374 3922 363430 3978
rect 363498 3922 363554 3978
rect 363622 3922 363678 3978
rect 363250 -216 363306 -160
rect 363374 -216 363430 -160
rect 363498 -216 363554 -160
rect 363622 -216 363678 -160
rect 363250 -340 363306 -284
rect 363374 -340 363430 -284
rect 363498 -340 363554 -284
rect 363622 -340 363678 -284
rect 363250 -464 363306 -408
rect 363374 -464 363430 -408
rect 363498 -464 363554 -408
rect 363622 -464 363678 -408
rect 363250 -588 363306 -532
rect 363374 -588 363430 -532
rect 363498 -588 363554 -532
rect 363622 -588 363678 -532
rect 366970 208294 367026 208350
rect 367094 208294 367150 208350
rect 367218 208294 367274 208350
rect 367342 208294 367398 208350
rect 366970 208170 367026 208226
rect 367094 208170 367150 208226
rect 367218 208170 367274 208226
rect 367342 208170 367398 208226
rect 366970 208046 367026 208102
rect 367094 208046 367150 208102
rect 367218 208046 367274 208102
rect 367342 208046 367398 208102
rect 366970 207922 367026 207978
rect 367094 207922 367150 207978
rect 367218 207922 367274 207978
rect 367342 207922 367398 207978
rect 373478 208294 373534 208350
rect 373602 208294 373658 208350
rect 373478 208170 373534 208226
rect 373602 208170 373658 208226
rect 373478 208046 373534 208102
rect 373602 208046 373658 208102
rect 373478 207922 373534 207978
rect 373602 207922 373658 207978
rect 366970 190294 367026 190350
rect 367094 190294 367150 190350
rect 367218 190294 367274 190350
rect 367342 190294 367398 190350
rect 366970 190170 367026 190226
rect 367094 190170 367150 190226
rect 367218 190170 367274 190226
rect 367342 190170 367398 190226
rect 366970 190046 367026 190102
rect 367094 190046 367150 190102
rect 367218 190046 367274 190102
rect 367342 190046 367398 190102
rect 366970 189922 367026 189978
rect 367094 189922 367150 189978
rect 367218 189922 367274 189978
rect 367342 189922 367398 189978
rect 366970 172294 367026 172350
rect 367094 172294 367150 172350
rect 367218 172294 367274 172350
rect 367342 172294 367398 172350
rect 366970 172170 367026 172226
rect 367094 172170 367150 172226
rect 367218 172170 367274 172226
rect 367342 172170 367398 172226
rect 366970 172046 367026 172102
rect 367094 172046 367150 172102
rect 367218 172046 367274 172102
rect 367342 172046 367398 172102
rect 366970 171922 367026 171978
rect 367094 171922 367150 171978
rect 367218 171922 367274 171978
rect 367342 171922 367398 171978
rect 366970 154294 367026 154350
rect 367094 154294 367150 154350
rect 367218 154294 367274 154350
rect 367342 154294 367398 154350
rect 366970 154170 367026 154226
rect 367094 154170 367150 154226
rect 367218 154170 367274 154226
rect 367342 154170 367398 154226
rect 366970 154046 367026 154102
rect 367094 154046 367150 154102
rect 367218 154046 367274 154102
rect 367342 154046 367398 154102
rect 366970 153922 367026 153978
rect 367094 153922 367150 153978
rect 367218 153922 367274 153978
rect 367342 153922 367398 153978
rect 366970 136294 367026 136350
rect 367094 136294 367150 136350
rect 367218 136294 367274 136350
rect 367342 136294 367398 136350
rect 366970 136170 367026 136226
rect 367094 136170 367150 136226
rect 367218 136170 367274 136226
rect 367342 136170 367398 136226
rect 366970 136046 367026 136102
rect 367094 136046 367150 136102
rect 367218 136046 367274 136102
rect 367342 136046 367398 136102
rect 366970 135922 367026 135978
rect 367094 135922 367150 135978
rect 367218 135922 367274 135978
rect 367342 135922 367398 135978
rect 366970 118294 367026 118350
rect 367094 118294 367150 118350
rect 367218 118294 367274 118350
rect 367342 118294 367398 118350
rect 366970 118170 367026 118226
rect 367094 118170 367150 118226
rect 367218 118170 367274 118226
rect 367342 118170 367398 118226
rect 366970 118046 367026 118102
rect 367094 118046 367150 118102
rect 367218 118046 367274 118102
rect 367342 118046 367398 118102
rect 366970 117922 367026 117978
rect 367094 117922 367150 117978
rect 367218 117922 367274 117978
rect 367342 117922 367398 117978
rect 366970 100294 367026 100350
rect 367094 100294 367150 100350
rect 367218 100294 367274 100350
rect 367342 100294 367398 100350
rect 366970 100170 367026 100226
rect 367094 100170 367150 100226
rect 367218 100170 367274 100226
rect 367342 100170 367398 100226
rect 366970 100046 367026 100102
rect 367094 100046 367150 100102
rect 367218 100046 367274 100102
rect 367342 100046 367398 100102
rect 366970 99922 367026 99978
rect 367094 99922 367150 99978
rect 367218 99922 367274 99978
rect 367342 99922 367398 99978
rect 366970 82294 367026 82350
rect 367094 82294 367150 82350
rect 367218 82294 367274 82350
rect 367342 82294 367398 82350
rect 366970 82170 367026 82226
rect 367094 82170 367150 82226
rect 367218 82170 367274 82226
rect 367342 82170 367398 82226
rect 366970 82046 367026 82102
rect 367094 82046 367150 82102
rect 367218 82046 367274 82102
rect 367342 82046 367398 82102
rect 366970 81922 367026 81978
rect 367094 81922 367150 81978
rect 367218 81922 367274 81978
rect 367342 81922 367398 81978
rect 366970 64294 367026 64350
rect 367094 64294 367150 64350
rect 367218 64294 367274 64350
rect 367342 64294 367398 64350
rect 366970 64170 367026 64226
rect 367094 64170 367150 64226
rect 367218 64170 367274 64226
rect 367342 64170 367398 64226
rect 366970 64046 367026 64102
rect 367094 64046 367150 64102
rect 367218 64046 367274 64102
rect 367342 64046 367398 64102
rect 366970 63922 367026 63978
rect 367094 63922 367150 63978
rect 367218 63922 367274 63978
rect 367342 63922 367398 63978
rect 366970 46294 367026 46350
rect 367094 46294 367150 46350
rect 367218 46294 367274 46350
rect 367342 46294 367398 46350
rect 366970 46170 367026 46226
rect 367094 46170 367150 46226
rect 367218 46170 367274 46226
rect 367342 46170 367398 46226
rect 366970 46046 367026 46102
rect 367094 46046 367150 46102
rect 367218 46046 367274 46102
rect 367342 46046 367398 46102
rect 366970 45922 367026 45978
rect 367094 45922 367150 45978
rect 367218 45922 367274 45978
rect 367342 45922 367398 45978
rect 366970 28294 367026 28350
rect 367094 28294 367150 28350
rect 367218 28294 367274 28350
rect 367342 28294 367398 28350
rect 366970 28170 367026 28226
rect 367094 28170 367150 28226
rect 367218 28170 367274 28226
rect 367342 28170 367398 28226
rect 366970 28046 367026 28102
rect 367094 28046 367150 28102
rect 367218 28046 367274 28102
rect 367342 28046 367398 28102
rect 366970 27922 367026 27978
rect 367094 27922 367150 27978
rect 367218 27922 367274 27978
rect 367342 27922 367398 27978
rect 366970 10294 367026 10350
rect 367094 10294 367150 10350
rect 367218 10294 367274 10350
rect 367342 10294 367398 10350
rect 366970 10170 367026 10226
rect 367094 10170 367150 10226
rect 367218 10170 367274 10226
rect 367342 10170 367398 10226
rect 366970 10046 367026 10102
rect 367094 10046 367150 10102
rect 367218 10046 367274 10102
rect 367342 10046 367398 10102
rect 366970 9922 367026 9978
rect 367094 9922 367150 9978
rect 367218 9922 367274 9978
rect 367342 9922 367398 9978
rect 366970 -1176 367026 -1120
rect 367094 -1176 367150 -1120
rect 367218 -1176 367274 -1120
rect 367342 -1176 367398 -1120
rect 366970 -1300 367026 -1244
rect 367094 -1300 367150 -1244
rect 367218 -1300 367274 -1244
rect 367342 -1300 367398 -1244
rect 366970 -1424 367026 -1368
rect 367094 -1424 367150 -1368
rect 367218 -1424 367274 -1368
rect 367342 -1424 367398 -1368
rect 366970 -1548 367026 -1492
rect 367094 -1548 367150 -1492
rect 367218 -1548 367274 -1492
rect 367342 -1548 367398 -1492
rect 381250 202294 381306 202350
rect 381374 202294 381430 202350
rect 381498 202294 381554 202350
rect 381622 202294 381678 202350
rect 381250 202170 381306 202226
rect 381374 202170 381430 202226
rect 381498 202170 381554 202226
rect 381622 202170 381678 202226
rect 381250 202046 381306 202102
rect 381374 202046 381430 202102
rect 381498 202046 381554 202102
rect 381622 202046 381678 202102
rect 381250 201922 381306 201978
rect 381374 201922 381430 201978
rect 381498 201922 381554 201978
rect 381622 201922 381678 201978
rect 381250 184294 381306 184350
rect 381374 184294 381430 184350
rect 381498 184294 381554 184350
rect 381622 184294 381678 184350
rect 381250 184170 381306 184226
rect 381374 184170 381430 184226
rect 381498 184170 381554 184226
rect 381622 184170 381678 184226
rect 381250 184046 381306 184102
rect 381374 184046 381430 184102
rect 381498 184046 381554 184102
rect 381622 184046 381678 184102
rect 381250 183922 381306 183978
rect 381374 183922 381430 183978
rect 381498 183922 381554 183978
rect 381622 183922 381678 183978
rect 381250 166294 381306 166350
rect 381374 166294 381430 166350
rect 381498 166294 381554 166350
rect 381622 166294 381678 166350
rect 381250 166170 381306 166226
rect 381374 166170 381430 166226
rect 381498 166170 381554 166226
rect 381622 166170 381678 166226
rect 381250 166046 381306 166102
rect 381374 166046 381430 166102
rect 381498 166046 381554 166102
rect 381622 166046 381678 166102
rect 381250 165922 381306 165978
rect 381374 165922 381430 165978
rect 381498 165922 381554 165978
rect 381622 165922 381678 165978
rect 381250 148294 381306 148350
rect 381374 148294 381430 148350
rect 381498 148294 381554 148350
rect 381622 148294 381678 148350
rect 381250 148170 381306 148226
rect 381374 148170 381430 148226
rect 381498 148170 381554 148226
rect 381622 148170 381678 148226
rect 381250 148046 381306 148102
rect 381374 148046 381430 148102
rect 381498 148046 381554 148102
rect 381622 148046 381678 148102
rect 381250 147922 381306 147978
rect 381374 147922 381430 147978
rect 381498 147922 381554 147978
rect 381622 147922 381678 147978
rect 381250 130294 381306 130350
rect 381374 130294 381430 130350
rect 381498 130294 381554 130350
rect 381622 130294 381678 130350
rect 381250 130170 381306 130226
rect 381374 130170 381430 130226
rect 381498 130170 381554 130226
rect 381622 130170 381678 130226
rect 381250 130046 381306 130102
rect 381374 130046 381430 130102
rect 381498 130046 381554 130102
rect 381622 130046 381678 130102
rect 381250 129922 381306 129978
rect 381374 129922 381430 129978
rect 381498 129922 381554 129978
rect 381622 129922 381678 129978
rect 381250 112294 381306 112350
rect 381374 112294 381430 112350
rect 381498 112294 381554 112350
rect 381622 112294 381678 112350
rect 381250 112170 381306 112226
rect 381374 112170 381430 112226
rect 381498 112170 381554 112226
rect 381622 112170 381678 112226
rect 381250 112046 381306 112102
rect 381374 112046 381430 112102
rect 381498 112046 381554 112102
rect 381622 112046 381678 112102
rect 381250 111922 381306 111978
rect 381374 111922 381430 111978
rect 381498 111922 381554 111978
rect 381622 111922 381678 111978
rect 381250 94294 381306 94350
rect 381374 94294 381430 94350
rect 381498 94294 381554 94350
rect 381622 94294 381678 94350
rect 381250 94170 381306 94226
rect 381374 94170 381430 94226
rect 381498 94170 381554 94226
rect 381622 94170 381678 94226
rect 381250 94046 381306 94102
rect 381374 94046 381430 94102
rect 381498 94046 381554 94102
rect 381622 94046 381678 94102
rect 381250 93922 381306 93978
rect 381374 93922 381430 93978
rect 381498 93922 381554 93978
rect 381622 93922 381678 93978
rect 381250 76294 381306 76350
rect 381374 76294 381430 76350
rect 381498 76294 381554 76350
rect 381622 76294 381678 76350
rect 381250 76170 381306 76226
rect 381374 76170 381430 76226
rect 381498 76170 381554 76226
rect 381622 76170 381678 76226
rect 381250 76046 381306 76102
rect 381374 76046 381430 76102
rect 381498 76046 381554 76102
rect 381622 76046 381678 76102
rect 381250 75922 381306 75978
rect 381374 75922 381430 75978
rect 381498 75922 381554 75978
rect 381622 75922 381678 75978
rect 381250 58294 381306 58350
rect 381374 58294 381430 58350
rect 381498 58294 381554 58350
rect 381622 58294 381678 58350
rect 381250 58170 381306 58226
rect 381374 58170 381430 58226
rect 381498 58170 381554 58226
rect 381622 58170 381678 58226
rect 381250 58046 381306 58102
rect 381374 58046 381430 58102
rect 381498 58046 381554 58102
rect 381622 58046 381678 58102
rect 381250 57922 381306 57978
rect 381374 57922 381430 57978
rect 381498 57922 381554 57978
rect 381622 57922 381678 57978
rect 381250 40294 381306 40350
rect 381374 40294 381430 40350
rect 381498 40294 381554 40350
rect 381622 40294 381678 40350
rect 381250 40170 381306 40226
rect 381374 40170 381430 40226
rect 381498 40170 381554 40226
rect 381622 40170 381678 40226
rect 381250 40046 381306 40102
rect 381374 40046 381430 40102
rect 381498 40046 381554 40102
rect 381622 40046 381678 40102
rect 381250 39922 381306 39978
rect 381374 39922 381430 39978
rect 381498 39922 381554 39978
rect 381622 39922 381678 39978
rect 381250 22294 381306 22350
rect 381374 22294 381430 22350
rect 381498 22294 381554 22350
rect 381622 22294 381678 22350
rect 381250 22170 381306 22226
rect 381374 22170 381430 22226
rect 381498 22170 381554 22226
rect 381622 22170 381678 22226
rect 381250 22046 381306 22102
rect 381374 22046 381430 22102
rect 381498 22046 381554 22102
rect 381622 22046 381678 22102
rect 381250 21922 381306 21978
rect 381374 21922 381430 21978
rect 381498 21922 381554 21978
rect 381622 21922 381678 21978
rect 381250 4294 381306 4350
rect 381374 4294 381430 4350
rect 381498 4294 381554 4350
rect 381622 4294 381678 4350
rect 381250 4170 381306 4226
rect 381374 4170 381430 4226
rect 381498 4170 381554 4226
rect 381622 4170 381678 4226
rect 381250 4046 381306 4102
rect 381374 4046 381430 4102
rect 381498 4046 381554 4102
rect 381622 4046 381678 4102
rect 381250 3922 381306 3978
rect 381374 3922 381430 3978
rect 381498 3922 381554 3978
rect 381622 3922 381678 3978
rect 381250 -216 381306 -160
rect 381374 -216 381430 -160
rect 381498 -216 381554 -160
rect 381622 -216 381678 -160
rect 381250 -340 381306 -284
rect 381374 -340 381430 -284
rect 381498 -340 381554 -284
rect 381622 -340 381678 -284
rect 381250 -464 381306 -408
rect 381374 -464 381430 -408
rect 381498 -464 381554 -408
rect 381622 -464 381678 -408
rect 381250 -588 381306 -532
rect 381374 -588 381430 -532
rect 381498 -588 381554 -532
rect 381622 -588 381678 -532
rect 384970 208294 385026 208350
rect 385094 208294 385150 208350
rect 385218 208294 385274 208350
rect 385342 208294 385398 208350
rect 384970 208170 385026 208226
rect 385094 208170 385150 208226
rect 385218 208170 385274 208226
rect 385342 208170 385398 208226
rect 384970 208046 385026 208102
rect 385094 208046 385150 208102
rect 385218 208046 385274 208102
rect 385342 208046 385398 208102
rect 384970 207922 385026 207978
rect 385094 207922 385150 207978
rect 385218 207922 385274 207978
rect 385342 207922 385398 207978
rect 384970 190294 385026 190350
rect 385094 190294 385150 190350
rect 385218 190294 385274 190350
rect 385342 190294 385398 190350
rect 384970 190170 385026 190226
rect 385094 190170 385150 190226
rect 385218 190170 385274 190226
rect 385342 190170 385398 190226
rect 384970 190046 385026 190102
rect 385094 190046 385150 190102
rect 385218 190046 385274 190102
rect 385342 190046 385398 190102
rect 384970 189922 385026 189978
rect 385094 189922 385150 189978
rect 385218 189922 385274 189978
rect 385342 189922 385398 189978
rect 384970 172294 385026 172350
rect 385094 172294 385150 172350
rect 385218 172294 385274 172350
rect 385342 172294 385398 172350
rect 384970 172170 385026 172226
rect 385094 172170 385150 172226
rect 385218 172170 385274 172226
rect 385342 172170 385398 172226
rect 384970 172046 385026 172102
rect 385094 172046 385150 172102
rect 385218 172046 385274 172102
rect 385342 172046 385398 172102
rect 384970 171922 385026 171978
rect 385094 171922 385150 171978
rect 385218 171922 385274 171978
rect 385342 171922 385398 171978
rect 384970 154294 385026 154350
rect 385094 154294 385150 154350
rect 385218 154294 385274 154350
rect 385342 154294 385398 154350
rect 384970 154170 385026 154226
rect 385094 154170 385150 154226
rect 385218 154170 385274 154226
rect 385342 154170 385398 154226
rect 384970 154046 385026 154102
rect 385094 154046 385150 154102
rect 385218 154046 385274 154102
rect 385342 154046 385398 154102
rect 384970 153922 385026 153978
rect 385094 153922 385150 153978
rect 385218 153922 385274 153978
rect 385342 153922 385398 153978
rect 384970 136294 385026 136350
rect 385094 136294 385150 136350
rect 385218 136294 385274 136350
rect 385342 136294 385398 136350
rect 384970 136170 385026 136226
rect 385094 136170 385150 136226
rect 385218 136170 385274 136226
rect 385342 136170 385398 136226
rect 384970 136046 385026 136102
rect 385094 136046 385150 136102
rect 385218 136046 385274 136102
rect 385342 136046 385398 136102
rect 384970 135922 385026 135978
rect 385094 135922 385150 135978
rect 385218 135922 385274 135978
rect 385342 135922 385398 135978
rect 384970 118294 385026 118350
rect 385094 118294 385150 118350
rect 385218 118294 385274 118350
rect 385342 118294 385398 118350
rect 384970 118170 385026 118226
rect 385094 118170 385150 118226
rect 385218 118170 385274 118226
rect 385342 118170 385398 118226
rect 384970 118046 385026 118102
rect 385094 118046 385150 118102
rect 385218 118046 385274 118102
rect 385342 118046 385398 118102
rect 384970 117922 385026 117978
rect 385094 117922 385150 117978
rect 385218 117922 385274 117978
rect 385342 117922 385398 117978
rect 384970 100294 385026 100350
rect 385094 100294 385150 100350
rect 385218 100294 385274 100350
rect 385342 100294 385398 100350
rect 384970 100170 385026 100226
rect 385094 100170 385150 100226
rect 385218 100170 385274 100226
rect 385342 100170 385398 100226
rect 384970 100046 385026 100102
rect 385094 100046 385150 100102
rect 385218 100046 385274 100102
rect 385342 100046 385398 100102
rect 384970 99922 385026 99978
rect 385094 99922 385150 99978
rect 385218 99922 385274 99978
rect 385342 99922 385398 99978
rect 384970 82294 385026 82350
rect 385094 82294 385150 82350
rect 385218 82294 385274 82350
rect 385342 82294 385398 82350
rect 384970 82170 385026 82226
rect 385094 82170 385150 82226
rect 385218 82170 385274 82226
rect 385342 82170 385398 82226
rect 384970 82046 385026 82102
rect 385094 82046 385150 82102
rect 385218 82046 385274 82102
rect 385342 82046 385398 82102
rect 384970 81922 385026 81978
rect 385094 81922 385150 81978
rect 385218 81922 385274 81978
rect 385342 81922 385398 81978
rect 384970 64294 385026 64350
rect 385094 64294 385150 64350
rect 385218 64294 385274 64350
rect 385342 64294 385398 64350
rect 384970 64170 385026 64226
rect 385094 64170 385150 64226
rect 385218 64170 385274 64226
rect 385342 64170 385398 64226
rect 384970 64046 385026 64102
rect 385094 64046 385150 64102
rect 385218 64046 385274 64102
rect 385342 64046 385398 64102
rect 384970 63922 385026 63978
rect 385094 63922 385150 63978
rect 385218 63922 385274 63978
rect 385342 63922 385398 63978
rect 384970 46294 385026 46350
rect 385094 46294 385150 46350
rect 385218 46294 385274 46350
rect 385342 46294 385398 46350
rect 384970 46170 385026 46226
rect 385094 46170 385150 46226
rect 385218 46170 385274 46226
rect 385342 46170 385398 46226
rect 384970 46046 385026 46102
rect 385094 46046 385150 46102
rect 385218 46046 385274 46102
rect 385342 46046 385398 46102
rect 384970 45922 385026 45978
rect 385094 45922 385150 45978
rect 385218 45922 385274 45978
rect 385342 45922 385398 45978
rect 384970 28294 385026 28350
rect 385094 28294 385150 28350
rect 385218 28294 385274 28350
rect 385342 28294 385398 28350
rect 384970 28170 385026 28226
rect 385094 28170 385150 28226
rect 385218 28170 385274 28226
rect 385342 28170 385398 28226
rect 384970 28046 385026 28102
rect 385094 28046 385150 28102
rect 385218 28046 385274 28102
rect 385342 28046 385398 28102
rect 384970 27922 385026 27978
rect 385094 27922 385150 27978
rect 385218 27922 385274 27978
rect 385342 27922 385398 27978
rect 384970 10294 385026 10350
rect 385094 10294 385150 10350
rect 385218 10294 385274 10350
rect 385342 10294 385398 10350
rect 384970 10170 385026 10226
rect 385094 10170 385150 10226
rect 385218 10170 385274 10226
rect 385342 10170 385398 10226
rect 384970 10046 385026 10102
rect 385094 10046 385150 10102
rect 385218 10046 385274 10102
rect 385342 10046 385398 10102
rect 384970 9922 385026 9978
rect 385094 9922 385150 9978
rect 385218 9922 385274 9978
rect 385342 9922 385398 9978
rect 384970 -1176 385026 -1120
rect 385094 -1176 385150 -1120
rect 385218 -1176 385274 -1120
rect 385342 -1176 385398 -1120
rect 384970 -1300 385026 -1244
rect 385094 -1300 385150 -1244
rect 385218 -1300 385274 -1244
rect 385342 -1300 385398 -1244
rect 384970 -1424 385026 -1368
rect 385094 -1424 385150 -1368
rect 385218 -1424 385274 -1368
rect 385342 -1424 385398 -1368
rect 384970 -1548 385026 -1492
rect 385094 -1548 385150 -1492
rect 385218 -1548 385274 -1492
rect 385342 -1548 385398 -1492
rect 399250 202294 399306 202350
rect 399374 202294 399430 202350
rect 399498 202294 399554 202350
rect 399622 202294 399678 202350
rect 399250 202170 399306 202226
rect 399374 202170 399430 202226
rect 399498 202170 399554 202226
rect 399622 202170 399678 202226
rect 399250 202046 399306 202102
rect 399374 202046 399430 202102
rect 399498 202046 399554 202102
rect 399622 202046 399678 202102
rect 399250 201922 399306 201978
rect 399374 201922 399430 201978
rect 399498 201922 399554 201978
rect 399622 201922 399678 201978
rect 399250 184294 399306 184350
rect 399374 184294 399430 184350
rect 399498 184294 399554 184350
rect 399622 184294 399678 184350
rect 399250 184170 399306 184226
rect 399374 184170 399430 184226
rect 399498 184170 399554 184226
rect 399622 184170 399678 184226
rect 399250 184046 399306 184102
rect 399374 184046 399430 184102
rect 399498 184046 399554 184102
rect 399622 184046 399678 184102
rect 399250 183922 399306 183978
rect 399374 183922 399430 183978
rect 399498 183922 399554 183978
rect 399622 183922 399678 183978
rect 399250 166294 399306 166350
rect 399374 166294 399430 166350
rect 399498 166294 399554 166350
rect 399622 166294 399678 166350
rect 399250 166170 399306 166226
rect 399374 166170 399430 166226
rect 399498 166170 399554 166226
rect 399622 166170 399678 166226
rect 399250 166046 399306 166102
rect 399374 166046 399430 166102
rect 399498 166046 399554 166102
rect 399622 166046 399678 166102
rect 399250 165922 399306 165978
rect 399374 165922 399430 165978
rect 399498 165922 399554 165978
rect 399622 165922 399678 165978
rect 399250 148294 399306 148350
rect 399374 148294 399430 148350
rect 399498 148294 399554 148350
rect 399622 148294 399678 148350
rect 399250 148170 399306 148226
rect 399374 148170 399430 148226
rect 399498 148170 399554 148226
rect 399622 148170 399678 148226
rect 399250 148046 399306 148102
rect 399374 148046 399430 148102
rect 399498 148046 399554 148102
rect 399622 148046 399678 148102
rect 399250 147922 399306 147978
rect 399374 147922 399430 147978
rect 399498 147922 399554 147978
rect 399622 147922 399678 147978
rect 399250 130294 399306 130350
rect 399374 130294 399430 130350
rect 399498 130294 399554 130350
rect 399622 130294 399678 130350
rect 399250 130170 399306 130226
rect 399374 130170 399430 130226
rect 399498 130170 399554 130226
rect 399622 130170 399678 130226
rect 399250 130046 399306 130102
rect 399374 130046 399430 130102
rect 399498 130046 399554 130102
rect 399622 130046 399678 130102
rect 399250 129922 399306 129978
rect 399374 129922 399430 129978
rect 399498 129922 399554 129978
rect 399622 129922 399678 129978
rect 399250 112294 399306 112350
rect 399374 112294 399430 112350
rect 399498 112294 399554 112350
rect 399622 112294 399678 112350
rect 399250 112170 399306 112226
rect 399374 112170 399430 112226
rect 399498 112170 399554 112226
rect 399622 112170 399678 112226
rect 399250 112046 399306 112102
rect 399374 112046 399430 112102
rect 399498 112046 399554 112102
rect 399622 112046 399678 112102
rect 399250 111922 399306 111978
rect 399374 111922 399430 111978
rect 399498 111922 399554 111978
rect 399622 111922 399678 111978
rect 399250 94294 399306 94350
rect 399374 94294 399430 94350
rect 399498 94294 399554 94350
rect 399622 94294 399678 94350
rect 399250 94170 399306 94226
rect 399374 94170 399430 94226
rect 399498 94170 399554 94226
rect 399622 94170 399678 94226
rect 399250 94046 399306 94102
rect 399374 94046 399430 94102
rect 399498 94046 399554 94102
rect 399622 94046 399678 94102
rect 399250 93922 399306 93978
rect 399374 93922 399430 93978
rect 399498 93922 399554 93978
rect 399622 93922 399678 93978
rect 399250 76294 399306 76350
rect 399374 76294 399430 76350
rect 399498 76294 399554 76350
rect 399622 76294 399678 76350
rect 399250 76170 399306 76226
rect 399374 76170 399430 76226
rect 399498 76170 399554 76226
rect 399622 76170 399678 76226
rect 399250 76046 399306 76102
rect 399374 76046 399430 76102
rect 399498 76046 399554 76102
rect 399622 76046 399678 76102
rect 399250 75922 399306 75978
rect 399374 75922 399430 75978
rect 399498 75922 399554 75978
rect 399622 75922 399678 75978
rect 399250 58294 399306 58350
rect 399374 58294 399430 58350
rect 399498 58294 399554 58350
rect 399622 58294 399678 58350
rect 399250 58170 399306 58226
rect 399374 58170 399430 58226
rect 399498 58170 399554 58226
rect 399622 58170 399678 58226
rect 399250 58046 399306 58102
rect 399374 58046 399430 58102
rect 399498 58046 399554 58102
rect 399622 58046 399678 58102
rect 399250 57922 399306 57978
rect 399374 57922 399430 57978
rect 399498 57922 399554 57978
rect 399622 57922 399678 57978
rect 399250 40294 399306 40350
rect 399374 40294 399430 40350
rect 399498 40294 399554 40350
rect 399622 40294 399678 40350
rect 399250 40170 399306 40226
rect 399374 40170 399430 40226
rect 399498 40170 399554 40226
rect 399622 40170 399678 40226
rect 399250 40046 399306 40102
rect 399374 40046 399430 40102
rect 399498 40046 399554 40102
rect 399622 40046 399678 40102
rect 399250 39922 399306 39978
rect 399374 39922 399430 39978
rect 399498 39922 399554 39978
rect 399622 39922 399678 39978
rect 399250 22294 399306 22350
rect 399374 22294 399430 22350
rect 399498 22294 399554 22350
rect 399622 22294 399678 22350
rect 399250 22170 399306 22226
rect 399374 22170 399430 22226
rect 399498 22170 399554 22226
rect 399622 22170 399678 22226
rect 399250 22046 399306 22102
rect 399374 22046 399430 22102
rect 399498 22046 399554 22102
rect 399622 22046 399678 22102
rect 399250 21922 399306 21978
rect 399374 21922 399430 21978
rect 399498 21922 399554 21978
rect 399622 21922 399678 21978
rect 399250 4294 399306 4350
rect 399374 4294 399430 4350
rect 399498 4294 399554 4350
rect 399622 4294 399678 4350
rect 399250 4170 399306 4226
rect 399374 4170 399430 4226
rect 399498 4170 399554 4226
rect 399622 4170 399678 4226
rect 399250 4046 399306 4102
rect 399374 4046 399430 4102
rect 399498 4046 399554 4102
rect 399622 4046 399678 4102
rect 399250 3922 399306 3978
rect 399374 3922 399430 3978
rect 399498 3922 399554 3978
rect 399622 3922 399678 3978
rect 399250 -216 399306 -160
rect 399374 -216 399430 -160
rect 399498 -216 399554 -160
rect 399622 -216 399678 -160
rect 399250 -340 399306 -284
rect 399374 -340 399430 -284
rect 399498 -340 399554 -284
rect 399622 -340 399678 -284
rect 399250 -464 399306 -408
rect 399374 -464 399430 -408
rect 399498 -464 399554 -408
rect 399622 -464 399678 -408
rect 399250 -588 399306 -532
rect 399374 -588 399430 -532
rect 399498 -588 399554 -532
rect 399622 -588 399678 -532
rect 402970 208294 403026 208350
rect 403094 208294 403150 208350
rect 403218 208294 403274 208350
rect 403342 208294 403398 208350
rect 402970 208170 403026 208226
rect 403094 208170 403150 208226
rect 403218 208170 403274 208226
rect 403342 208170 403398 208226
rect 402970 208046 403026 208102
rect 403094 208046 403150 208102
rect 403218 208046 403274 208102
rect 403342 208046 403398 208102
rect 402970 207922 403026 207978
rect 403094 207922 403150 207978
rect 403218 207922 403274 207978
rect 403342 207922 403398 207978
rect 404198 208294 404254 208350
rect 404322 208294 404378 208350
rect 404198 208170 404254 208226
rect 404322 208170 404378 208226
rect 404198 208046 404254 208102
rect 404322 208046 404378 208102
rect 404198 207922 404254 207978
rect 404322 207922 404378 207978
rect 402970 190294 403026 190350
rect 403094 190294 403150 190350
rect 403218 190294 403274 190350
rect 403342 190294 403398 190350
rect 402970 190170 403026 190226
rect 403094 190170 403150 190226
rect 403218 190170 403274 190226
rect 403342 190170 403398 190226
rect 402970 190046 403026 190102
rect 403094 190046 403150 190102
rect 403218 190046 403274 190102
rect 403342 190046 403398 190102
rect 402970 189922 403026 189978
rect 403094 189922 403150 189978
rect 403218 189922 403274 189978
rect 403342 189922 403398 189978
rect 402970 172294 403026 172350
rect 403094 172294 403150 172350
rect 403218 172294 403274 172350
rect 403342 172294 403398 172350
rect 402970 172170 403026 172226
rect 403094 172170 403150 172226
rect 403218 172170 403274 172226
rect 403342 172170 403398 172226
rect 402970 172046 403026 172102
rect 403094 172046 403150 172102
rect 403218 172046 403274 172102
rect 403342 172046 403398 172102
rect 402970 171922 403026 171978
rect 403094 171922 403150 171978
rect 403218 171922 403274 171978
rect 403342 171922 403398 171978
rect 402970 154294 403026 154350
rect 403094 154294 403150 154350
rect 403218 154294 403274 154350
rect 403342 154294 403398 154350
rect 402970 154170 403026 154226
rect 403094 154170 403150 154226
rect 403218 154170 403274 154226
rect 403342 154170 403398 154226
rect 402970 154046 403026 154102
rect 403094 154046 403150 154102
rect 403218 154046 403274 154102
rect 403342 154046 403398 154102
rect 402970 153922 403026 153978
rect 403094 153922 403150 153978
rect 403218 153922 403274 153978
rect 403342 153922 403398 153978
rect 402970 136294 403026 136350
rect 403094 136294 403150 136350
rect 403218 136294 403274 136350
rect 403342 136294 403398 136350
rect 402970 136170 403026 136226
rect 403094 136170 403150 136226
rect 403218 136170 403274 136226
rect 403342 136170 403398 136226
rect 402970 136046 403026 136102
rect 403094 136046 403150 136102
rect 403218 136046 403274 136102
rect 403342 136046 403398 136102
rect 402970 135922 403026 135978
rect 403094 135922 403150 135978
rect 403218 135922 403274 135978
rect 403342 135922 403398 135978
rect 402970 118294 403026 118350
rect 403094 118294 403150 118350
rect 403218 118294 403274 118350
rect 403342 118294 403398 118350
rect 402970 118170 403026 118226
rect 403094 118170 403150 118226
rect 403218 118170 403274 118226
rect 403342 118170 403398 118226
rect 402970 118046 403026 118102
rect 403094 118046 403150 118102
rect 403218 118046 403274 118102
rect 403342 118046 403398 118102
rect 402970 117922 403026 117978
rect 403094 117922 403150 117978
rect 403218 117922 403274 117978
rect 403342 117922 403398 117978
rect 402970 100294 403026 100350
rect 403094 100294 403150 100350
rect 403218 100294 403274 100350
rect 403342 100294 403398 100350
rect 402970 100170 403026 100226
rect 403094 100170 403150 100226
rect 403218 100170 403274 100226
rect 403342 100170 403398 100226
rect 402970 100046 403026 100102
rect 403094 100046 403150 100102
rect 403218 100046 403274 100102
rect 403342 100046 403398 100102
rect 402970 99922 403026 99978
rect 403094 99922 403150 99978
rect 403218 99922 403274 99978
rect 403342 99922 403398 99978
rect 402970 82294 403026 82350
rect 403094 82294 403150 82350
rect 403218 82294 403274 82350
rect 403342 82294 403398 82350
rect 402970 82170 403026 82226
rect 403094 82170 403150 82226
rect 403218 82170 403274 82226
rect 403342 82170 403398 82226
rect 402970 82046 403026 82102
rect 403094 82046 403150 82102
rect 403218 82046 403274 82102
rect 403342 82046 403398 82102
rect 402970 81922 403026 81978
rect 403094 81922 403150 81978
rect 403218 81922 403274 81978
rect 403342 81922 403398 81978
rect 402970 64294 403026 64350
rect 403094 64294 403150 64350
rect 403218 64294 403274 64350
rect 403342 64294 403398 64350
rect 402970 64170 403026 64226
rect 403094 64170 403150 64226
rect 403218 64170 403274 64226
rect 403342 64170 403398 64226
rect 402970 64046 403026 64102
rect 403094 64046 403150 64102
rect 403218 64046 403274 64102
rect 403342 64046 403398 64102
rect 402970 63922 403026 63978
rect 403094 63922 403150 63978
rect 403218 63922 403274 63978
rect 403342 63922 403398 63978
rect 402970 46294 403026 46350
rect 403094 46294 403150 46350
rect 403218 46294 403274 46350
rect 403342 46294 403398 46350
rect 402970 46170 403026 46226
rect 403094 46170 403150 46226
rect 403218 46170 403274 46226
rect 403342 46170 403398 46226
rect 402970 46046 403026 46102
rect 403094 46046 403150 46102
rect 403218 46046 403274 46102
rect 403342 46046 403398 46102
rect 402970 45922 403026 45978
rect 403094 45922 403150 45978
rect 403218 45922 403274 45978
rect 403342 45922 403398 45978
rect 402970 28294 403026 28350
rect 403094 28294 403150 28350
rect 403218 28294 403274 28350
rect 403342 28294 403398 28350
rect 402970 28170 403026 28226
rect 403094 28170 403150 28226
rect 403218 28170 403274 28226
rect 403342 28170 403398 28226
rect 402970 28046 403026 28102
rect 403094 28046 403150 28102
rect 403218 28046 403274 28102
rect 403342 28046 403398 28102
rect 402970 27922 403026 27978
rect 403094 27922 403150 27978
rect 403218 27922 403274 27978
rect 403342 27922 403398 27978
rect 402970 10294 403026 10350
rect 403094 10294 403150 10350
rect 403218 10294 403274 10350
rect 403342 10294 403398 10350
rect 402970 10170 403026 10226
rect 403094 10170 403150 10226
rect 403218 10170 403274 10226
rect 403342 10170 403398 10226
rect 402970 10046 403026 10102
rect 403094 10046 403150 10102
rect 403218 10046 403274 10102
rect 403342 10046 403398 10102
rect 402970 9922 403026 9978
rect 403094 9922 403150 9978
rect 403218 9922 403274 9978
rect 403342 9922 403398 9978
rect 402970 -1176 403026 -1120
rect 403094 -1176 403150 -1120
rect 403218 -1176 403274 -1120
rect 403342 -1176 403398 -1120
rect 402970 -1300 403026 -1244
rect 403094 -1300 403150 -1244
rect 403218 -1300 403274 -1244
rect 403342 -1300 403398 -1244
rect 402970 -1424 403026 -1368
rect 403094 -1424 403150 -1368
rect 403218 -1424 403274 -1368
rect 403342 -1424 403398 -1368
rect 402970 -1548 403026 -1492
rect 403094 -1548 403150 -1492
rect 403218 -1548 403274 -1492
rect 403342 -1548 403398 -1492
rect 417250 202294 417306 202350
rect 417374 202294 417430 202350
rect 417498 202294 417554 202350
rect 417622 202294 417678 202350
rect 417250 202170 417306 202226
rect 417374 202170 417430 202226
rect 417498 202170 417554 202226
rect 417622 202170 417678 202226
rect 417250 202046 417306 202102
rect 417374 202046 417430 202102
rect 417498 202046 417554 202102
rect 417622 202046 417678 202102
rect 417250 201922 417306 201978
rect 417374 201922 417430 201978
rect 417498 201922 417554 201978
rect 417622 201922 417678 201978
rect 417250 184294 417306 184350
rect 417374 184294 417430 184350
rect 417498 184294 417554 184350
rect 417622 184294 417678 184350
rect 417250 184170 417306 184226
rect 417374 184170 417430 184226
rect 417498 184170 417554 184226
rect 417622 184170 417678 184226
rect 417250 184046 417306 184102
rect 417374 184046 417430 184102
rect 417498 184046 417554 184102
rect 417622 184046 417678 184102
rect 417250 183922 417306 183978
rect 417374 183922 417430 183978
rect 417498 183922 417554 183978
rect 417622 183922 417678 183978
rect 417250 166294 417306 166350
rect 417374 166294 417430 166350
rect 417498 166294 417554 166350
rect 417622 166294 417678 166350
rect 417250 166170 417306 166226
rect 417374 166170 417430 166226
rect 417498 166170 417554 166226
rect 417622 166170 417678 166226
rect 417250 166046 417306 166102
rect 417374 166046 417430 166102
rect 417498 166046 417554 166102
rect 417622 166046 417678 166102
rect 417250 165922 417306 165978
rect 417374 165922 417430 165978
rect 417498 165922 417554 165978
rect 417622 165922 417678 165978
rect 417250 148294 417306 148350
rect 417374 148294 417430 148350
rect 417498 148294 417554 148350
rect 417622 148294 417678 148350
rect 417250 148170 417306 148226
rect 417374 148170 417430 148226
rect 417498 148170 417554 148226
rect 417622 148170 417678 148226
rect 417250 148046 417306 148102
rect 417374 148046 417430 148102
rect 417498 148046 417554 148102
rect 417622 148046 417678 148102
rect 417250 147922 417306 147978
rect 417374 147922 417430 147978
rect 417498 147922 417554 147978
rect 417622 147922 417678 147978
rect 417250 130294 417306 130350
rect 417374 130294 417430 130350
rect 417498 130294 417554 130350
rect 417622 130294 417678 130350
rect 417250 130170 417306 130226
rect 417374 130170 417430 130226
rect 417498 130170 417554 130226
rect 417622 130170 417678 130226
rect 417250 130046 417306 130102
rect 417374 130046 417430 130102
rect 417498 130046 417554 130102
rect 417622 130046 417678 130102
rect 417250 129922 417306 129978
rect 417374 129922 417430 129978
rect 417498 129922 417554 129978
rect 417622 129922 417678 129978
rect 417250 112294 417306 112350
rect 417374 112294 417430 112350
rect 417498 112294 417554 112350
rect 417622 112294 417678 112350
rect 417250 112170 417306 112226
rect 417374 112170 417430 112226
rect 417498 112170 417554 112226
rect 417622 112170 417678 112226
rect 417250 112046 417306 112102
rect 417374 112046 417430 112102
rect 417498 112046 417554 112102
rect 417622 112046 417678 112102
rect 417250 111922 417306 111978
rect 417374 111922 417430 111978
rect 417498 111922 417554 111978
rect 417622 111922 417678 111978
rect 417250 94294 417306 94350
rect 417374 94294 417430 94350
rect 417498 94294 417554 94350
rect 417622 94294 417678 94350
rect 417250 94170 417306 94226
rect 417374 94170 417430 94226
rect 417498 94170 417554 94226
rect 417622 94170 417678 94226
rect 417250 94046 417306 94102
rect 417374 94046 417430 94102
rect 417498 94046 417554 94102
rect 417622 94046 417678 94102
rect 417250 93922 417306 93978
rect 417374 93922 417430 93978
rect 417498 93922 417554 93978
rect 417622 93922 417678 93978
rect 417250 76294 417306 76350
rect 417374 76294 417430 76350
rect 417498 76294 417554 76350
rect 417622 76294 417678 76350
rect 417250 76170 417306 76226
rect 417374 76170 417430 76226
rect 417498 76170 417554 76226
rect 417622 76170 417678 76226
rect 417250 76046 417306 76102
rect 417374 76046 417430 76102
rect 417498 76046 417554 76102
rect 417622 76046 417678 76102
rect 417250 75922 417306 75978
rect 417374 75922 417430 75978
rect 417498 75922 417554 75978
rect 417622 75922 417678 75978
rect 417250 58294 417306 58350
rect 417374 58294 417430 58350
rect 417498 58294 417554 58350
rect 417622 58294 417678 58350
rect 417250 58170 417306 58226
rect 417374 58170 417430 58226
rect 417498 58170 417554 58226
rect 417622 58170 417678 58226
rect 417250 58046 417306 58102
rect 417374 58046 417430 58102
rect 417498 58046 417554 58102
rect 417622 58046 417678 58102
rect 417250 57922 417306 57978
rect 417374 57922 417430 57978
rect 417498 57922 417554 57978
rect 417622 57922 417678 57978
rect 417250 40294 417306 40350
rect 417374 40294 417430 40350
rect 417498 40294 417554 40350
rect 417622 40294 417678 40350
rect 417250 40170 417306 40226
rect 417374 40170 417430 40226
rect 417498 40170 417554 40226
rect 417622 40170 417678 40226
rect 417250 40046 417306 40102
rect 417374 40046 417430 40102
rect 417498 40046 417554 40102
rect 417622 40046 417678 40102
rect 417250 39922 417306 39978
rect 417374 39922 417430 39978
rect 417498 39922 417554 39978
rect 417622 39922 417678 39978
rect 417250 22294 417306 22350
rect 417374 22294 417430 22350
rect 417498 22294 417554 22350
rect 417622 22294 417678 22350
rect 417250 22170 417306 22226
rect 417374 22170 417430 22226
rect 417498 22170 417554 22226
rect 417622 22170 417678 22226
rect 417250 22046 417306 22102
rect 417374 22046 417430 22102
rect 417498 22046 417554 22102
rect 417622 22046 417678 22102
rect 417250 21922 417306 21978
rect 417374 21922 417430 21978
rect 417498 21922 417554 21978
rect 417622 21922 417678 21978
rect 417250 4294 417306 4350
rect 417374 4294 417430 4350
rect 417498 4294 417554 4350
rect 417622 4294 417678 4350
rect 417250 4170 417306 4226
rect 417374 4170 417430 4226
rect 417498 4170 417554 4226
rect 417622 4170 417678 4226
rect 417250 4046 417306 4102
rect 417374 4046 417430 4102
rect 417498 4046 417554 4102
rect 417622 4046 417678 4102
rect 417250 3922 417306 3978
rect 417374 3922 417430 3978
rect 417498 3922 417554 3978
rect 417622 3922 417678 3978
rect 417250 -216 417306 -160
rect 417374 -216 417430 -160
rect 417498 -216 417554 -160
rect 417622 -216 417678 -160
rect 417250 -340 417306 -284
rect 417374 -340 417430 -284
rect 417498 -340 417554 -284
rect 417622 -340 417678 -284
rect 417250 -464 417306 -408
rect 417374 -464 417430 -408
rect 417498 -464 417554 -408
rect 417622 -464 417678 -408
rect 417250 -588 417306 -532
rect 417374 -588 417430 -532
rect 417498 -588 417554 -532
rect 417622 -588 417678 -532
rect 420970 208294 421026 208350
rect 421094 208294 421150 208350
rect 421218 208294 421274 208350
rect 421342 208294 421398 208350
rect 420970 208170 421026 208226
rect 421094 208170 421150 208226
rect 421218 208170 421274 208226
rect 421342 208170 421398 208226
rect 420970 208046 421026 208102
rect 421094 208046 421150 208102
rect 421218 208046 421274 208102
rect 421342 208046 421398 208102
rect 420970 207922 421026 207978
rect 421094 207922 421150 207978
rect 421218 207922 421274 207978
rect 421342 207922 421398 207978
rect 434918 208294 434974 208350
rect 435042 208294 435098 208350
rect 434918 208170 434974 208226
rect 435042 208170 435098 208226
rect 434918 208046 434974 208102
rect 435042 208046 435098 208102
rect 434918 207922 434974 207978
rect 435042 207922 435098 207978
rect 438970 208294 439026 208350
rect 439094 208294 439150 208350
rect 439218 208294 439274 208350
rect 439342 208294 439398 208350
rect 438970 208170 439026 208226
rect 439094 208170 439150 208226
rect 439218 208170 439274 208226
rect 439342 208170 439398 208226
rect 438970 208046 439026 208102
rect 439094 208046 439150 208102
rect 439218 208046 439274 208102
rect 439342 208046 439398 208102
rect 438970 207922 439026 207978
rect 439094 207922 439150 207978
rect 439218 207922 439274 207978
rect 439342 207922 439398 207978
rect 420970 190294 421026 190350
rect 421094 190294 421150 190350
rect 421218 190294 421274 190350
rect 421342 190294 421398 190350
rect 420970 190170 421026 190226
rect 421094 190170 421150 190226
rect 421218 190170 421274 190226
rect 421342 190170 421398 190226
rect 420970 190046 421026 190102
rect 421094 190046 421150 190102
rect 421218 190046 421274 190102
rect 421342 190046 421398 190102
rect 420970 189922 421026 189978
rect 421094 189922 421150 189978
rect 421218 189922 421274 189978
rect 421342 189922 421398 189978
rect 420970 172294 421026 172350
rect 421094 172294 421150 172350
rect 421218 172294 421274 172350
rect 421342 172294 421398 172350
rect 420970 172170 421026 172226
rect 421094 172170 421150 172226
rect 421218 172170 421274 172226
rect 421342 172170 421398 172226
rect 420970 172046 421026 172102
rect 421094 172046 421150 172102
rect 421218 172046 421274 172102
rect 421342 172046 421398 172102
rect 420970 171922 421026 171978
rect 421094 171922 421150 171978
rect 421218 171922 421274 171978
rect 421342 171922 421398 171978
rect 420970 154294 421026 154350
rect 421094 154294 421150 154350
rect 421218 154294 421274 154350
rect 421342 154294 421398 154350
rect 420970 154170 421026 154226
rect 421094 154170 421150 154226
rect 421218 154170 421274 154226
rect 421342 154170 421398 154226
rect 420970 154046 421026 154102
rect 421094 154046 421150 154102
rect 421218 154046 421274 154102
rect 421342 154046 421398 154102
rect 420970 153922 421026 153978
rect 421094 153922 421150 153978
rect 421218 153922 421274 153978
rect 421342 153922 421398 153978
rect 420970 136294 421026 136350
rect 421094 136294 421150 136350
rect 421218 136294 421274 136350
rect 421342 136294 421398 136350
rect 420970 136170 421026 136226
rect 421094 136170 421150 136226
rect 421218 136170 421274 136226
rect 421342 136170 421398 136226
rect 420970 136046 421026 136102
rect 421094 136046 421150 136102
rect 421218 136046 421274 136102
rect 421342 136046 421398 136102
rect 420970 135922 421026 135978
rect 421094 135922 421150 135978
rect 421218 135922 421274 135978
rect 421342 135922 421398 135978
rect 420970 118294 421026 118350
rect 421094 118294 421150 118350
rect 421218 118294 421274 118350
rect 421342 118294 421398 118350
rect 420970 118170 421026 118226
rect 421094 118170 421150 118226
rect 421218 118170 421274 118226
rect 421342 118170 421398 118226
rect 420970 118046 421026 118102
rect 421094 118046 421150 118102
rect 421218 118046 421274 118102
rect 421342 118046 421398 118102
rect 420970 117922 421026 117978
rect 421094 117922 421150 117978
rect 421218 117922 421274 117978
rect 421342 117922 421398 117978
rect 420970 100294 421026 100350
rect 421094 100294 421150 100350
rect 421218 100294 421274 100350
rect 421342 100294 421398 100350
rect 420970 100170 421026 100226
rect 421094 100170 421150 100226
rect 421218 100170 421274 100226
rect 421342 100170 421398 100226
rect 420970 100046 421026 100102
rect 421094 100046 421150 100102
rect 421218 100046 421274 100102
rect 421342 100046 421398 100102
rect 420970 99922 421026 99978
rect 421094 99922 421150 99978
rect 421218 99922 421274 99978
rect 421342 99922 421398 99978
rect 420970 82294 421026 82350
rect 421094 82294 421150 82350
rect 421218 82294 421274 82350
rect 421342 82294 421398 82350
rect 420970 82170 421026 82226
rect 421094 82170 421150 82226
rect 421218 82170 421274 82226
rect 421342 82170 421398 82226
rect 420970 82046 421026 82102
rect 421094 82046 421150 82102
rect 421218 82046 421274 82102
rect 421342 82046 421398 82102
rect 420970 81922 421026 81978
rect 421094 81922 421150 81978
rect 421218 81922 421274 81978
rect 421342 81922 421398 81978
rect 420970 64294 421026 64350
rect 421094 64294 421150 64350
rect 421218 64294 421274 64350
rect 421342 64294 421398 64350
rect 420970 64170 421026 64226
rect 421094 64170 421150 64226
rect 421218 64170 421274 64226
rect 421342 64170 421398 64226
rect 420970 64046 421026 64102
rect 421094 64046 421150 64102
rect 421218 64046 421274 64102
rect 421342 64046 421398 64102
rect 420970 63922 421026 63978
rect 421094 63922 421150 63978
rect 421218 63922 421274 63978
rect 421342 63922 421398 63978
rect 420970 46294 421026 46350
rect 421094 46294 421150 46350
rect 421218 46294 421274 46350
rect 421342 46294 421398 46350
rect 420970 46170 421026 46226
rect 421094 46170 421150 46226
rect 421218 46170 421274 46226
rect 421342 46170 421398 46226
rect 420970 46046 421026 46102
rect 421094 46046 421150 46102
rect 421218 46046 421274 46102
rect 421342 46046 421398 46102
rect 420970 45922 421026 45978
rect 421094 45922 421150 45978
rect 421218 45922 421274 45978
rect 421342 45922 421398 45978
rect 420970 28294 421026 28350
rect 421094 28294 421150 28350
rect 421218 28294 421274 28350
rect 421342 28294 421398 28350
rect 420970 28170 421026 28226
rect 421094 28170 421150 28226
rect 421218 28170 421274 28226
rect 421342 28170 421398 28226
rect 420970 28046 421026 28102
rect 421094 28046 421150 28102
rect 421218 28046 421274 28102
rect 421342 28046 421398 28102
rect 420970 27922 421026 27978
rect 421094 27922 421150 27978
rect 421218 27922 421274 27978
rect 421342 27922 421398 27978
rect 420970 10294 421026 10350
rect 421094 10294 421150 10350
rect 421218 10294 421274 10350
rect 421342 10294 421398 10350
rect 420970 10170 421026 10226
rect 421094 10170 421150 10226
rect 421218 10170 421274 10226
rect 421342 10170 421398 10226
rect 420970 10046 421026 10102
rect 421094 10046 421150 10102
rect 421218 10046 421274 10102
rect 421342 10046 421398 10102
rect 420970 9922 421026 9978
rect 421094 9922 421150 9978
rect 421218 9922 421274 9978
rect 421342 9922 421398 9978
rect 420970 -1176 421026 -1120
rect 421094 -1176 421150 -1120
rect 421218 -1176 421274 -1120
rect 421342 -1176 421398 -1120
rect 420970 -1300 421026 -1244
rect 421094 -1300 421150 -1244
rect 421218 -1300 421274 -1244
rect 421342 -1300 421398 -1244
rect 420970 -1424 421026 -1368
rect 421094 -1424 421150 -1368
rect 421218 -1424 421274 -1368
rect 421342 -1424 421398 -1368
rect 420970 -1548 421026 -1492
rect 421094 -1548 421150 -1492
rect 421218 -1548 421274 -1492
rect 421342 -1548 421398 -1492
rect 435250 184294 435306 184350
rect 435374 184294 435430 184350
rect 435498 184294 435554 184350
rect 435622 184294 435678 184350
rect 435250 184170 435306 184226
rect 435374 184170 435430 184226
rect 435498 184170 435554 184226
rect 435622 184170 435678 184226
rect 435250 184046 435306 184102
rect 435374 184046 435430 184102
rect 435498 184046 435554 184102
rect 435622 184046 435678 184102
rect 435250 183922 435306 183978
rect 435374 183922 435430 183978
rect 435498 183922 435554 183978
rect 435622 183922 435678 183978
rect 435250 166294 435306 166350
rect 435374 166294 435430 166350
rect 435498 166294 435554 166350
rect 435622 166294 435678 166350
rect 435250 166170 435306 166226
rect 435374 166170 435430 166226
rect 435498 166170 435554 166226
rect 435622 166170 435678 166226
rect 435250 166046 435306 166102
rect 435374 166046 435430 166102
rect 435498 166046 435554 166102
rect 435622 166046 435678 166102
rect 435250 165922 435306 165978
rect 435374 165922 435430 165978
rect 435498 165922 435554 165978
rect 435622 165922 435678 165978
rect 435250 148294 435306 148350
rect 435374 148294 435430 148350
rect 435498 148294 435554 148350
rect 435622 148294 435678 148350
rect 435250 148170 435306 148226
rect 435374 148170 435430 148226
rect 435498 148170 435554 148226
rect 435622 148170 435678 148226
rect 435250 148046 435306 148102
rect 435374 148046 435430 148102
rect 435498 148046 435554 148102
rect 435622 148046 435678 148102
rect 435250 147922 435306 147978
rect 435374 147922 435430 147978
rect 435498 147922 435554 147978
rect 435622 147922 435678 147978
rect 435250 130294 435306 130350
rect 435374 130294 435430 130350
rect 435498 130294 435554 130350
rect 435622 130294 435678 130350
rect 435250 130170 435306 130226
rect 435374 130170 435430 130226
rect 435498 130170 435554 130226
rect 435622 130170 435678 130226
rect 435250 130046 435306 130102
rect 435374 130046 435430 130102
rect 435498 130046 435554 130102
rect 435622 130046 435678 130102
rect 435250 129922 435306 129978
rect 435374 129922 435430 129978
rect 435498 129922 435554 129978
rect 435622 129922 435678 129978
rect 435250 112294 435306 112350
rect 435374 112294 435430 112350
rect 435498 112294 435554 112350
rect 435622 112294 435678 112350
rect 435250 112170 435306 112226
rect 435374 112170 435430 112226
rect 435498 112170 435554 112226
rect 435622 112170 435678 112226
rect 435250 112046 435306 112102
rect 435374 112046 435430 112102
rect 435498 112046 435554 112102
rect 435622 112046 435678 112102
rect 435250 111922 435306 111978
rect 435374 111922 435430 111978
rect 435498 111922 435554 111978
rect 435622 111922 435678 111978
rect 435250 94294 435306 94350
rect 435374 94294 435430 94350
rect 435498 94294 435554 94350
rect 435622 94294 435678 94350
rect 435250 94170 435306 94226
rect 435374 94170 435430 94226
rect 435498 94170 435554 94226
rect 435622 94170 435678 94226
rect 435250 94046 435306 94102
rect 435374 94046 435430 94102
rect 435498 94046 435554 94102
rect 435622 94046 435678 94102
rect 435250 93922 435306 93978
rect 435374 93922 435430 93978
rect 435498 93922 435554 93978
rect 435622 93922 435678 93978
rect 435250 76294 435306 76350
rect 435374 76294 435430 76350
rect 435498 76294 435554 76350
rect 435622 76294 435678 76350
rect 435250 76170 435306 76226
rect 435374 76170 435430 76226
rect 435498 76170 435554 76226
rect 435622 76170 435678 76226
rect 435250 76046 435306 76102
rect 435374 76046 435430 76102
rect 435498 76046 435554 76102
rect 435622 76046 435678 76102
rect 435250 75922 435306 75978
rect 435374 75922 435430 75978
rect 435498 75922 435554 75978
rect 435622 75922 435678 75978
rect 435250 58294 435306 58350
rect 435374 58294 435430 58350
rect 435498 58294 435554 58350
rect 435622 58294 435678 58350
rect 435250 58170 435306 58226
rect 435374 58170 435430 58226
rect 435498 58170 435554 58226
rect 435622 58170 435678 58226
rect 435250 58046 435306 58102
rect 435374 58046 435430 58102
rect 435498 58046 435554 58102
rect 435622 58046 435678 58102
rect 435250 57922 435306 57978
rect 435374 57922 435430 57978
rect 435498 57922 435554 57978
rect 435622 57922 435678 57978
rect 435250 40294 435306 40350
rect 435374 40294 435430 40350
rect 435498 40294 435554 40350
rect 435622 40294 435678 40350
rect 435250 40170 435306 40226
rect 435374 40170 435430 40226
rect 435498 40170 435554 40226
rect 435622 40170 435678 40226
rect 435250 40046 435306 40102
rect 435374 40046 435430 40102
rect 435498 40046 435554 40102
rect 435622 40046 435678 40102
rect 435250 39922 435306 39978
rect 435374 39922 435430 39978
rect 435498 39922 435554 39978
rect 435622 39922 435678 39978
rect 435250 22294 435306 22350
rect 435374 22294 435430 22350
rect 435498 22294 435554 22350
rect 435622 22294 435678 22350
rect 435250 22170 435306 22226
rect 435374 22170 435430 22226
rect 435498 22170 435554 22226
rect 435622 22170 435678 22226
rect 435250 22046 435306 22102
rect 435374 22046 435430 22102
rect 435498 22046 435554 22102
rect 435622 22046 435678 22102
rect 435250 21922 435306 21978
rect 435374 21922 435430 21978
rect 435498 21922 435554 21978
rect 435622 21922 435678 21978
rect 435250 4294 435306 4350
rect 435374 4294 435430 4350
rect 435498 4294 435554 4350
rect 435622 4294 435678 4350
rect 435250 4170 435306 4226
rect 435374 4170 435430 4226
rect 435498 4170 435554 4226
rect 435622 4170 435678 4226
rect 435250 4046 435306 4102
rect 435374 4046 435430 4102
rect 435498 4046 435554 4102
rect 435622 4046 435678 4102
rect 435250 3922 435306 3978
rect 435374 3922 435430 3978
rect 435498 3922 435554 3978
rect 435622 3922 435678 3978
rect 435250 -216 435306 -160
rect 435374 -216 435430 -160
rect 435498 -216 435554 -160
rect 435622 -216 435678 -160
rect 435250 -340 435306 -284
rect 435374 -340 435430 -284
rect 435498 -340 435554 -284
rect 435622 -340 435678 -284
rect 435250 -464 435306 -408
rect 435374 -464 435430 -408
rect 435498 -464 435554 -408
rect 435622 -464 435678 -408
rect 435250 -588 435306 -532
rect 435374 -588 435430 -532
rect 435498 -588 435554 -532
rect 435622 -588 435678 -532
rect 438970 190294 439026 190350
rect 439094 190294 439150 190350
rect 439218 190294 439274 190350
rect 439342 190294 439398 190350
rect 438970 190170 439026 190226
rect 439094 190170 439150 190226
rect 439218 190170 439274 190226
rect 439342 190170 439398 190226
rect 438970 190046 439026 190102
rect 439094 190046 439150 190102
rect 439218 190046 439274 190102
rect 439342 190046 439398 190102
rect 438970 189922 439026 189978
rect 439094 189922 439150 189978
rect 439218 189922 439274 189978
rect 439342 189922 439398 189978
rect 438970 172294 439026 172350
rect 439094 172294 439150 172350
rect 439218 172294 439274 172350
rect 439342 172294 439398 172350
rect 438970 172170 439026 172226
rect 439094 172170 439150 172226
rect 439218 172170 439274 172226
rect 439342 172170 439398 172226
rect 438970 172046 439026 172102
rect 439094 172046 439150 172102
rect 439218 172046 439274 172102
rect 439342 172046 439398 172102
rect 438970 171922 439026 171978
rect 439094 171922 439150 171978
rect 439218 171922 439274 171978
rect 439342 171922 439398 171978
rect 438970 154294 439026 154350
rect 439094 154294 439150 154350
rect 439218 154294 439274 154350
rect 439342 154294 439398 154350
rect 438970 154170 439026 154226
rect 439094 154170 439150 154226
rect 439218 154170 439274 154226
rect 439342 154170 439398 154226
rect 438970 154046 439026 154102
rect 439094 154046 439150 154102
rect 439218 154046 439274 154102
rect 439342 154046 439398 154102
rect 438970 153922 439026 153978
rect 439094 153922 439150 153978
rect 439218 153922 439274 153978
rect 439342 153922 439398 153978
rect 438970 136294 439026 136350
rect 439094 136294 439150 136350
rect 439218 136294 439274 136350
rect 439342 136294 439398 136350
rect 438970 136170 439026 136226
rect 439094 136170 439150 136226
rect 439218 136170 439274 136226
rect 439342 136170 439398 136226
rect 438970 136046 439026 136102
rect 439094 136046 439150 136102
rect 439218 136046 439274 136102
rect 439342 136046 439398 136102
rect 438970 135922 439026 135978
rect 439094 135922 439150 135978
rect 439218 135922 439274 135978
rect 439342 135922 439398 135978
rect 438970 118294 439026 118350
rect 439094 118294 439150 118350
rect 439218 118294 439274 118350
rect 439342 118294 439398 118350
rect 438970 118170 439026 118226
rect 439094 118170 439150 118226
rect 439218 118170 439274 118226
rect 439342 118170 439398 118226
rect 438970 118046 439026 118102
rect 439094 118046 439150 118102
rect 439218 118046 439274 118102
rect 439342 118046 439398 118102
rect 438970 117922 439026 117978
rect 439094 117922 439150 117978
rect 439218 117922 439274 117978
rect 439342 117922 439398 117978
rect 438970 100294 439026 100350
rect 439094 100294 439150 100350
rect 439218 100294 439274 100350
rect 439342 100294 439398 100350
rect 438970 100170 439026 100226
rect 439094 100170 439150 100226
rect 439218 100170 439274 100226
rect 439342 100170 439398 100226
rect 438970 100046 439026 100102
rect 439094 100046 439150 100102
rect 439218 100046 439274 100102
rect 439342 100046 439398 100102
rect 438970 99922 439026 99978
rect 439094 99922 439150 99978
rect 439218 99922 439274 99978
rect 439342 99922 439398 99978
rect 438970 82294 439026 82350
rect 439094 82294 439150 82350
rect 439218 82294 439274 82350
rect 439342 82294 439398 82350
rect 438970 82170 439026 82226
rect 439094 82170 439150 82226
rect 439218 82170 439274 82226
rect 439342 82170 439398 82226
rect 438970 82046 439026 82102
rect 439094 82046 439150 82102
rect 439218 82046 439274 82102
rect 439342 82046 439398 82102
rect 438970 81922 439026 81978
rect 439094 81922 439150 81978
rect 439218 81922 439274 81978
rect 439342 81922 439398 81978
rect 438970 64294 439026 64350
rect 439094 64294 439150 64350
rect 439218 64294 439274 64350
rect 439342 64294 439398 64350
rect 438970 64170 439026 64226
rect 439094 64170 439150 64226
rect 439218 64170 439274 64226
rect 439342 64170 439398 64226
rect 438970 64046 439026 64102
rect 439094 64046 439150 64102
rect 439218 64046 439274 64102
rect 439342 64046 439398 64102
rect 438970 63922 439026 63978
rect 439094 63922 439150 63978
rect 439218 63922 439274 63978
rect 439342 63922 439398 63978
rect 438970 46294 439026 46350
rect 439094 46294 439150 46350
rect 439218 46294 439274 46350
rect 439342 46294 439398 46350
rect 438970 46170 439026 46226
rect 439094 46170 439150 46226
rect 439218 46170 439274 46226
rect 439342 46170 439398 46226
rect 438970 46046 439026 46102
rect 439094 46046 439150 46102
rect 439218 46046 439274 46102
rect 439342 46046 439398 46102
rect 438970 45922 439026 45978
rect 439094 45922 439150 45978
rect 439218 45922 439274 45978
rect 439342 45922 439398 45978
rect 438970 28294 439026 28350
rect 439094 28294 439150 28350
rect 439218 28294 439274 28350
rect 439342 28294 439398 28350
rect 438970 28170 439026 28226
rect 439094 28170 439150 28226
rect 439218 28170 439274 28226
rect 439342 28170 439398 28226
rect 438970 28046 439026 28102
rect 439094 28046 439150 28102
rect 439218 28046 439274 28102
rect 439342 28046 439398 28102
rect 438970 27922 439026 27978
rect 439094 27922 439150 27978
rect 439218 27922 439274 27978
rect 439342 27922 439398 27978
rect 438970 10294 439026 10350
rect 439094 10294 439150 10350
rect 439218 10294 439274 10350
rect 439342 10294 439398 10350
rect 438970 10170 439026 10226
rect 439094 10170 439150 10226
rect 439218 10170 439274 10226
rect 439342 10170 439398 10226
rect 438970 10046 439026 10102
rect 439094 10046 439150 10102
rect 439218 10046 439274 10102
rect 439342 10046 439398 10102
rect 438970 9922 439026 9978
rect 439094 9922 439150 9978
rect 439218 9922 439274 9978
rect 439342 9922 439398 9978
rect 438970 -1176 439026 -1120
rect 439094 -1176 439150 -1120
rect 439218 -1176 439274 -1120
rect 439342 -1176 439398 -1120
rect 438970 -1300 439026 -1244
rect 439094 -1300 439150 -1244
rect 439218 -1300 439274 -1244
rect 439342 -1300 439398 -1244
rect 438970 -1424 439026 -1368
rect 439094 -1424 439150 -1368
rect 439218 -1424 439274 -1368
rect 439342 -1424 439398 -1368
rect 438970 -1548 439026 -1492
rect 439094 -1548 439150 -1492
rect 439218 -1548 439274 -1492
rect 439342 -1548 439398 -1492
rect 453250 202294 453306 202350
rect 453374 202294 453430 202350
rect 453498 202294 453554 202350
rect 453622 202294 453678 202350
rect 453250 202170 453306 202226
rect 453374 202170 453430 202226
rect 453498 202170 453554 202226
rect 453622 202170 453678 202226
rect 453250 202046 453306 202102
rect 453374 202046 453430 202102
rect 453498 202046 453554 202102
rect 453622 202046 453678 202102
rect 453250 201922 453306 201978
rect 453374 201922 453430 201978
rect 453498 201922 453554 201978
rect 453622 201922 453678 201978
rect 453250 184294 453306 184350
rect 453374 184294 453430 184350
rect 453498 184294 453554 184350
rect 453622 184294 453678 184350
rect 453250 184170 453306 184226
rect 453374 184170 453430 184226
rect 453498 184170 453554 184226
rect 453622 184170 453678 184226
rect 453250 184046 453306 184102
rect 453374 184046 453430 184102
rect 453498 184046 453554 184102
rect 453622 184046 453678 184102
rect 453250 183922 453306 183978
rect 453374 183922 453430 183978
rect 453498 183922 453554 183978
rect 453622 183922 453678 183978
rect 453250 166294 453306 166350
rect 453374 166294 453430 166350
rect 453498 166294 453554 166350
rect 453622 166294 453678 166350
rect 453250 166170 453306 166226
rect 453374 166170 453430 166226
rect 453498 166170 453554 166226
rect 453622 166170 453678 166226
rect 453250 166046 453306 166102
rect 453374 166046 453430 166102
rect 453498 166046 453554 166102
rect 453622 166046 453678 166102
rect 453250 165922 453306 165978
rect 453374 165922 453430 165978
rect 453498 165922 453554 165978
rect 453622 165922 453678 165978
rect 453250 148294 453306 148350
rect 453374 148294 453430 148350
rect 453498 148294 453554 148350
rect 453622 148294 453678 148350
rect 453250 148170 453306 148226
rect 453374 148170 453430 148226
rect 453498 148170 453554 148226
rect 453622 148170 453678 148226
rect 453250 148046 453306 148102
rect 453374 148046 453430 148102
rect 453498 148046 453554 148102
rect 453622 148046 453678 148102
rect 453250 147922 453306 147978
rect 453374 147922 453430 147978
rect 453498 147922 453554 147978
rect 453622 147922 453678 147978
rect 453250 130294 453306 130350
rect 453374 130294 453430 130350
rect 453498 130294 453554 130350
rect 453622 130294 453678 130350
rect 453250 130170 453306 130226
rect 453374 130170 453430 130226
rect 453498 130170 453554 130226
rect 453622 130170 453678 130226
rect 453250 130046 453306 130102
rect 453374 130046 453430 130102
rect 453498 130046 453554 130102
rect 453622 130046 453678 130102
rect 453250 129922 453306 129978
rect 453374 129922 453430 129978
rect 453498 129922 453554 129978
rect 453622 129922 453678 129978
rect 453250 112294 453306 112350
rect 453374 112294 453430 112350
rect 453498 112294 453554 112350
rect 453622 112294 453678 112350
rect 453250 112170 453306 112226
rect 453374 112170 453430 112226
rect 453498 112170 453554 112226
rect 453622 112170 453678 112226
rect 453250 112046 453306 112102
rect 453374 112046 453430 112102
rect 453498 112046 453554 112102
rect 453622 112046 453678 112102
rect 453250 111922 453306 111978
rect 453374 111922 453430 111978
rect 453498 111922 453554 111978
rect 453622 111922 453678 111978
rect 453250 94294 453306 94350
rect 453374 94294 453430 94350
rect 453498 94294 453554 94350
rect 453622 94294 453678 94350
rect 453250 94170 453306 94226
rect 453374 94170 453430 94226
rect 453498 94170 453554 94226
rect 453622 94170 453678 94226
rect 453250 94046 453306 94102
rect 453374 94046 453430 94102
rect 453498 94046 453554 94102
rect 453622 94046 453678 94102
rect 453250 93922 453306 93978
rect 453374 93922 453430 93978
rect 453498 93922 453554 93978
rect 453622 93922 453678 93978
rect 453250 76294 453306 76350
rect 453374 76294 453430 76350
rect 453498 76294 453554 76350
rect 453622 76294 453678 76350
rect 453250 76170 453306 76226
rect 453374 76170 453430 76226
rect 453498 76170 453554 76226
rect 453622 76170 453678 76226
rect 453250 76046 453306 76102
rect 453374 76046 453430 76102
rect 453498 76046 453554 76102
rect 453622 76046 453678 76102
rect 453250 75922 453306 75978
rect 453374 75922 453430 75978
rect 453498 75922 453554 75978
rect 453622 75922 453678 75978
rect 453250 58294 453306 58350
rect 453374 58294 453430 58350
rect 453498 58294 453554 58350
rect 453622 58294 453678 58350
rect 453250 58170 453306 58226
rect 453374 58170 453430 58226
rect 453498 58170 453554 58226
rect 453622 58170 453678 58226
rect 453250 58046 453306 58102
rect 453374 58046 453430 58102
rect 453498 58046 453554 58102
rect 453622 58046 453678 58102
rect 453250 57922 453306 57978
rect 453374 57922 453430 57978
rect 453498 57922 453554 57978
rect 453622 57922 453678 57978
rect 453250 40294 453306 40350
rect 453374 40294 453430 40350
rect 453498 40294 453554 40350
rect 453622 40294 453678 40350
rect 453250 40170 453306 40226
rect 453374 40170 453430 40226
rect 453498 40170 453554 40226
rect 453622 40170 453678 40226
rect 453250 40046 453306 40102
rect 453374 40046 453430 40102
rect 453498 40046 453554 40102
rect 453622 40046 453678 40102
rect 453250 39922 453306 39978
rect 453374 39922 453430 39978
rect 453498 39922 453554 39978
rect 453622 39922 453678 39978
rect 453250 22294 453306 22350
rect 453374 22294 453430 22350
rect 453498 22294 453554 22350
rect 453622 22294 453678 22350
rect 453250 22170 453306 22226
rect 453374 22170 453430 22226
rect 453498 22170 453554 22226
rect 453622 22170 453678 22226
rect 453250 22046 453306 22102
rect 453374 22046 453430 22102
rect 453498 22046 453554 22102
rect 453622 22046 453678 22102
rect 453250 21922 453306 21978
rect 453374 21922 453430 21978
rect 453498 21922 453554 21978
rect 453622 21922 453678 21978
rect 453250 4294 453306 4350
rect 453374 4294 453430 4350
rect 453498 4294 453554 4350
rect 453622 4294 453678 4350
rect 453250 4170 453306 4226
rect 453374 4170 453430 4226
rect 453498 4170 453554 4226
rect 453622 4170 453678 4226
rect 453250 4046 453306 4102
rect 453374 4046 453430 4102
rect 453498 4046 453554 4102
rect 453622 4046 453678 4102
rect 453250 3922 453306 3978
rect 453374 3922 453430 3978
rect 453498 3922 453554 3978
rect 453622 3922 453678 3978
rect 453250 -216 453306 -160
rect 453374 -216 453430 -160
rect 453498 -216 453554 -160
rect 453622 -216 453678 -160
rect 453250 -340 453306 -284
rect 453374 -340 453430 -284
rect 453498 -340 453554 -284
rect 453622 -340 453678 -284
rect 453250 -464 453306 -408
rect 453374 -464 453430 -408
rect 453498 -464 453554 -408
rect 453622 -464 453678 -408
rect 453250 -588 453306 -532
rect 453374 -588 453430 -532
rect 453498 -588 453554 -532
rect 453622 -588 453678 -532
rect 456970 208294 457026 208350
rect 457094 208294 457150 208350
rect 457218 208294 457274 208350
rect 457342 208294 457398 208350
rect 456970 208170 457026 208226
rect 457094 208170 457150 208226
rect 457218 208170 457274 208226
rect 457342 208170 457398 208226
rect 456970 208046 457026 208102
rect 457094 208046 457150 208102
rect 457218 208046 457274 208102
rect 457342 208046 457398 208102
rect 456970 207922 457026 207978
rect 457094 207922 457150 207978
rect 457218 207922 457274 207978
rect 457342 207922 457398 207978
rect 465638 208294 465694 208350
rect 465762 208294 465818 208350
rect 465638 208170 465694 208226
rect 465762 208170 465818 208226
rect 465638 208046 465694 208102
rect 465762 208046 465818 208102
rect 465638 207922 465694 207978
rect 465762 207922 465818 207978
rect 456970 190294 457026 190350
rect 457094 190294 457150 190350
rect 457218 190294 457274 190350
rect 457342 190294 457398 190350
rect 456970 190170 457026 190226
rect 457094 190170 457150 190226
rect 457218 190170 457274 190226
rect 457342 190170 457398 190226
rect 456970 190046 457026 190102
rect 457094 190046 457150 190102
rect 457218 190046 457274 190102
rect 457342 190046 457398 190102
rect 456970 189922 457026 189978
rect 457094 189922 457150 189978
rect 457218 189922 457274 189978
rect 457342 189922 457398 189978
rect 456970 172294 457026 172350
rect 457094 172294 457150 172350
rect 457218 172294 457274 172350
rect 457342 172294 457398 172350
rect 456970 172170 457026 172226
rect 457094 172170 457150 172226
rect 457218 172170 457274 172226
rect 457342 172170 457398 172226
rect 456970 172046 457026 172102
rect 457094 172046 457150 172102
rect 457218 172046 457274 172102
rect 457342 172046 457398 172102
rect 456970 171922 457026 171978
rect 457094 171922 457150 171978
rect 457218 171922 457274 171978
rect 457342 171922 457398 171978
rect 456970 154294 457026 154350
rect 457094 154294 457150 154350
rect 457218 154294 457274 154350
rect 457342 154294 457398 154350
rect 456970 154170 457026 154226
rect 457094 154170 457150 154226
rect 457218 154170 457274 154226
rect 457342 154170 457398 154226
rect 456970 154046 457026 154102
rect 457094 154046 457150 154102
rect 457218 154046 457274 154102
rect 457342 154046 457398 154102
rect 456970 153922 457026 153978
rect 457094 153922 457150 153978
rect 457218 153922 457274 153978
rect 457342 153922 457398 153978
rect 456970 136294 457026 136350
rect 457094 136294 457150 136350
rect 457218 136294 457274 136350
rect 457342 136294 457398 136350
rect 456970 136170 457026 136226
rect 457094 136170 457150 136226
rect 457218 136170 457274 136226
rect 457342 136170 457398 136226
rect 456970 136046 457026 136102
rect 457094 136046 457150 136102
rect 457218 136046 457274 136102
rect 457342 136046 457398 136102
rect 456970 135922 457026 135978
rect 457094 135922 457150 135978
rect 457218 135922 457274 135978
rect 457342 135922 457398 135978
rect 456970 118294 457026 118350
rect 457094 118294 457150 118350
rect 457218 118294 457274 118350
rect 457342 118294 457398 118350
rect 456970 118170 457026 118226
rect 457094 118170 457150 118226
rect 457218 118170 457274 118226
rect 457342 118170 457398 118226
rect 456970 118046 457026 118102
rect 457094 118046 457150 118102
rect 457218 118046 457274 118102
rect 457342 118046 457398 118102
rect 456970 117922 457026 117978
rect 457094 117922 457150 117978
rect 457218 117922 457274 117978
rect 457342 117922 457398 117978
rect 456970 100294 457026 100350
rect 457094 100294 457150 100350
rect 457218 100294 457274 100350
rect 457342 100294 457398 100350
rect 456970 100170 457026 100226
rect 457094 100170 457150 100226
rect 457218 100170 457274 100226
rect 457342 100170 457398 100226
rect 456970 100046 457026 100102
rect 457094 100046 457150 100102
rect 457218 100046 457274 100102
rect 457342 100046 457398 100102
rect 456970 99922 457026 99978
rect 457094 99922 457150 99978
rect 457218 99922 457274 99978
rect 457342 99922 457398 99978
rect 456970 82294 457026 82350
rect 457094 82294 457150 82350
rect 457218 82294 457274 82350
rect 457342 82294 457398 82350
rect 456970 82170 457026 82226
rect 457094 82170 457150 82226
rect 457218 82170 457274 82226
rect 457342 82170 457398 82226
rect 456970 82046 457026 82102
rect 457094 82046 457150 82102
rect 457218 82046 457274 82102
rect 457342 82046 457398 82102
rect 456970 81922 457026 81978
rect 457094 81922 457150 81978
rect 457218 81922 457274 81978
rect 457342 81922 457398 81978
rect 456970 64294 457026 64350
rect 457094 64294 457150 64350
rect 457218 64294 457274 64350
rect 457342 64294 457398 64350
rect 456970 64170 457026 64226
rect 457094 64170 457150 64226
rect 457218 64170 457274 64226
rect 457342 64170 457398 64226
rect 456970 64046 457026 64102
rect 457094 64046 457150 64102
rect 457218 64046 457274 64102
rect 457342 64046 457398 64102
rect 456970 63922 457026 63978
rect 457094 63922 457150 63978
rect 457218 63922 457274 63978
rect 457342 63922 457398 63978
rect 456970 46294 457026 46350
rect 457094 46294 457150 46350
rect 457218 46294 457274 46350
rect 457342 46294 457398 46350
rect 456970 46170 457026 46226
rect 457094 46170 457150 46226
rect 457218 46170 457274 46226
rect 457342 46170 457398 46226
rect 456970 46046 457026 46102
rect 457094 46046 457150 46102
rect 457218 46046 457274 46102
rect 457342 46046 457398 46102
rect 456970 45922 457026 45978
rect 457094 45922 457150 45978
rect 457218 45922 457274 45978
rect 457342 45922 457398 45978
rect 456970 28294 457026 28350
rect 457094 28294 457150 28350
rect 457218 28294 457274 28350
rect 457342 28294 457398 28350
rect 456970 28170 457026 28226
rect 457094 28170 457150 28226
rect 457218 28170 457274 28226
rect 457342 28170 457398 28226
rect 456970 28046 457026 28102
rect 457094 28046 457150 28102
rect 457218 28046 457274 28102
rect 457342 28046 457398 28102
rect 456970 27922 457026 27978
rect 457094 27922 457150 27978
rect 457218 27922 457274 27978
rect 457342 27922 457398 27978
rect 456970 10294 457026 10350
rect 457094 10294 457150 10350
rect 457218 10294 457274 10350
rect 457342 10294 457398 10350
rect 456970 10170 457026 10226
rect 457094 10170 457150 10226
rect 457218 10170 457274 10226
rect 457342 10170 457398 10226
rect 456970 10046 457026 10102
rect 457094 10046 457150 10102
rect 457218 10046 457274 10102
rect 457342 10046 457398 10102
rect 456970 9922 457026 9978
rect 457094 9922 457150 9978
rect 457218 9922 457274 9978
rect 457342 9922 457398 9978
rect 456970 -1176 457026 -1120
rect 457094 -1176 457150 -1120
rect 457218 -1176 457274 -1120
rect 457342 -1176 457398 -1120
rect 456970 -1300 457026 -1244
rect 457094 -1300 457150 -1244
rect 457218 -1300 457274 -1244
rect 457342 -1300 457398 -1244
rect 456970 -1424 457026 -1368
rect 457094 -1424 457150 -1368
rect 457218 -1424 457274 -1368
rect 457342 -1424 457398 -1368
rect 456970 -1548 457026 -1492
rect 457094 -1548 457150 -1492
rect 457218 -1548 457274 -1492
rect 457342 -1548 457398 -1492
rect 471250 202294 471306 202350
rect 471374 202294 471430 202350
rect 471498 202294 471554 202350
rect 471622 202294 471678 202350
rect 471250 202170 471306 202226
rect 471374 202170 471430 202226
rect 471498 202170 471554 202226
rect 471622 202170 471678 202226
rect 471250 202046 471306 202102
rect 471374 202046 471430 202102
rect 471498 202046 471554 202102
rect 471622 202046 471678 202102
rect 471250 201922 471306 201978
rect 471374 201922 471430 201978
rect 471498 201922 471554 201978
rect 471622 201922 471678 201978
rect 471250 184294 471306 184350
rect 471374 184294 471430 184350
rect 471498 184294 471554 184350
rect 471622 184294 471678 184350
rect 471250 184170 471306 184226
rect 471374 184170 471430 184226
rect 471498 184170 471554 184226
rect 471622 184170 471678 184226
rect 471250 184046 471306 184102
rect 471374 184046 471430 184102
rect 471498 184046 471554 184102
rect 471622 184046 471678 184102
rect 471250 183922 471306 183978
rect 471374 183922 471430 183978
rect 471498 183922 471554 183978
rect 471622 183922 471678 183978
rect 471250 166294 471306 166350
rect 471374 166294 471430 166350
rect 471498 166294 471554 166350
rect 471622 166294 471678 166350
rect 471250 166170 471306 166226
rect 471374 166170 471430 166226
rect 471498 166170 471554 166226
rect 471622 166170 471678 166226
rect 471250 166046 471306 166102
rect 471374 166046 471430 166102
rect 471498 166046 471554 166102
rect 471622 166046 471678 166102
rect 471250 165922 471306 165978
rect 471374 165922 471430 165978
rect 471498 165922 471554 165978
rect 471622 165922 471678 165978
rect 471250 148294 471306 148350
rect 471374 148294 471430 148350
rect 471498 148294 471554 148350
rect 471622 148294 471678 148350
rect 471250 148170 471306 148226
rect 471374 148170 471430 148226
rect 471498 148170 471554 148226
rect 471622 148170 471678 148226
rect 471250 148046 471306 148102
rect 471374 148046 471430 148102
rect 471498 148046 471554 148102
rect 471622 148046 471678 148102
rect 471250 147922 471306 147978
rect 471374 147922 471430 147978
rect 471498 147922 471554 147978
rect 471622 147922 471678 147978
rect 471250 130294 471306 130350
rect 471374 130294 471430 130350
rect 471498 130294 471554 130350
rect 471622 130294 471678 130350
rect 471250 130170 471306 130226
rect 471374 130170 471430 130226
rect 471498 130170 471554 130226
rect 471622 130170 471678 130226
rect 471250 130046 471306 130102
rect 471374 130046 471430 130102
rect 471498 130046 471554 130102
rect 471622 130046 471678 130102
rect 471250 129922 471306 129978
rect 471374 129922 471430 129978
rect 471498 129922 471554 129978
rect 471622 129922 471678 129978
rect 471250 112294 471306 112350
rect 471374 112294 471430 112350
rect 471498 112294 471554 112350
rect 471622 112294 471678 112350
rect 471250 112170 471306 112226
rect 471374 112170 471430 112226
rect 471498 112170 471554 112226
rect 471622 112170 471678 112226
rect 471250 112046 471306 112102
rect 471374 112046 471430 112102
rect 471498 112046 471554 112102
rect 471622 112046 471678 112102
rect 471250 111922 471306 111978
rect 471374 111922 471430 111978
rect 471498 111922 471554 111978
rect 471622 111922 471678 111978
rect 471250 94294 471306 94350
rect 471374 94294 471430 94350
rect 471498 94294 471554 94350
rect 471622 94294 471678 94350
rect 471250 94170 471306 94226
rect 471374 94170 471430 94226
rect 471498 94170 471554 94226
rect 471622 94170 471678 94226
rect 471250 94046 471306 94102
rect 471374 94046 471430 94102
rect 471498 94046 471554 94102
rect 471622 94046 471678 94102
rect 471250 93922 471306 93978
rect 471374 93922 471430 93978
rect 471498 93922 471554 93978
rect 471622 93922 471678 93978
rect 471250 76294 471306 76350
rect 471374 76294 471430 76350
rect 471498 76294 471554 76350
rect 471622 76294 471678 76350
rect 471250 76170 471306 76226
rect 471374 76170 471430 76226
rect 471498 76170 471554 76226
rect 471622 76170 471678 76226
rect 471250 76046 471306 76102
rect 471374 76046 471430 76102
rect 471498 76046 471554 76102
rect 471622 76046 471678 76102
rect 471250 75922 471306 75978
rect 471374 75922 471430 75978
rect 471498 75922 471554 75978
rect 471622 75922 471678 75978
rect 471250 58294 471306 58350
rect 471374 58294 471430 58350
rect 471498 58294 471554 58350
rect 471622 58294 471678 58350
rect 471250 58170 471306 58226
rect 471374 58170 471430 58226
rect 471498 58170 471554 58226
rect 471622 58170 471678 58226
rect 471250 58046 471306 58102
rect 471374 58046 471430 58102
rect 471498 58046 471554 58102
rect 471622 58046 471678 58102
rect 471250 57922 471306 57978
rect 471374 57922 471430 57978
rect 471498 57922 471554 57978
rect 471622 57922 471678 57978
rect 471250 40294 471306 40350
rect 471374 40294 471430 40350
rect 471498 40294 471554 40350
rect 471622 40294 471678 40350
rect 471250 40170 471306 40226
rect 471374 40170 471430 40226
rect 471498 40170 471554 40226
rect 471622 40170 471678 40226
rect 471250 40046 471306 40102
rect 471374 40046 471430 40102
rect 471498 40046 471554 40102
rect 471622 40046 471678 40102
rect 471250 39922 471306 39978
rect 471374 39922 471430 39978
rect 471498 39922 471554 39978
rect 471622 39922 471678 39978
rect 471250 22294 471306 22350
rect 471374 22294 471430 22350
rect 471498 22294 471554 22350
rect 471622 22294 471678 22350
rect 471250 22170 471306 22226
rect 471374 22170 471430 22226
rect 471498 22170 471554 22226
rect 471622 22170 471678 22226
rect 471250 22046 471306 22102
rect 471374 22046 471430 22102
rect 471498 22046 471554 22102
rect 471622 22046 471678 22102
rect 471250 21922 471306 21978
rect 471374 21922 471430 21978
rect 471498 21922 471554 21978
rect 471622 21922 471678 21978
rect 471250 4294 471306 4350
rect 471374 4294 471430 4350
rect 471498 4294 471554 4350
rect 471622 4294 471678 4350
rect 471250 4170 471306 4226
rect 471374 4170 471430 4226
rect 471498 4170 471554 4226
rect 471622 4170 471678 4226
rect 471250 4046 471306 4102
rect 471374 4046 471430 4102
rect 471498 4046 471554 4102
rect 471622 4046 471678 4102
rect 471250 3922 471306 3978
rect 471374 3922 471430 3978
rect 471498 3922 471554 3978
rect 471622 3922 471678 3978
rect 471250 -216 471306 -160
rect 471374 -216 471430 -160
rect 471498 -216 471554 -160
rect 471622 -216 471678 -160
rect 471250 -340 471306 -284
rect 471374 -340 471430 -284
rect 471498 -340 471554 -284
rect 471622 -340 471678 -284
rect 471250 -464 471306 -408
rect 471374 -464 471430 -408
rect 471498 -464 471554 -408
rect 471622 -464 471678 -408
rect 471250 -588 471306 -532
rect 471374 -588 471430 -532
rect 471498 -588 471554 -532
rect 471622 -588 471678 -532
rect 474970 208294 475026 208350
rect 475094 208294 475150 208350
rect 475218 208294 475274 208350
rect 475342 208294 475398 208350
rect 474970 208170 475026 208226
rect 475094 208170 475150 208226
rect 475218 208170 475274 208226
rect 475342 208170 475398 208226
rect 474970 208046 475026 208102
rect 475094 208046 475150 208102
rect 475218 208046 475274 208102
rect 475342 208046 475398 208102
rect 474970 207922 475026 207978
rect 475094 207922 475150 207978
rect 475218 207922 475274 207978
rect 475342 207922 475398 207978
rect 474970 190294 475026 190350
rect 475094 190294 475150 190350
rect 475218 190294 475274 190350
rect 475342 190294 475398 190350
rect 474970 190170 475026 190226
rect 475094 190170 475150 190226
rect 475218 190170 475274 190226
rect 475342 190170 475398 190226
rect 474970 190046 475026 190102
rect 475094 190046 475150 190102
rect 475218 190046 475274 190102
rect 475342 190046 475398 190102
rect 474970 189922 475026 189978
rect 475094 189922 475150 189978
rect 475218 189922 475274 189978
rect 475342 189922 475398 189978
rect 474970 172294 475026 172350
rect 475094 172294 475150 172350
rect 475218 172294 475274 172350
rect 475342 172294 475398 172350
rect 474970 172170 475026 172226
rect 475094 172170 475150 172226
rect 475218 172170 475274 172226
rect 475342 172170 475398 172226
rect 474970 172046 475026 172102
rect 475094 172046 475150 172102
rect 475218 172046 475274 172102
rect 475342 172046 475398 172102
rect 474970 171922 475026 171978
rect 475094 171922 475150 171978
rect 475218 171922 475274 171978
rect 475342 171922 475398 171978
rect 474970 154294 475026 154350
rect 475094 154294 475150 154350
rect 475218 154294 475274 154350
rect 475342 154294 475398 154350
rect 474970 154170 475026 154226
rect 475094 154170 475150 154226
rect 475218 154170 475274 154226
rect 475342 154170 475398 154226
rect 474970 154046 475026 154102
rect 475094 154046 475150 154102
rect 475218 154046 475274 154102
rect 475342 154046 475398 154102
rect 474970 153922 475026 153978
rect 475094 153922 475150 153978
rect 475218 153922 475274 153978
rect 475342 153922 475398 153978
rect 474970 136294 475026 136350
rect 475094 136294 475150 136350
rect 475218 136294 475274 136350
rect 475342 136294 475398 136350
rect 474970 136170 475026 136226
rect 475094 136170 475150 136226
rect 475218 136170 475274 136226
rect 475342 136170 475398 136226
rect 474970 136046 475026 136102
rect 475094 136046 475150 136102
rect 475218 136046 475274 136102
rect 475342 136046 475398 136102
rect 474970 135922 475026 135978
rect 475094 135922 475150 135978
rect 475218 135922 475274 135978
rect 475342 135922 475398 135978
rect 474970 118294 475026 118350
rect 475094 118294 475150 118350
rect 475218 118294 475274 118350
rect 475342 118294 475398 118350
rect 474970 118170 475026 118226
rect 475094 118170 475150 118226
rect 475218 118170 475274 118226
rect 475342 118170 475398 118226
rect 474970 118046 475026 118102
rect 475094 118046 475150 118102
rect 475218 118046 475274 118102
rect 475342 118046 475398 118102
rect 474970 117922 475026 117978
rect 475094 117922 475150 117978
rect 475218 117922 475274 117978
rect 475342 117922 475398 117978
rect 474970 100294 475026 100350
rect 475094 100294 475150 100350
rect 475218 100294 475274 100350
rect 475342 100294 475398 100350
rect 474970 100170 475026 100226
rect 475094 100170 475150 100226
rect 475218 100170 475274 100226
rect 475342 100170 475398 100226
rect 474970 100046 475026 100102
rect 475094 100046 475150 100102
rect 475218 100046 475274 100102
rect 475342 100046 475398 100102
rect 474970 99922 475026 99978
rect 475094 99922 475150 99978
rect 475218 99922 475274 99978
rect 475342 99922 475398 99978
rect 474970 82294 475026 82350
rect 475094 82294 475150 82350
rect 475218 82294 475274 82350
rect 475342 82294 475398 82350
rect 474970 82170 475026 82226
rect 475094 82170 475150 82226
rect 475218 82170 475274 82226
rect 475342 82170 475398 82226
rect 474970 82046 475026 82102
rect 475094 82046 475150 82102
rect 475218 82046 475274 82102
rect 475342 82046 475398 82102
rect 474970 81922 475026 81978
rect 475094 81922 475150 81978
rect 475218 81922 475274 81978
rect 475342 81922 475398 81978
rect 474970 64294 475026 64350
rect 475094 64294 475150 64350
rect 475218 64294 475274 64350
rect 475342 64294 475398 64350
rect 474970 64170 475026 64226
rect 475094 64170 475150 64226
rect 475218 64170 475274 64226
rect 475342 64170 475398 64226
rect 474970 64046 475026 64102
rect 475094 64046 475150 64102
rect 475218 64046 475274 64102
rect 475342 64046 475398 64102
rect 474970 63922 475026 63978
rect 475094 63922 475150 63978
rect 475218 63922 475274 63978
rect 475342 63922 475398 63978
rect 474970 46294 475026 46350
rect 475094 46294 475150 46350
rect 475218 46294 475274 46350
rect 475342 46294 475398 46350
rect 474970 46170 475026 46226
rect 475094 46170 475150 46226
rect 475218 46170 475274 46226
rect 475342 46170 475398 46226
rect 474970 46046 475026 46102
rect 475094 46046 475150 46102
rect 475218 46046 475274 46102
rect 475342 46046 475398 46102
rect 474970 45922 475026 45978
rect 475094 45922 475150 45978
rect 475218 45922 475274 45978
rect 475342 45922 475398 45978
rect 474970 28294 475026 28350
rect 475094 28294 475150 28350
rect 475218 28294 475274 28350
rect 475342 28294 475398 28350
rect 474970 28170 475026 28226
rect 475094 28170 475150 28226
rect 475218 28170 475274 28226
rect 475342 28170 475398 28226
rect 474970 28046 475026 28102
rect 475094 28046 475150 28102
rect 475218 28046 475274 28102
rect 475342 28046 475398 28102
rect 474970 27922 475026 27978
rect 475094 27922 475150 27978
rect 475218 27922 475274 27978
rect 475342 27922 475398 27978
rect 474970 10294 475026 10350
rect 475094 10294 475150 10350
rect 475218 10294 475274 10350
rect 475342 10294 475398 10350
rect 474970 10170 475026 10226
rect 475094 10170 475150 10226
rect 475218 10170 475274 10226
rect 475342 10170 475398 10226
rect 474970 10046 475026 10102
rect 475094 10046 475150 10102
rect 475218 10046 475274 10102
rect 475342 10046 475398 10102
rect 474970 9922 475026 9978
rect 475094 9922 475150 9978
rect 475218 9922 475274 9978
rect 475342 9922 475398 9978
rect 474970 -1176 475026 -1120
rect 475094 -1176 475150 -1120
rect 475218 -1176 475274 -1120
rect 475342 -1176 475398 -1120
rect 474970 -1300 475026 -1244
rect 475094 -1300 475150 -1244
rect 475218 -1300 475274 -1244
rect 475342 -1300 475398 -1244
rect 474970 -1424 475026 -1368
rect 475094 -1424 475150 -1368
rect 475218 -1424 475274 -1368
rect 475342 -1424 475398 -1368
rect 474970 -1548 475026 -1492
rect 475094 -1548 475150 -1492
rect 475218 -1548 475274 -1492
rect 475342 -1548 475398 -1492
rect 489250 202294 489306 202350
rect 489374 202294 489430 202350
rect 489498 202294 489554 202350
rect 489622 202294 489678 202350
rect 489250 202170 489306 202226
rect 489374 202170 489430 202226
rect 489498 202170 489554 202226
rect 489622 202170 489678 202226
rect 489250 202046 489306 202102
rect 489374 202046 489430 202102
rect 489498 202046 489554 202102
rect 489622 202046 489678 202102
rect 489250 201922 489306 201978
rect 489374 201922 489430 201978
rect 489498 201922 489554 201978
rect 489622 201922 489678 201978
rect 489250 184294 489306 184350
rect 489374 184294 489430 184350
rect 489498 184294 489554 184350
rect 489622 184294 489678 184350
rect 489250 184170 489306 184226
rect 489374 184170 489430 184226
rect 489498 184170 489554 184226
rect 489622 184170 489678 184226
rect 489250 184046 489306 184102
rect 489374 184046 489430 184102
rect 489498 184046 489554 184102
rect 489622 184046 489678 184102
rect 489250 183922 489306 183978
rect 489374 183922 489430 183978
rect 489498 183922 489554 183978
rect 489622 183922 489678 183978
rect 489250 166294 489306 166350
rect 489374 166294 489430 166350
rect 489498 166294 489554 166350
rect 489622 166294 489678 166350
rect 489250 166170 489306 166226
rect 489374 166170 489430 166226
rect 489498 166170 489554 166226
rect 489622 166170 489678 166226
rect 489250 166046 489306 166102
rect 489374 166046 489430 166102
rect 489498 166046 489554 166102
rect 489622 166046 489678 166102
rect 489250 165922 489306 165978
rect 489374 165922 489430 165978
rect 489498 165922 489554 165978
rect 489622 165922 489678 165978
rect 489250 148294 489306 148350
rect 489374 148294 489430 148350
rect 489498 148294 489554 148350
rect 489622 148294 489678 148350
rect 489250 148170 489306 148226
rect 489374 148170 489430 148226
rect 489498 148170 489554 148226
rect 489622 148170 489678 148226
rect 489250 148046 489306 148102
rect 489374 148046 489430 148102
rect 489498 148046 489554 148102
rect 489622 148046 489678 148102
rect 489250 147922 489306 147978
rect 489374 147922 489430 147978
rect 489498 147922 489554 147978
rect 489622 147922 489678 147978
rect 489250 130294 489306 130350
rect 489374 130294 489430 130350
rect 489498 130294 489554 130350
rect 489622 130294 489678 130350
rect 489250 130170 489306 130226
rect 489374 130170 489430 130226
rect 489498 130170 489554 130226
rect 489622 130170 489678 130226
rect 489250 130046 489306 130102
rect 489374 130046 489430 130102
rect 489498 130046 489554 130102
rect 489622 130046 489678 130102
rect 489250 129922 489306 129978
rect 489374 129922 489430 129978
rect 489498 129922 489554 129978
rect 489622 129922 489678 129978
rect 489250 112294 489306 112350
rect 489374 112294 489430 112350
rect 489498 112294 489554 112350
rect 489622 112294 489678 112350
rect 489250 112170 489306 112226
rect 489374 112170 489430 112226
rect 489498 112170 489554 112226
rect 489622 112170 489678 112226
rect 489250 112046 489306 112102
rect 489374 112046 489430 112102
rect 489498 112046 489554 112102
rect 489622 112046 489678 112102
rect 489250 111922 489306 111978
rect 489374 111922 489430 111978
rect 489498 111922 489554 111978
rect 489622 111922 489678 111978
rect 489250 94294 489306 94350
rect 489374 94294 489430 94350
rect 489498 94294 489554 94350
rect 489622 94294 489678 94350
rect 489250 94170 489306 94226
rect 489374 94170 489430 94226
rect 489498 94170 489554 94226
rect 489622 94170 489678 94226
rect 489250 94046 489306 94102
rect 489374 94046 489430 94102
rect 489498 94046 489554 94102
rect 489622 94046 489678 94102
rect 489250 93922 489306 93978
rect 489374 93922 489430 93978
rect 489498 93922 489554 93978
rect 489622 93922 489678 93978
rect 489250 76294 489306 76350
rect 489374 76294 489430 76350
rect 489498 76294 489554 76350
rect 489622 76294 489678 76350
rect 489250 76170 489306 76226
rect 489374 76170 489430 76226
rect 489498 76170 489554 76226
rect 489622 76170 489678 76226
rect 489250 76046 489306 76102
rect 489374 76046 489430 76102
rect 489498 76046 489554 76102
rect 489622 76046 489678 76102
rect 489250 75922 489306 75978
rect 489374 75922 489430 75978
rect 489498 75922 489554 75978
rect 489622 75922 489678 75978
rect 489250 58294 489306 58350
rect 489374 58294 489430 58350
rect 489498 58294 489554 58350
rect 489622 58294 489678 58350
rect 489250 58170 489306 58226
rect 489374 58170 489430 58226
rect 489498 58170 489554 58226
rect 489622 58170 489678 58226
rect 489250 58046 489306 58102
rect 489374 58046 489430 58102
rect 489498 58046 489554 58102
rect 489622 58046 489678 58102
rect 489250 57922 489306 57978
rect 489374 57922 489430 57978
rect 489498 57922 489554 57978
rect 489622 57922 489678 57978
rect 489250 40294 489306 40350
rect 489374 40294 489430 40350
rect 489498 40294 489554 40350
rect 489622 40294 489678 40350
rect 489250 40170 489306 40226
rect 489374 40170 489430 40226
rect 489498 40170 489554 40226
rect 489622 40170 489678 40226
rect 489250 40046 489306 40102
rect 489374 40046 489430 40102
rect 489498 40046 489554 40102
rect 489622 40046 489678 40102
rect 489250 39922 489306 39978
rect 489374 39922 489430 39978
rect 489498 39922 489554 39978
rect 489622 39922 489678 39978
rect 489250 22294 489306 22350
rect 489374 22294 489430 22350
rect 489498 22294 489554 22350
rect 489622 22294 489678 22350
rect 489250 22170 489306 22226
rect 489374 22170 489430 22226
rect 489498 22170 489554 22226
rect 489622 22170 489678 22226
rect 489250 22046 489306 22102
rect 489374 22046 489430 22102
rect 489498 22046 489554 22102
rect 489622 22046 489678 22102
rect 489250 21922 489306 21978
rect 489374 21922 489430 21978
rect 489498 21922 489554 21978
rect 489622 21922 489678 21978
rect 489250 4294 489306 4350
rect 489374 4294 489430 4350
rect 489498 4294 489554 4350
rect 489622 4294 489678 4350
rect 489250 4170 489306 4226
rect 489374 4170 489430 4226
rect 489498 4170 489554 4226
rect 489622 4170 489678 4226
rect 489250 4046 489306 4102
rect 489374 4046 489430 4102
rect 489498 4046 489554 4102
rect 489622 4046 489678 4102
rect 489250 3922 489306 3978
rect 489374 3922 489430 3978
rect 489498 3922 489554 3978
rect 489622 3922 489678 3978
rect 489250 -216 489306 -160
rect 489374 -216 489430 -160
rect 489498 -216 489554 -160
rect 489622 -216 489678 -160
rect 489250 -340 489306 -284
rect 489374 -340 489430 -284
rect 489498 -340 489554 -284
rect 489622 -340 489678 -284
rect 489250 -464 489306 -408
rect 489374 -464 489430 -408
rect 489498 -464 489554 -408
rect 489622 -464 489678 -408
rect 489250 -588 489306 -532
rect 489374 -588 489430 -532
rect 489498 -588 489554 -532
rect 489622 -588 489678 -532
rect 492970 208294 493026 208350
rect 493094 208294 493150 208350
rect 493218 208294 493274 208350
rect 493342 208294 493398 208350
rect 492970 208170 493026 208226
rect 493094 208170 493150 208226
rect 493218 208170 493274 208226
rect 493342 208170 493398 208226
rect 492970 208046 493026 208102
rect 493094 208046 493150 208102
rect 493218 208046 493274 208102
rect 493342 208046 493398 208102
rect 492970 207922 493026 207978
rect 493094 207922 493150 207978
rect 493218 207922 493274 207978
rect 493342 207922 493398 207978
rect 496358 208294 496414 208350
rect 496482 208294 496538 208350
rect 496358 208170 496414 208226
rect 496482 208170 496538 208226
rect 496358 208046 496414 208102
rect 496482 208046 496538 208102
rect 496358 207922 496414 207978
rect 496482 207922 496538 207978
rect 492970 190294 493026 190350
rect 493094 190294 493150 190350
rect 493218 190294 493274 190350
rect 493342 190294 493398 190350
rect 492970 190170 493026 190226
rect 493094 190170 493150 190226
rect 493218 190170 493274 190226
rect 493342 190170 493398 190226
rect 492970 190046 493026 190102
rect 493094 190046 493150 190102
rect 493218 190046 493274 190102
rect 493342 190046 493398 190102
rect 492970 189922 493026 189978
rect 493094 189922 493150 189978
rect 493218 189922 493274 189978
rect 493342 189922 493398 189978
rect 492970 172294 493026 172350
rect 493094 172294 493150 172350
rect 493218 172294 493274 172350
rect 493342 172294 493398 172350
rect 492970 172170 493026 172226
rect 493094 172170 493150 172226
rect 493218 172170 493274 172226
rect 493342 172170 493398 172226
rect 492970 172046 493026 172102
rect 493094 172046 493150 172102
rect 493218 172046 493274 172102
rect 493342 172046 493398 172102
rect 492970 171922 493026 171978
rect 493094 171922 493150 171978
rect 493218 171922 493274 171978
rect 493342 171922 493398 171978
rect 492970 154294 493026 154350
rect 493094 154294 493150 154350
rect 493218 154294 493274 154350
rect 493342 154294 493398 154350
rect 492970 154170 493026 154226
rect 493094 154170 493150 154226
rect 493218 154170 493274 154226
rect 493342 154170 493398 154226
rect 492970 154046 493026 154102
rect 493094 154046 493150 154102
rect 493218 154046 493274 154102
rect 493342 154046 493398 154102
rect 492970 153922 493026 153978
rect 493094 153922 493150 153978
rect 493218 153922 493274 153978
rect 493342 153922 493398 153978
rect 492970 136294 493026 136350
rect 493094 136294 493150 136350
rect 493218 136294 493274 136350
rect 493342 136294 493398 136350
rect 492970 136170 493026 136226
rect 493094 136170 493150 136226
rect 493218 136170 493274 136226
rect 493342 136170 493398 136226
rect 492970 136046 493026 136102
rect 493094 136046 493150 136102
rect 493218 136046 493274 136102
rect 493342 136046 493398 136102
rect 492970 135922 493026 135978
rect 493094 135922 493150 135978
rect 493218 135922 493274 135978
rect 493342 135922 493398 135978
rect 492970 118294 493026 118350
rect 493094 118294 493150 118350
rect 493218 118294 493274 118350
rect 493342 118294 493398 118350
rect 492970 118170 493026 118226
rect 493094 118170 493150 118226
rect 493218 118170 493274 118226
rect 493342 118170 493398 118226
rect 492970 118046 493026 118102
rect 493094 118046 493150 118102
rect 493218 118046 493274 118102
rect 493342 118046 493398 118102
rect 492970 117922 493026 117978
rect 493094 117922 493150 117978
rect 493218 117922 493274 117978
rect 493342 117922 493398 117978
rect 492970 100294 493026 100350
rect 493094 100294 493150 100350
rect 493218 100294 493274 100350
rect 493342 100294 493398 100350
rect 492970 100170 493026 100226
rect 493094 100170 493150 100226
rect 493218 100170 493274 100226
rect 493342 100170 493398 100226
rect 492970 100046 493026 100102
rect 493094 100046 493150 100102
rect 493218 100046 493274 100102
rect 493342 100046 493398 100102
rect 492970 99922 493026 99978
rect 493094 99922 493150 99978
rect 493218 99922 493274 99978
rect 493342 99922 493398 99978
rect 492970 82294 493026 82350
rect 493094 82294 493150 82350
rect 493218 82294 493274 82350
rect 493342 82294 493398 82350
rect 492970 82170 493026 82226
rect 493094 82170 493150 82226
rect 493218 82170 493274 82226
rect 493342 82170 493398 82226
rect 492970 82046 493026 82102
rect 493094 82046 493150 82102
rect 493218 82046 493274 82102
rect 493342 82046 493398 82102
rect 492970 81922 493026 81978
rect 493094 81922 493150 81978
rect 493218 81922 493274 81978
rect 493342 81922 493398 81978
rect 492970 64294 493026 64350
rect 493094 64294 493150 64350
rect 493218 64294 493274 64350
rect 493342 64294 493398 64350
rect 492970 64170 493026 64226
rect 493094 64170 493150 64226
rect 493218 64170 493274 64226
rect 493342 64170 493398 64226
rect 492970 64046 493026 64102
rect 493094 64046 493150 64102
rect 493218 64046 493274 64102
rect 493342 64046 493398 64102
rect 492970 63922 493026 63978
rect 493094 63922 493150 63978
rect 493218 63922 493274 63978
rect 493342 63922 493398 63978
rect 492970 46294 493026 46350
rect 493094 46294 493150 46350
rect 493218 46294 493274 46350
rect 493342 46294 493398 46350
rect 492970 46170 493026 46226
rect 493094 46170 493150 46226
rect 493218 46170 493274 46226
rect 493342 46170 493398 46226
rect 492970 46046 493026 46102
rect 493094 46046 493150 46102
rect 493218 46046 493274 46102
rect 493342 46046 493398 46102
rect 492970 45922 493026 45978
rect 493094 45922 493150 45978
rect 493218 45922 493274 45978
rect 493342 45922 493398 45978
rect 492970 28294 493026 28350
rect 493094 28294 493150 28350
rect 493218 28294 493274 28350
rect 493342 28294 493398 28350
rect 492970 28170 493026 28226
rect 493094 28170 493150 28226
rect 493218 28170 493274 28226
rect 493342 28170 493398 28226
rect 492970 28046 493026 28102
rect 493094 28046 493150 28102
rect 493218 28046 493274 28102
rect 493342 28046 493398 28102
rect 492970 27922 493026 27978
rect 493094 27922 493150 27978
rect 493218 27922 493274 27978
rect 493342 27922 493398 27978
rect 492970 10294 493026 10350
rect 493094 10294 493150 10350
rect 493218 10294 493274 10350
rect 493342 10294 493398 10350
rect 492970 10170 493026 10226
rect 493094 10170 493150 10226
rect 493218 10170 493274 10226
rect 493342 10170 493398 10226
rect 492970 10046 493026 10102
rect 493094 10046 493150 10102
rect 493218 10046 493274 10102
rect 493342 10046 493398 10102
rect 492970 9922 493026 9978
rect 493094 9922 493150 9978
rect 493218 9922 493274 9978
rect 493342 9922 493398 9978
rect 492970 -1176 493026 -1120
rect 493094 -1176 493150 -1120
rect 493218 -1176 493274 -1120
rect 493342 -1176 493398 -1120
rect 492970 -1300 493026 -1244
rect 493094 -1300 493150 -1244
rect 493218 -1300 493274 -1244
rect 493342 -1300 493398 -1244
rect 492970 -1424 493026 -1368
rect 493094 -1424 493150 -1368
rect 493218 -1424 493274 -1368
rect 493342 -1424 493398 -1368
rect 492970 -1548 493026 -1492
rect 493094 -1548 493150 -1492
rect 493218 -1548 493274 -1492
rect 493342 -1548 493398 -1492
rect 507250 202294 507306 202350
rect 507374 202294 507430 202350
rect 507498 202294 507554 202350
rect 507622 202294 507678 202350
rect 507250 202170 507306 202226
rect 507374 202170 507430 202226
rect 507498 202170 507554 202226
rect 507622 202170 507678 202226
rect 507250 202046 507306 202102
rect 507374 202046 507430 202102
rect 507498 202046 507554 202102
rect 507622 202046 507678 202102
rect 507250 201922 507306 201978
rect 507374 201922 507430 201978
rect 507498 201922 507554 201978
rect 507622 201922 507678 201978
rect 507250 184294 507306 184350
rect 507374 184294 507430 184350
rect 507498 184294 507554 184350
rect 507622 184294 507678 184350
rect 507250 184170 507306 184226
rect 507374 184170 507430 184226
rect 507498 184170 507554 184226
rect 507622 184170 507678 184226
rect 507250 184046 507306 184102
rect 507374 184046 507430 184102
rect 507498 184046 507554 184102
rect 507622 184046 507678 184102
rect 507250 183922 507306 183978
rect 507374 183922 507430 183978
rect 507498 183922 507554 183978
rect 507622 183922 507678 183978
rect 507250 166294 507306 166350
rect 507374 166294 507430 166350
rect 507498 166294 507554 166350
rect 507622 166294 507678 166350
rect 507250 166170 507306 166226
rect 507374 166170 507430 166226
rect 507498 166170 507554 166226
rect 507622 166170 507678 166226
rect 507250 166046 507306 166102
rect 507374 166046 507430 166102
rect 507498 166046 507554 166102
rect 507622 166046 507678 166102
rect 507250 165922 507306 165978
rect 507374 165922 507430 165978
rect 507498 165922 507554 165978
rect 507622 165922 507678 165978
rect 507250 148294 507306 148350
rect 507374 148294 507430 148350
rect 507498 148294 507554 148350
rect 507622 148294 507678 148350
rect 507250 148170 507306 148226
rect 507374 148170 507430 148226
rect 507498 148170 507554 148226
rect 507622 148170 507678 148226
rect 507250 148046 507306 148102
rect 507374 148046 507430 148102
rect 507498 148046 507554 148102
rect 507622 148046 507678 148102
rect 507250 147922 507306 147978
rect 507374 147922 507430 147978
rect 507498 147922 507554 147978
rect 507622 147922 507678 147978
rect 507250 130294 507306 130350
rect 507374 130294 507430 130350
rect 507498 130294 507554 130350
rect 507622 130294 507678 130350
rect 507250 130170 507306 130226
rect 507374 130170 507430 130226
rect 507498 130170 507554 130226
rect 507622 130170 507678 130226
rect 507250 130046 507306 130102
rect 507374 130046 507430 130102
rect 507498 130046 507554 130102
rect 507622 130046 507678 130102
rect 507250 129922 507306 129978
rect 507374 129922 507430 129978
rect 507498 129922 507554 129978
rect 507622 129922 507678 129978
rect 507250 112294 507306 112350
rect 507374 112294 507430 112350
rect 507498 112294 507554 112350
rect 507622 112294 507678 112350
rect 507250 112170 507306 112226
rect 507374 112170 507430 112226
rect 507498 112170 507554 112226
rect 507622 112170 507678 112226
rect 507250 112046 507306 112102
rect 507374 112046 507430 112102
rect 507498 112046 507554 112102
rect 507622 112046 507678 112102
rect 507250 111922 507306 111978
rect 507374 111922 507430 111978
rect 507498 111922 507554 111978
rect 507622 111922 507678 111978
rect 507250 94294 507306 94350
rect 507374 94294 507430 94350
rect 507498 94294 507554 94350
rect 507622 94294 507678 94350
rect 507250 94170 507306 94226
rect 507374 94170 507430 94226
rect 507498 94170 507554 94226
rect 507622 94170 507678 94226
rect 507250 94046 507306 94102
rect 507374 94046 507430 94102
rect 507498 94046 507554 94102
rect 507622 94046 507678 94102
rect 507250 93922 507306 93978
rect 507374 93922 507430 93978
rect 507498 93922 507554 93978
rect 507622 93922 507678 93978
rect 507250 76294 507306 76350
rect 507374 76294 507430 76350
rect 507498 76294 507554 76350
rect 507622 76294 507678 76350
rect 507250 76170 507306 76226
rect 507374 76170 507430 76226
rect 507498 76170 507554 76226
rect 507622 76170 507678 76226
rect 507250 76046 507306 76102
rect 507374 76046 507430 76102
rect 507498 76046 507554 76102
rect 507622 76046 507678 76102
rect 507250 75922 507306 75978
rect 507374 75922 507430 75978
rect 507498 75922 507554 75978
rect 507622 75922 507678 75978
rect 507250 58294 507306 58350
rect 507374 58294 507430 58350
rect 507498 58294 507554 58350
rect 507622 58294 507678 58350
rect 507250 58170 507306 58226
rect 507374 58170 507430 58226
rect 507498 58170 507554 58226
rect 507622 58170 507678 58226
rect 507250 58046 507306 58102
rect 507374 58046 507430 58102
rect 507498 58046 507554 58102
rect 507622 58046 507678 58102
rect 507250 57922 507306 57978
rect 507374 57922 507430 57978
rect 507498 57922 507554 57978
rect 507622 57922 507678 57978
rect 507250 40294 507306 40350
rect 507374 40294 507430 40350
rect 507498 40294 507554 40350
rect 507622 40294 507678 40350
rect 507250 40170 507306 40226
rect 507374 40170 507430 40226
rect 507498 40170 507554 40226
rect 507622 40170 507678 40226
rect 507250 40046 507306 40102
rect 507374 40046 507430 40102
rect 507498 40046 507554 40102
rect 507622 40046 507678 40102
rect 507250 39922 507306 39978
rect 507374 39922 507430 39978
rect 507498 39922 507554 39978
rect 507622 39922 507678 39978
rect 507250 22294 507306 22350
rect 507374 22294 507430 22350
rect 507498 22294 507554 22350
rect 507622 22294 507678 22350
rect 507250 22170 507306 22226
rect 507374 22170 507430 22226
rect 507498 22170 507554 22226
rect 507622 22170 507678 22226
rect 507250 22046 507306 22102
rect 507374 22046 507430 22102
rect 507498 22046 507554 22102
rect 507622 22046 507678 22102
rect 507250 21922 507306 21978
rect 507374 21922 507430 21978
rect 507498 21922 507554 21978
rect 507622 21922 507678 21978
rect 507250 4294 507306 4350
rect 507374 4294 507430 4350
rect 507498 4294 507554 4350
rect 507622 4294 507678 4350
rect 507250 4170 507306 4226
rect 507374 4170 507430 4226
rect 507498 4170 507554 4226
rect 507622 4170 507678 4226
rect 507250 4046 507306 4102
rect 507374 4046 507430 4102
rect 507498 4046 507554 4102
rect 507622 4046 507678 4102
rect 507250 3922 507306 3978
rect 507374 3922 507430 3978
rect 507498 3922 507554 3978
rect 507622 3922 507678 3978
rect 507250 -216 507306 -160
rect 507374 -216 507430 -160
rect 507498 -216 507554 -160
rect 507622 -216 507678 -160
rect 507250 -340 507306 -284
rect 507374 -340 507430 -284
rect 507498 -340 507554 -284
rect 507622 -340 507678 -284
rect 507250 -464 507306 -408
rect 507374 -464 507430 -408
rect 507498 -464 507554 -408
rect 507622 -464 507678 -408
rect 507250 -588 507306 -532
rect 507374 -588 507430 -532
rect 507498 -588 507554 -532
rect 507622 -588 507678 -532
rect 510970 598116 511026 598172
rect 511094 598116 511150 598172
rect 511218 598116 511274 598172
rect 511342 598116 511398 598172
rect 510970 597992 511026 598048
rect 511094 597992 511150 598048
rect 511218 597992 511274 598048
rect 511342 597992 511398 598048
rect 510970 597868 511026 597924
rect 511094 597868 511150 597924
rect 511218 597868 511274 597924
rect 511342 597868 511398 597924
rect 510970 597744 511026 597800
rect 511094 597744 511150 597800
rect 511218 597744 511274 597800
rect 511342 597744 511398 597800
rect 510970 586294 511026 586350
rect 511094 586294 511150 586350
rect 511218 586294 511274 586350
rect 511342 586294 511398 586350
rect 510970 586170 511026 586226
rect 511094 586170 511150 586226
rect 511218 586170 511274 586226
rect 511342 586170 511398 586226
rect 510970 586046 511026 586102
rect 511094 586046 511150 586102
rect 511218 586046 511274 586102
rect 511342 586046 511398 586102
rect 510970 585922 511026 585978
rect 511094 585922 511150 585978
rect 511218 585922 511274 585978
rect 511342 585922 511398 585978
rect 510970 568294 511026 568350
rect 511094 568294 511150 568350
rect 511218 568294 511274 568350
rect 511342 568294 511398 568350
rect 510970 568170 511026 568226
rect 511094 568170 511150 568226
rect 511218 568170 511274 568226
rect 511342 568170 511398 568226
rect 510970 568046 511026 568102
rect 511094 568046 511150 568102
rect 511218 568046 511274 568102
rect 511342 568046 511398 568102
rect 510970 567922 511026 567978
rect 511094 567922 511150 567978
rect 511218 567922 511274 567978
rect 511342 567922 511398 567978
rect 510970 550294 511026 550350
rect 511094 550294 511150 550350
rect 511218 550294 511274 550350
rect 511342 550294 511398 550350
rect 510970 550170 511026 550226
rect 511094 550170 511150 550226
rect 511218 550170 511274 550226
rect 511342 550170 511398 550226
rect 510970 550046 511026 550102
rect 511094 550046 511150 550102
rect 511218 550046 511274 550102
rect 511342 550046 511398 550102
rect 510970 549922 511026 549978
rect 511094 549922 511150 549978
rect 511218 549922 511274 549978
rect 511342 549922 511398 549978
rect 510970 532294 511026 532350
rect 511094 532294 511150 532350
rect 511218 532294 511274 532350
rect 511342 532294 511398 532350
rect 510970 532170 511026 532226
rect 511094 532170 511150 532226
rect 511218 532170 511274 532226
rect 511342 532170 511398 532226
rect 510970 532046 511026 532102
rect 511094 532046 511150 532102
rect 511218 532046 511274 532102
rect 511342 532046 511398 532102
rect 510970 531922 511026 531978
rect 511094 531922 511150 531978
rect 511218 531922 511274 531978
rect 511342 531922 511398 531978
rect 510970 514294 511026 514350
rect 511094 514294 511150 514350
rect 511218 514294 511274 514350
rect 511342 514294 511398 514350
rect 510970 514170 511026 514226
rect 511094 514170 511150 514226
rect 511218 514170 511274 514226
rect 511342 514170 511398 514226
rect 510970 514046 511026 514102
rect 511094 514046 511150 514102
rect 511218 514046 511274 514102
rect 511342 514046 511398 514102
rect 510970 513922 511026 513978
rect 511094 513922 511150 513978
rect 511218 513922 511274 513978
rect 511342 513922 511398 513978
rect 510970 496294 511026 496350
rect 511094 496294 511150 496350
rect 511218 496294 511274 496350
rect 511342 496294 511398 496350
rect 510970 496170 511026 496226
rect 511094 496170 511150 496226
rect 511218 496170 511274 496226
rect 511342 496170 511398 496226
rect 510970 496046 511026 496102
rect 511094 496046 511150 496102
rect 511218 496046 511274 496102
rect 511342 496046 511398 496102
rect 510970 495922 511026 495978
rect 511094 495922 511150 495978
rect 511218 495922 511274 495978
rect 511342 495922 511398 495978
rect 510970 478294 511026 478350
rect 511094 478294 511150 478350
rect 511218 478294 511274 478350
rect 511342 478294 511398 478350
rect 510970 478170 511026 478226
rect 511094 478170 511150 478226
rect 511218 478170 511274 478226
rect 511342 478170 511398 478226
rect 510970 478046 511026 478102
rect 511094 478046 511150 478102
rect 511218 478046 511274 478102
rect 511342 478046 511398 478102
rect 510970 477922 511026 477978
rect 511094 477922 511150 477978
rect 511218 477922 511274 477978
rect 511342 477922 511398 477978
rect 510970 460294 511026 460350
rect 511094 460294 511150 460350
rect 511218 460294 511274 460350
rect 511342 460294 511398 460350
rect 510970 460170 511026 460226
rect 511094 460170 511150 460226
rect 511218 460170 511274 460226
rect 511342 460170 511398 460226
rect 510970 460046 511026 460102
rect 511094 460046 511150 460102
rect 511218 460046 511274 460102
rect 511342 460046 511398 460102
rect 510970 459922 511026 459978
rect 511094 459922 511150 459978
rect 511218 459922 511274 459978
rect 511342 459922 511398 459978
rect 510970 442294 511026 442350
rect 511094 442294 511150 442350
rect 511218 442294 511274 442350
rect 511342 442294 511398 442350
rect 510970 442170 511026 442226
rect 511094 442170 511150 442226
rect 511218 442170 511274 442226
rect 511342 442170 511398 442226
rect 510970 442046 511026 442102
rect 511094 442046 511150 442102
rect 511218 442046 511274 442102
rect 511342 442046 511398 442102
rect 510970 441922 511026 441978
rect 511094 441922 511150 441978
rect 511218 441922 511274 441978
rect 511342 441922 511398 441978
rect 510970 424294 511026 424350
rect 511094 424294 511150 424350
rect 511218 424294 511274 424350
rect 511342 424294 511398 424350
rect 510970 424170 511026 424226
rect 511094 424170 511150 424226
rect 511218 424170 511274 424226
rect 511342 424170 511398 424226
rect 510970 424046 511026 424102
rect 511094 424046 511150 424102
rect 511218 424046 511274 424102
rect 511342 424046 511398 424102
rect 510970 423922 511026 423978
rect 511094 423922 511150 423978
rect 511218 423922 511274 423978
rect 511342 423922 511398 423978
rect 510970 406294 511026 406350
rect 511094 406294 511150 406350
rect 511218 406294 511274 406350
rect 511342 406294 511398 406350
rect 510970 406170 511026 406226
rect 511094 406170 511150 406226
rect 511218 406170 511274 406226
rect 511342 406170 511398 406226
rect 510970 406046 511026 406102
rect 511094 406046 511150 406102
rect 511218 406046 511274 406102
rect 511342 406046 511398 406102
rect 510970 405922 511026 405978
rect 511094 405922 511150 405978
rect 511218 405922 511274 405978
rect 511342 405922 511398 405978
rect 510970 388294 511026 388350
rect 511094 388294 511150 388350
rect 511218 388294 511274 388350
rect 511342 388294 511398 388350
rect 510970 388170 511026 388226
rect 511094 388170 511150 388226
rect 511218 388170 511274 388226
rect 511342 388170 511398 388226
rect 510970 388046 511026 388102
rect 511094 388046 511150 388102
rect 511218 388046 511274 388102
rect 511342 388046 511398 388102
rect 510970 387922 511026 387978
rect 511094 387922 511150 387978
rect 511218 387922 511274 387978
rect 511342 387922 511398 387978
rect 510970 370294 511026 370350
rect 511094 370294 511150 370350
rect 511218 370294 511274 370350
rect 511342 370294 511398 370350
rect 510970 370170 511026 370226
rect 511094 370170 511150 370226
rect 511218 370170 511274 370226
rect 511342 370170 511398 370226
rect 510970 370046 511026 370102
rect 511094 370046 511150 370102
rect 511218 370046 511274 370102
rect 511342 370046 511398 370102
rect 510970 369922 511026 369978
rect 511094 369922 511150 369978
rect 511218 369922 511274 369978
rect 511342 369922 511398 369978
rect 510970 352294 511026 352350
rect 511094 352294 511150 352350
rect 511218 352294 511274 352350
rect 511342 352294 511398 352350
rect 510970 352170 511026 352226
rect 511094 352170 511150 352226
rect 511218 352170 511274 352226
rect 511342 352170 511398 352226
rect 510970 352046 511026 352102
rect 511094 352046 511150 352102
rect 511218 352046 511274 352102
rect 511342 352046 511398 352102
rect 510970 351922 511026 351978
rect 511094 351922 511150 351978
rect 511218 351922 511274 351978
rect 511342 351922 511398 351978
rect 510970 334294 511026 334350
rect 511094 334294 511150 334350
rect 511218 334294 511274 334350
rect 511342 334294 511398 334350
rect 510970 334170 511026 334226
rect 511094 334170 511150 334226
rect 511218 334170 511274 334226
rect 511342 334170 511398 334226
rect 510970 334046 511026 334102
rect 511094 334046 511150 334102
rect 511218 334046 511274 334102
rect 511342 334046 511398 334102
rect 510970 333922 511026 333978
rect 511094 333922 511150 333978
rect 511218 333922 511274 333978
rect 511342 333922 511398 333978
rect 510970 316294 511026 316350
rect 511094 316294 511150 316350
rect 511218 316294 511274 316350
rect 511342 316294 511398 316350
rect 510970 316170 511026 316226
rect 511094 316170 511150 316226
rect 511218 316170 511274 316226
rect 511342 316170 511398 316226
rect 510970 316046 511026 316102
rect 511094 316046 511150 316102
rect 511218 316046 511274 316102
rect 511342 316046 511398 316102
rect 510970 315922 511026 315978
rect 511094 315922 511150 315978
rect 511218 315922 511274 315978
rect 511342 315922 511398 315978
rect 510970 298294 511026 298350
rect 511094 298294 511150 298350
rect 511218 298294 511274 298350
rect 511342 298294 511398 298350
rect 510970 298170 511026 298226
rect 511094 298170 511150 298226
rect 511218 298170 511274 298226
rect 511342 298170 511398 298226
rect 510970 298046 511026 298102
rect 511094 298046 511150 298102
rect 511218 298046 511274 298102
rect 511342 298046 511398 298102
rect 510970 297922 511026 297978
rect 511094 297922 511150 297978
rect 511218 297922 511274 297978
rect 511342 297922 511398 297978
rect 510970 280294 511026 280350
rect 511094 280294 511150 280350
rect 511218 280294 511274 280350
rect 511342 280294 511398 280350
rect 510970 280170 511026 280226
rect 511094 280170 511150 280226
rect 511218 280170 511274 280226
rect 511342 280170 511398 280226
rect 510970 280046 511026 280102
rect 511094 280046 511150 280102
rect 511218 280046 511274 280102
rect 511342 280046 511398 280102
rect 510970 279922 511026 279978
rect 511094 279922 511150 279978
rect 511218 279922 511274 279978
rect 511342 279922 511398 279978
rect 510970 262294 511026 262350
rect 511094 262294 511150 262350
rect 511218 262294 511274 262350
rect 511342 262294 511398 262350
rect 510970 262170 511026 262226
rect 511094 262170 511150 262226
rect 511218 262170 511274 262226
rect 511342 262170 511398 262226
rect 510970 262046 511026 262102
rect 511094 262046 511150 262102
rect 511218 262046 511274 262102
rect 511342 262046 511398 262102
rect 510970 261922 511026 261978
rect 511094 261922 511150 261978
rect 511218 261922 511274 261978
rect 511342 261922 511398 261978
rect 510970 244294 511026 244350
rect 511094 244294 511150 244350
rect 511218 244294 511274 244350
rect 511342 244294 511398 244350
rect 510970 244170 511026 244226
rect 511094 244170 511150 244226
rect 511218 244170 511274 244226
rect 511342 244170 511398 244226
rect 510970 244046 511026 244102
rect 511094 244046 511150 244102
rect 511218 244046 511274 244102
rect 511342 244046 511398 244102
rect 510970 243922 511026 243978
rect 511094 243922 511150 243978
rect 511218 243922 511274 243978
rect 511342 243922 511398 243978
rect 510970 226294 511026 226350
rect 511094 226294 511150 226350
rect 511218 226294 511274 226350
rect 511342 226294 511398 226350
rect 510970 226170 511026 226226
rect 511094 226170 511150 226226
rect 511218 226170 511274 226226
rect 511342 226170 511398 226226
rect 510970 226046 511026 226102
rect 511094 226046 511150 226102
rect 511218 226046 511274 226102
rect 511342 226046 511398 226102
rect 510970 225922 511026 225978
rect 511094 225922 511150 225978
rect 511218 225922 511274 225978
rect 511342 225922 511398 225978
rect 510970 208294 511026 208350
rect 511094 208294 511150 208350
rect 511218 208294 511274 208350
rect 511342 208294 511398 208350
rect 510970 208170 511026 208226
rect 511094 208170 511150 208226
rect 511218 208170 511274 208226
rect 511342 208170 511398 208226
rect 510970 208046 511026 208102
rect 511094 208046 511150 208102
rect 511218 208046 511274 208102
rect 511342 208046 511398 208102
rect 510970 207922 511026 207978
rect 511094 207922 511150 207978
rect 511218 207922 511274 207978
rect 511342 207922 511398 207978
rect 510970 190294 511026 190350
rect 511094 190294 511150 190350
rect 511218 190294 511274 190350
rect 511342 190294 511398 190350
rect 510970 190170 511026 190226
rect 511094 190170 511150 190226
rect 511218 190170 511274 190226
rect 511342 190170 511398 190226
rect 510970 190046 511026 190102
rect 511094 190046 511150 190102
rect 511218 190046 511274 190102
rect 511342 190046 511398 190102
rect 510970 189922 511026 189978
rect 511094 189922 511150 189978
rect 511218 189922 511274 189978
rect 511342 189922 511398 189978
rect 510970 172294 511026 172350
rect 511094 172294 511150 172350
rect 511218 172294 511274 172350
rect 511342 172294 511398 172350
rect 510970 172170 511026 172226
rect 511094 172170 511150 172226
rect 511218 172170 511274 172226
rect 511342 172170 511398 172226
rect 510970 172046 511026 172102
rect 511094 172046 511150 172102
rect 511218 172046 511274 172102
rect 511342 172046 511398 172102
rect 510970 171922 511026 171978
rect 511094 171922 511150 171978
rect 511218 171922 511274 171978
rect 511342 171922 511398 171978
rect 510970 154294 511026 154350
rect 511094 154294 511150 154350
rect 511218 154294 511274 154350
rect 511342 154294 511398 154350
rect 510970 154170 511026 154226
rect 511094 154170 511150 154226
rect 511218 154170 511274 154226
rect 511342 154170 511398 154226
rect 510970 154046 511026 154102
rect 511094 154046 511150 154102
rect 511218 154046 511274 154102
rect 511342 154046 511398 154102
rect 510970 153922 511026 153978
rect 511094 153922 511150 153978
rect 511218 153922 511274 153978
rect 511342 153922 511398 153978
rect 510970 136294 511026 136350
rect 511094 136294 511150 136350
rect 511218 136294 511274 136350
rect 511342 136294 511398 136350
rect 510970 136170 511026 136226
rect 511094 136170 511150 136226
rect 511218 136170 511274 136226
rect 511342 136170 511398 136226
rect 510970 136046 511026 136102
rect 511094 136046 511150 136102
rect 511218 136046 511274 136102
rect 511342 136046 511398 136102
rect 510970 135922 511026 135978
rect 511094 135922 511150 135978
rect 511218 135922 511274 135978
rect 511342 135922 511398 135978
rect 510970 118294 511026 118350
rect 511094 118294 511150 118350
rect 511218 118294 511274 118350
rect 511342 118294 511398 118350
rect 510970 118170 511026 118226
rect 511094 118170 511150 118226
rect 511218 118170 511274 118226
rect 511342 118170 511398 118226
rect 510970 118046 511026 118102
rect 511094 118046 511150 118102
rect 511218 118046 511274 118102
rect 511342 118046 511398 118102
rect 510970 117922 511026 117978
rect 511094 117922 511150 117978
rect 511218 117922 511274 117978
rect 511342 117922 511398 117978
rect 510970 100294 511026 100350
rect 511094 100294 511150 100350
rect 511218 100294 511274 100350
rect 511342 100294 511398 100350
rect 510970 100170 511026 100226
rect 511094 100170 511150 100226
rect 511218 100170 511274 100226
rect 511342 100170 511398 100226
rect 510970 100046 511026 100102
rect 511094 100046 511150 100102
rect 511218 100046 511274 100102
rect 511342 100046 511398 100102
rect 510970 99922 511026 99978
rect 511094 99922 511150 99978
rect 511218 99922 511274 99978
rect 511342 99922 511398 99978
rect 510970 82294 511026 82350
rect 511094 82294 511150 82350
rect 511218 82294 511274 82350
rect 511342 82294 511398 82350
rect 510970 82170 511026 82226
rect 511094 82170 511150 82226
rect 511218 82170 511274 82226
rect 511342 82170 511398 82226
rect 510970 82046 511026 82102
rect 511094 82046 511150 82102
rect 511218 82046 511274 82102
rect 511342 82046 511398 82102
rect 510970 81922 511026 81978
rect 511094 81922 511150 81978
rect 511218 81922 511274 81978
rect 511342 81922 511398 81978
rect 510970 64294 511026 64350
rect 511094 64294 511150 64350
rect 511218 64294 511274 64350
rect 511342 64294 511398 64350
rect 510970 64170 511026 64226
rect 511094 64170 511150 64226
rect 511218 64170 511274 64226
rect 511342 64170 511398 64226
rect 510970 64046 511026 64102
rect 511094 64046 511150 64102
rect 511218 64046 511274 64102
rect 511342 64046 511398 64102
rect 510970 63922 511026 63978
rect 511094 63922 511150 63978
rect 511218 63922 511274 63978
rect 511342 63922 511398 63978
rect 510970 46294 511026 46350
rect 511094 46294 511150 46350
rect 511218 46294 511274 46350
rect 511342 46294 511398 46350
rect 510970 46170 511026 46226
rect 511094 46170 511150 46226
rect 511218 46170 511274 46226
rect 511342 46170 511398 46226
rect 510970 46046 511026 46102
rect 511094 46046 511150 46102
rect 511218 46046 511274 46102
rect 511342 46046 511398 46102
rect 510970 45922 511026 45978
rect 511094 45922 511150 45978
rect 511218 45922 511274 45978
rect 511342 45922 511398 45978
rect 510970 28294 511026 28350
rect 511094 28294 511150 28350
rect 511218 28294 511274 28350
rect 511342 28294 511398 28350
rect 510970 28170 511026 28226
rect 511094 28170 511150 28226
rect 511218 28170 511274 28226
rect 511342 28170 511398 28226
rect 510970 28046 511026 28102
rect 511094 28046 511150 28102
rect 511218 28046 511274 28102
rect 511342 28046 511398 28102
rect 510970 27922 511026 27978
rect 511094 27922 511150 27978
rect 511218 27922 511274 27978
rect 511342 27922 511398 27978
rect 510970 10294 511026 10350
rect 511094 10294 511150 10350
rect 511218 10294 511274 10350
rect 511342 10294 511398 10350
rect 510970 10170 511026 10226
rect 511094 10170 511150 10226
rect 511218 10170 511274 10226
rect 511342 10170 511398 10226
rect 510970 10046 511026 10102
rect 511094 10046 511150 10102
rect 511218 10046 511274 10102
rect 511342 10046 511398 10102
rect 510970 9922 511026 9978
rect 511094 9922 511150 9978
rect 511218 9922 511274 9978
rect 511342 9922 511398 9978
rect 510970 -1176 511026 -1120
rect 511094 -1176 511150 -1120
rect 511218 -1176 511274 -1120
rect 511342 -1176 511398 -1120
rect 510970 -1300 511026 -1244
rect 511094 -1300 511150 -1244
rect 511218 -1300 511274 -1244
rect 511342 -1300 511398 -1244
rect 510970 -1424 511026 -1368
rect 511094 -1424 511150 -1368
rect 511218 -1424 511274 -1368
rect 511342 -1424 511398 -1368
rect 510970 -1548 511026 -1492
rect 511094 -1548 511150 -1492
rect 511218 -1548 511274 -1492
rect 511342 -1548 511398 -1492
rect 525250 597156 525306 597212
rect 525374 597156 525430 597212
rect 525498 597156 525554 597212
rect 525622 597156 525678 597212
rect 525250 597032 525306 597088
rect 525374 597032 525430 597088
rect 525498 597032 525554 597088
rect 525622 597032 525678 597088
rect 525250 596908 525306 596964
rect 525374 596908 525430 596964
rect 525498 596908 525554 596964
rect 525622 596908 525678 596964
rect 525250 596784 525306 596840
rect 525374 596784 525430 596840
rect 525498 596784 525554 596840
rect 525622 596784 525678 596840
rect 525250 580294 525306 580350
rect 525374 580294 525430 580350
rect 525498 580294 525554 580350
rect 525622 580294 525678 580350
rect 525250 580170 525306 580226
rect 525374 580170 525430 580226
rect 525498 580170 525554 580226
rect 525622 580170 525678 580226
rect 525250 580046 525306 580102
rect 525374 580046 525430 580102
rect 525498 580046 525554 580102
rect 525622 580046 525678 580102
rect 525250 579922 525306 579978
rect 525374 579922 525430 579978
rect 525498 579922 525554 579978
rect 525622 579922 525678 579978
rect 525250 562294 525306 562350
rect 525374 562294 525430 562350
rect 525498 562294 525554 562350
rect 525622 562294 525678 562350
rect 525250 562170 525306 562226
rect 525374 562170 525430 562226
rect 525498 562170 525554 562226
rect 525622 562170 525678 562226
rect 525250 562046 525306 562102
rect 525374 562046 525430 562102
rect 525498 562046 525554 562102
rect 525622 562046 525678 562102
rect 525250 561922 525306 561978
rect 525374 561922 525430 561978
rect 525498 561922 525554 561978
rect 525622 561922 525678 561978
rect 525250 544294 525306 544350
rect 525374 544294 525430 544350
rect 525498 544294 525554 544350
rect 525622 544294 525678 544350
rect 525250 544170 525306 544226
rect 525374 544170 525430 544226
rect 525498 544170 525554 544226
rect 525622 544170 525678 544226
rect 525250 544046 525306 544102
rect 525374 544046 525430 544102
rect 525498 544046 525554 544102
rect 525622 544046 525678 544102
rect 525250 543922 525306 543978
rect 525374 543922 525430 543978
rect 525498 543922 525554 543978
rect 525622 543922 525678 543978
rect 525250 526294 525306 526350
rect 525374 526294 525430 526350
rect 525498 526294 525554 526350
rect 525622 526294 525678 526350
rect 525250 526170 525306 526226
rect 525374 526170 525430 526226
rect 525498 526170 525554 526226
rect 525622 526170 525678 526226
rect 525250 526046 525306 526102
rect 525374 526046 525430 526102
rect 525498 526046 525554 526102
rect 525622 526046 525678 526102
rect 525250 525922 525306 525978
rect 525374 525922 525430 525978
rect 525498 525922 525554 525978
rect 525622 525922 525678 525978
rect 525250 508294 525306 508350
rect 525374 508294 525430 508350
rect 525498 508294 525554 508350
rect 525622 508294 525678 508350
rect 525250 508170 525306 508226
rect 525374 508170 525430 508226
rect 525498 508170 525554 508226
rect 525622 508170 525678 508226
rect 525250 508046 525306 508102
rect 525374 508046 525430 508102
rect 525498 508046 525554 508102
rect 525622 508046 525678 508102
rect 525250 507922 525306 507978
rect 525374 507922 525430 507978
rect 525498 507922 525554 507978
rect 525622 507922 525678 507978
rect 525250 490294 525306 490350
rect 525374 490294 525430 490350
rect 525498 490294 525554 490350
rect 525622 490294 525678 490350
rect 525250 490170 525306 490226
rect 525374 490170 525430 490226
rect 525498 490170 525554 490226
rect 525622 490170 525678 490226
rect 525250 490046 525306 490102
rect 525374 490046 525430 490102
rect 525498 490046 525554 490102
rect 525622 490046 525678 490102
rect 525250 489922 525306 489978
rect 525374 489922 525430 489978
rect 525498 489922 525554 489978
rect 525622 489922 525678 489978
rect 525250 472294 525306 472350
rect 525374 472294 525430 472350
rect 525498 472294 525554 472350
rect 525622 472294 525678 472350
rect 525250 472170 525306 472226
rect 525374 472170 525430 472226
rect 525498 472170 525554 472226
rect 525622 472170 525678 472226
rect 525250 472046 525306 472102
rect 525374 472046 525430 472102
rect 525498 472046 525554 472102
rect 525622 472046 525678 472102
rect 525250 471922 525306 471978
rect 525374 471922 525430 471978
rect 525498 471922 525554 471978
rect 525622 471922 525678 471978
rect 525250 454294 525306 454350
rect 525374 454294 525430 454350
rect 525498 454294 525554 454350
rect 525622 454294 525678 454350
rect 525250 454170 525306 454226
rect 525374 454170 525430 454226
rect 525498 454170 525554 454226
rect 525622 454170 525678 454226
rect 525250 454046 525306 454102
rect 525374 454046 525430 454102
rect 525498 454046 525554 454102
rect 525622 454046 525678 454102
rect 525250 453922 525306 453978
rect 525374 453922 525430 453978
rect 525498 453922 525554 453978
rect 525622 453922 525678 453978
rect 525250 436294 525306 436350
rect 525374 436294 525430 436350
rect 525498 436294 525554 436350
rect 525622 436294 525678 436350
rect 525250 436170 525306 436226
rect 525374 436170 525430 436226
rect 525498 436170 525554 436226
rect 525622 436170 525678 436226
rect 525250 436046 525306 436102
rect 525374 436046 525430 436102
rect 525498 436046 525554 436102
rect 525622 436046 525678 436102
rect 525250 435922 525306 435978
rect 525374 435922 525430 435978
rect 525498 435922 525554 435978
rect 525622 435922 525678 435978
rect 525250 418294 525306 418350
rect 525374 418294 525430 418350
rect 525498 418294 525554 418350
rect 525622 418294 525678 418350
rect 525250 418170 525306 418226
rect 525374 418170 525430 418226
rect 525498 418170 525554 418226
rect 525622 418170 525678 418226
rect 525250 418046 525306 418102
rect 525374 418046 525430 418102
rect 525498 418046 525554 418102
rect 525622 418046 525678 418102
rect 525250 417922 525306 417978
rect 525374 417922 525430 417978
rect 525498 417922 525554 417978
rect 525622 417922 525678 417978
rect 525250 400294 525306 400350
rect 525374 400294 525430 400350
rect 525498 400294 525554 400350
rect 525622 400294 525678 400350
rect 525250 400170 525306 400226
rect 525374 400170 525430 400226
rect 525498 400170 525554 400226
rect 525622 400170 525678 400226
rect 525250 400046 525306 400102
rect 525374 400046 525430 400102
rect 525498 400046 525554 400102
rect 525622 400046 525678 400102
rect 525250 399922 525306 399978
rect 525374 399922 525430 399978
rect 525498 399922 525554 399978
rect 525622 399922 525678 399978
rect 525250 382294 525306 382350
rect 525374 382294 525430 382350
rect 525498 382294 525554 382350
rect 525622 382294 525678 382350
rect 525250 382170 525306 382226
rect 525374 382170 525430 382226
rect 525498 382170 525554 382226
rect 525622 382170 525678 382226
rect 525250 382046 525306 382102
rect 525374 382046 525430 382102
rect 525498 382046 525554 382102
rect 525622 382046 525678 382102
rect 525250 381922 525306 381978
rect 525374 381922 525430 381978
rect 525498 381922 525554 381978
rect 525622 381922 525678 381978
rect 525250 364294 525306 364350
rect 525374 364294 525430 364350
rect 525498 364294 525554 364350
rect 525622 364294 525678 364350
rect 525250 364170 525306 364226
rect 525374 364170 525430 364226
rect 525498 364170 525554 364226
rect 525622 364170 525678 364226
rect 525250 364046 525306 364102
rect 525374 364046 525430 364102
rect 525498 364046 525554 364102
rect 525622 364046 525678 364102
rect 525250 363922 525306 363978
rect 525374 363922 525430 363978
rect 525498 363922 525554 363978
rect 525622 363922 525678 363978
rect 525250 346294 525306 346350
rect 525374 346294 525430 346350
rect 525498 346294 525554 346350
rect 525622 346294 525678 346350
rect 525250 346170 525306 346226
rect 525374 346170 525430 346226
rect 525498 346170 525554 346226
rect 525622 346170 525678 346226
rect 525250 346046 525306 346102
rect 525374 346046 525430 346102
rect 525498 346046 525554 346102
rect 525622 346046 525678 346102
rect 525250 345922 525306 345978
rect 525374 345922 525430 345978
rect 525498 345922 525554 345978
rect 525622 345922 525678 345978
rect 525250 328294 525306 328350
rect 525374 328294 525430 328350
rect 525498 328294 525554 328350
rect 525622 328294 525678 328350
rect 525250 328170 525306 328226
rect 525374 328170 525430 328226
rect 525498 328170 525554 328226
rect 525622 328170 525678 328226
rect 525250 328046 525306 328102
rect 525374 328046 525430 328102
rect 525498 328046 525554 328102
rect 525622 328046 525678 328102
rect 525250 327922 525306 327978
rect 525374 327922 525430 327978
rect 525498 327922 525554 327978
rect 525622 327922 525678 327978
rect 525250 310294 525306 310350
rect 525374 310294 525430 310350
rect 525498 310294 525554 310350
rect 525622 310294 525678 310350
rect 525250 310170 525306 310226
rect 525374 310170 525430 310226
rect 525498 310170 525554 310226
rect 525622 310170 525678 310226
rect 525250 310046 525306 310102
rect 525374 310046 525430 310102
rect 525498 310046 525554 310102
rect 525622 310046 525678 310102
rect 525250 309922 525306 309978
rect 525374 309922 525430 309978
rect 525498 309922 525554 309978
rect 525622 309922 525678 309978
rect 525250 292294 525306 292350
rect 525374 292294 525430 292350
rect 525498 292294 525554 292350
rect 525622 292294 525678 292350
rect 525250 292170 525306 292226
rect 525374 292170 525430 292226
rect 525498 292170 525554 292226
rect 525622 292170 525678 292226
rect 525250 292046 525306 292102
rect 525374 292046 525430 292102
rect 525498 292046 525554 292102
rect 525622 292046 525678 292102
rect 525250 291922 525306 291978
rect 525374 291922 525430 291978
rect 525498 291922 525554 291978
rect 525622 291922 525678 291978
rect 525250 274294 525306 274350
rect 525374 274294 525430 274350
rect 525498 274294 525554 274350
rect 525622 274294 525678 274350
rect 525250 274170 525306 274226
rect 525374 274170 525430 274226
rect 525498 274170 525554 274226
rect 525622 274170 525678 274226
rect 525250 274046 525306 274102
rect 525374 274046 525430 274102
rect 525498 274046 525554 274102
rect 525622 274046 525678 274102
rect 525250 273922 525306 273978
rect 525374 273922 525430 273978
rect 525498 273922 525554 273978
rect 525622 273922 525678 273978
rect 525250 256294 525306 256350
rect 525374 256294 525430 256350
rect 525498 256294 525554 256350
rect 525622 256294 525678 256350
rect 525250 256170 525306 256226
rect 525374 256170 525430 256226
rect 525498 256170 525554 256226
rect 525622 256170 525678 256226
rect 525250 256046 525306 256102
rect 525374 256046 525430 256102
rect 525498 256046 525554 256102
rect 525622 256046 525678 256102
rect 525250 255922 525306 255978
rect 525374 255922 525430 255978
rect 525498 255922 525554 255978
rect 525622 255922 525678 255978
rect 525250 238294 525306 238350
rect 525374 238294 525430 238350
rect 525498 238294 525554 238350
rect 525622 238294 525678 238350
rect 525250 238170 525306 238226
rect 525374 238170 525430 238226
rect 525498 238170 525554 238226
rect 525622 238170 525678 238226
rect 525250 238046 525306 238102
rect 525374 238046 525430 238102
rect 525498 238046 525554 238102
rect 525622 238046 525678 238102
rect 525250 237922 525306 237978
rect 525374 237922 525430 237978
rect 525498 237922 525554 237978
rect 525622 237922 525678 237978
rect 525250 220294 525306 220350
rect 525374 220294 525430 220350
rect 525498 220294 525554 220350
rect 525622 220294 525678 220350
rect 525250 220170 525306 220226
rect 525374 220170 525430 220226
rect 525498 220170 525554 220226
rect 525622 220170 525678 220226
rect 525250 220046 525306 220102
rect 525374 220046 525430 220102
rect 525498 220046 525554 220102
rect 525622 220046 525678 220102
rect 525250 219922 525306 219978
rect 525374 219922 525430 219978
rect 525498 219922 525554 219978
rect 525622 219922 525678 219978
rect 525250 202294 525306 202350
rect 525374 202294 525430 202350
rect 525498 202294 525554 202350
rect 525622 202294 525678 202350
rect 525250 202170 525306 202226
rect 525374 202170 525430 202226
rect 525498 202170 525554 202226
rect 525622 202170 525678 202226
rect 525250 202046 525306 202102
rect 525374 202046 525430 202102
rect 525498 202046 525554 202102
rect 525622 202046 525678 202102
rect 525250 201922 525306 201978
rect 525374 201922 525430 201978
rect 525498 201922 525554 201978
rect 525622 201922 525678 201978
rect 525250 184294 525306 184350
rect 525374 184294 525430 184350
rect 525498 184294 525554 184350
rect 525622 184294 525678 184350
rect 525250 184170 525306 184226
rect 525374 184170 525430 184226
rect 525498 184170 525554 184226
rect 525622 184170 525678 184226
rect 525250 184046 525306 184102
rect 525374 184046 525430 184102
rect 525498 184046 525554 184102
rect 525622 184046 525678 184102
rect 525250 183922 525306 183978
rect 525374 183922 525430 183978
rect 525498 183922 525554 183978
rect 525622 183922 525678 183978
rect 525250 166294 525306 166350
rect 525374 166294 525430 166350
rect 525498 166294 525554 166350
rect 525622 166294 525678 166350
rect 525250 166170 525306 166226
rect 525374 166170 525430 166226
rect 525498 166170 525554 166226
rect 525622 166170 525678 166226
rect 525250 166046 525306 166102
rect 525374 166046 525430 166102
rect 525498 166046 525554 166102
rect 525622 166046 525678 166102
rect 525250 165922 525306 165978
rect 525374 165922 525430 165978
rect 525498 165922 525554 165978
rect 525622 165922 525678 165978
rect 525250 148294 525306 148350
rect 525374 148294 525430 148350
rect 525498 148294 525554 148350
rect 525622 148294 525678 148350
rect 525250 148170 525306 148226
rect 525374 148170 525430 148226
rect 525498 148170 525554 148226
rect 525622 148170 525678 148226
rect 525250 148046 525306 148102
rect 525374 148046 525430 148102
rect 525498 148046 525554 148102
rect 525622 148046 525678 148102
rect 525250 147922 525306 147978
rect 525374 147922 525430 147978
rect 525498 147922 525554 147978
rect 525622 147922 525678 147978
rect 525250 130294 525306 130350
rect 525374 130294 525430 130350
rect 525498 130294 525554 130350
rect 525622 130294 525678 130350
rect 525250 130170 525306 130226
rect 525374 130170 525430 130226
rect 525498 130170 525554 130226
rect 525622 130170 525678 130226
rect 525250 130046 525306 130102
rect 525374 130046 525430 130102
rect 525498 130046 525554 130102
rect 525622 130046 525678 130102
rect 525250 129922 525306 129978
rect 525374 129922 525430 129978
rect 525498 129922 525554 129978
rect 525622 129922 525678 129978
rect 525250 112294 525306 112350
rect 525374 112294 525430 112350
rect 525498 112294 525554 112350
rect 525622 112294 525678 112350
rect 525250 112170 525306 112226
rect 525374 112170 525430 112226
rect 525498 112170 525554 112226
rect 525622 112170 525678 112226
rect 525250 112046 525306 112102
rect 525374 112046 525430 112102
rect 525498 112046 525554 112102
rect 525622 112046 525678 112102
rect 525250 111922 525306 111978
rect 525374 111922 525430 111978
rect 525498 111922 525554 111978
rect 525622 111922 525678 111978
rect 525250 94294 525306 94350
rect 525374 94294 525430 94350
rect 525498 94294 525554 94350
rect 525622 94294 525678 94350
rect 525250 94170 525306 94226
rect 525374 94170 525430 94226
rect 525498 94170 525554 94226
rect 525622 94170 525678 94226
rect 525250 94046 525306 94102
rect 525374 94046 525430 94102
rect 525498 94046 525554 94102
rect 525622 94046 525678 94102
rect 525250 93922 525306 93978
rect 525374 93922 525430 93978
rect 525498 93922 525554 93978
rect 525622 93922 525678 93978
rect 525250 76294 525306 76350
rect 525374 76294 525430 76350
rect 525498 76294 525554 76350
rect 525622 76294 525678 76350
rect 525250 76170 525306 76226
rect 525374 76170 525430 76226
rect 525498 76170 525554 76226
rect 525622 76170 525678 76226
rect 525250 76046 525306 76102
rect 525374 76046 525430 76102
rect 525498 76046 525554 76102
rect 525622 76046 525678 76102
rect 525250 75922 525306 75978
rect 525374 75922 525430 75978
rect 525498 75922 525554 75978
rect 525622 75922 525678 75978
rect 525250 58294 525306 58350
rect 525374 58294 525430 58350
rect 525498 58294 525554 58350
rect 525622 58294 525678 58350
rect 525250 58170 525306 58226
rect 525374 58170 525430 58226
rect 525498 58170 525554 58226
rect 525622 58170 525678 58226
rect 525250 58046 525306 58102
rect 525374 58046 525430 58102
rect 525498 58046 525554 58102
rect 525622 58046 525678 58102
rect 525250 57922 525306 57978
rect 525374 57922 525430 57978
rect 525498 57922 525554 57978
rect 525622 57922 525678 57978
rect 525250 40294 525306 40350
rect 525374 40294 525430 40350
rect 525498 40294 525554 40350
rect 525622 40294 525678 40350
rect 525250 40170 525306 40226
rect 525374 40170 525430 40226
rect 525498 40170 525554 40226
rect 525622 40170 525678 40226
rect 525250 40046 525306 40102
rect 525374 40046 525430 40102
rect 525498 40046 525554 40102
rect 525622 40046 525678 40102
rect 525250 39922 525306 39978
rect 525374 39922 525430 39978
rect 525498 39922 525554 39978
rect 525622 39922 525678 39978
rect 525250 22294 525306 22350
rect 525374 22294 525430 22350
rect 525498 22294 525554 22350
rect 525622 22294 525678 22350
rect 525250 22170 525306 22226
rect 525374 22170 525430 22226
rect 525498 22170 525554 22226
rect 525622 22170 525678 22226
rect 525250 22046 525306 22102
rect 525374 22046 525430 22102
rect 525498 22046 525554 22102
rect 525622 22046 525678 22102
rect 525250 21922 525306 21978
rect 525374 21922 525430 21978
rect 525498 21922 525554 21978
rect 525622 21922 525678 21978
rect 525250 4294 525306 4350
rect 525374 4294 525430 4350
rect 525498 4294 525554 4350
rect 525622 4294 525678 4350
rect 525250 4170 525306 4226
rect 525374 4170 525430 4226
rect 525498 4170 525554 4226
rect 525622 4170 525678 4226
rect 525250 4046 525306 4102
rect 525374 4046 525430 4102
rect 525498 4046 525554 4102
rect 525622 4046 525678 4102
rect 525250 3922 525306 3978
rect 525374 3922 525430 3978
rect 525498 3922 525554 3978
rect 525622 3922 525678 3978
rect 525250 -216 525306 -160
rect 525374 -216 525430 -160
rect 525498 -216 525554 -160
rect 525622 -216 525678 -160
rect 525250 -340 525306 -284
rect 525374 -340 525430 -284
rect 525498 -340 525554 -284
rect 525622 -340 525678 -284
rect 525250 -464 525306 -408
rect 525374 -464 525430 -408
rect 525498 -464 525554 -408
rect 525622 -464 525678 -408
rect 525250 -588 525306 -532
rect 525374 -588 525430 -532
rect 525498 -588 525554 -532
rect 525622 -588 525678 -532
rect 528970 598116 529026 598172
rect 529094 598116 529150 598172
rect 529218 598116 529274 598172
rect 529342 598116 529398 598172
rect 528970 597992 529026 598048
rect 529094 597992 529150 598048
rect 529218 597992 529274 598048
rect 529342 597992 529398 598048
rect 528970 597868 529026 597924
rect 529094 597868 529150 597924
rect 529218 597868 529274 597924
rect 529342 597868 529398 597924
rect 528970 597744 529026 597800
rect 529094 597744 529150 597800
rect 529218 597744 529274 597800
rect 529342 597744 529398 597800
rect 528970 586294 529026 586350
rect 529094 586294 529150 586350
rect 529218 586294 529274 586350
rect 529342 586294 529398 586350
rect 528970 586170 529026 586226
rect 529094 586170 529150 586226
rect 529218 586170 529274 586226
rect 529342 586170 529398 586226
rect 528970 586046 529026 586102
rect 529094 586046 529150 586102
rect 529218 586046 529274 586102
rect 529342 586046 529398 586102
rect 528970 585922 529026 585978
rect 529094 585922 529150 585978
rect 529218 585922 529274 585978
rect 529342 585922 529398 585978
rect 528970 568294 529026 568350
rect 529094 568294 529150 568350
rect 529218 568294 529274 568350
rect 529342 568294 529398 568350
rect 528970 568170 529026 568226
rect 529094 568170 529150 568226
rect 529218 568170 529274 568226
rect 529342 568170 529398 568226
rect 528970 568046 529026 568102
rect 529094 568046 529150 568102
rect 529218 568046 529274 568102
rect 529342 568046 529398 568102
rect 528970 567922 529026 567978
rect 529094 567922 529150 567978
rect 529218 567922 529274 567978
rect 529342 567922 529398 567978
rect 528970 550294 529026 550350
rect 529094 550294 529150 550350
rect 529218 550294 529274 550350
rect 529342 550294 529398 550350
rect 528970 550170 529026 550226
rect 529094 550170 529150 550226
rect 529218 550170 529274 550226
rect 529342 550170 529398 550226
rect 528970 550046 529026 550102
rect 529094 550046 529150 550102
rect 529218 550046 529274 550102
rect 529342 550046 529398 550102
rect 528970 549922 529026 549978
rect 529094 549922 529150 549978
rect 529218 549922 529274 549978
rect 529342 549922 529398 549978
rect 528970 532294 529026 532350
rect 529094 532294 529150 532350
rect 529218 532294 529274 532350
rect 529342 532294 529398 532350
rect 528970 532170 529026 532226
rect 529094 532170 529150 532226
rect 529218 532170 529274 532226
rect 529342 532170 529398 532226
rect 528970 532046 529026 532102
rect 529094 532046 529150 532102
rect 529218 532046 529274 532102
rect 529342 532046 529398 532102
rect 528970 531922 529026 531978
rect 529094 531922 529150 531978
rect 529218 531922 529274 531978
rect 529342 531922 529398 531978
rect 528970 514294 529026 514350
rect 529094 514294 529150 514350
rect 529218 514294 529274 514350
rect 529342 514294 529398 514350
rect 528970 514170 529026 514226
rect 529094 514170 529150 514226
rect 529218 514170 529274 514226
rect 529342 514170 529398 514226
rect 528970 514046 529026 514102
rect 529094 514046 529150 514102
rect 529218 514046 529274 514102
rect 529342 514046 529398 514102
rect 528970 513922 529026 513978
rect 529094 513922 529150 513978
rect 529218 513922 529274 513978
rect 529342 513922 529398 513978
rect 528970 496294 529026 496350
rect 529094 496294 529150 496350
rect 529218 496294 529274 496350
rect 529342 496294 529398 496350
rect 528970 496170 529026 496226
rect 529094 496170 529150 496226
rect 529218 496170 529274 496226
rect 529342 496170 529398 496226
rect 528970 496046 529026 496102
rect 529094 496046 529150 496102
rect 529218 496046 529274 496102
rect 529342 496046 529398 496102
rect 528970 495922 529026 495978
rect 529094 495922 529150 495978
rect 529218 495922 529274 495978
rect 529342 495922 529398 495978
rect 528970 478294 529026 478350
rect 529094 478294 529150 478350
rect 529218 478294 529274 478350
rect 529342 478294 529398 478350
rect 528970 478170 529026 478226
rect 529094 478170 529150 478226
rect 529218 478170 529274 478226
rect 529342 478170 529398 478226
rect 528970 478046 529026 478102
rect 529094 478046 529150 478102
rect 529218 478046 529274 478102
rect 529342 478046 529398 478102
rect 528970 477922 529026 477978
rect 529094 477922 529150 477978
rect 529218 477922 529274 477978
rect 529342 477922 529398 477978
rect 528970 460294 529026 460350
rect 529094 460294 529150 460350
rect 529218 460294 529274 460350
rect 529342 460294 529398 460350
rect 528970 460170 529026 460226
rect 529094 460170 529150 460226
rect 529218 460170 529274 460226
rect 529342 460170 529398 460226
rect 528970 460046 529026 460102
rect 529094 460046 529150 460102
rect 529218 460046 529274 460102
rect 529342 460046 529398 460102
rect 528970 459922 529026 459978
rect 529094 459922 529150 459978
rect 529218 459922 529274 459978
rect 529342 459922 529398 459978
rect 528970 442294 529026 442350
rect 529094 442294 529150 442350
rect 529218 442294 529274 442350
rect 529342 442294 529398 442350
rect 528970 442170 529026 442226
rect 529094 442170 529150 442226
rect 529218 442170 529274 442226
rect 529342 442170 529398 442226
rect 528970 442046 529026 442102
rect 529094 442046 529150 442102
rect 529218 442046 529274 442102
rect 529342 442046 529398 442102
rect 528970 441922 529026 441978
rect 529094 441922 529150 441978
rect 529218 441922 529274 441978
rect 529342 441922 529398 441978
rect 528970 424294 529026 424350
rect 529094 424294 529150 424350
rect 529218 424294 529274 424350
rect 529342 424294 529398 424350
rect 528970 424170 529026 424226
rect 529094 424170 529150 424226
rect 529218 424170 529274 424226
rect 529342 424170 529398 424226
rect 528970 424046 529026 424102
rect 529094 424046 529150 424102
rect 529218 424046 529274 424102
rect 529342 424046 529398 424102
rect 528970 423922 529026 423978
rect 529094 423922 529150 423978
rect 529218 423922 529274 423978
rect 529342 423922 529398 423978
rect 528970 406294 529026 406350
rect 529094 406294 529150 406350
rect 529218 406294 529274 406350
rect 529342 406294 529398 406350
rect 528970 406170 529026 406226
rect 529094 406170 529150 406226
rect 529218 406170 529274 406226
rect 529342 406170 529398 406226
rect 528970 406046 529026 406102
rect 529094 406046 529150 406102
rect 529218 406046 529274 406102
rect 529342 406046 529398 406102
rect 528970 405922 529026 405978
rect 529094 405922 529150 405978
rect 529218 405922 529274 405978
rect 529342 405922 529398 405978
rect 528970 388294 529026 388350
rect 529094 388294 529150 388350
rect 529218 388294 529274 388350
rect 529342 388294 529398 388350
rect 528970 388170 529026 388226
rect 529094 388170 529150 388226
rect 529218 388170 529274 388226
rect 529342 388170 529398 388226
rect 528970 388046 529026 388102
rect 529094 388046 529150 388102
rect 529218 388046 529274 388102
rect 529342 388046 529398 388102
rect 528970 387922 529026 387978
rect 529094 387922 529150 387978
rect 529218 387922 529274 387978
rect 529342 387922 529398 387978
rect 528970 370294 529026 370350
rect 529094 370294 529150 370350
rect 529218 370294 529274 370350
rect 529342 370294 529398 370350
rect 528970 370170 529026 370226
rect 529094 370170 529150 370226
rect 529218 370170 529274 370226
rect 529342 370170 529398 370226
rect 528970 370046 529026 370102
rect 529094 370046 529150 370102
rect 529218 370046 529274 370102
rect 529342 370046 529398 370102
rect 528970 369922 529026 369978
rect 529094 369922 529150 369978
rect 529218 369922 529274 369978
rect 529342 369922 529398 369978
rect 528970 352294 529026 352350
rect 529094 352294 529150 352350
rect 529218 352294 529274 352350
rect 529342 352294 529398 352350
rect 528970 352170 529026 352226
rect 529094 352170 529150 352226
rect 529218 352170 529274 352226
rect 529342 352170 529398 352226
rect 528970 352046 529026 352102
rect 529094 352046 529150 352102
rect 529218 352046 529274 352102
rect 529342 352046 529398 352102
rect 528970 351922 529026 351978
rect 529094 351922 529150 351978
rect 529218 351922 529274 351978
rect 529342 351922 529398 351978
rect 528970 334294 529026 334350
rect 529094 334294 529150 334350
rect 529218 334294 529274 334350
rect 529342 334294 529398 334350
rect 528970 334170 529026 334226
rect 529094 334170 529150 334226
rect 529218 334170 529274 334226
rect 529342 334170 529398 334226
rect 528970 334046 529026 334102
rect 529094 334046 529150 334102
rect 529218 334046 529274 334102
rect 529342 334046 529398 334102
rect 528970 333922 529026 333978
rect 529094 333922 529150 333978
rect 529218 333922 529274 333978
rect 529342 333922 529398 333978
rect 528970 316294 529026 316350
rect 529094 316294 529150 316350
rect 529218 316294 529274 316350
rect 529342 316294 529398 316350
rect 528970 316170 529026 316226
rect 529094 316170 529150 316226
rect 529218 316170 529274 316226
rect 529342 316170 529398 316226
rect 528970 316046 529026 316102
rect 529094 316046 529150 316102
rect 529218 316046 529274 316102
rect 529342 316046 529398 316102
rect 528970 315922 529026 315978
rect 529094 315922 529150 315978
rect 529218 315922 529274 315978
rect 529342 315922 529398 315978
rect 528970 298294 529026 298350
rect 529094 298294 529150 298350
rect 529218 298294 529274 298350
rect 529342 298294 529398 298350
rect 528970 298170 529026 298226
rect 529094 298170 529150 298226
rect 529218 298170 529274 298226
rect 529342 298170 529398 298226
rect 528970 298046 529026 298102
rect 529094 298046 529150 298102
rect 529218 298046 529274 298102
rect 529342 298046 529398 298102
rect 528970 297922 529026 297978
rect 529094 297922 529150 297978
rect 529218 297922 529274 297978
rect 529342 297922 529398 297978
rect 528970 280294 529026 280350
rect 529094 280294 529150 280350
rect 529218 280294 529274 280350
rect 529342 280294 529398 280350
rect 528970 280170 529026 280226
rect 529094 280170 529150 280226
rect 529218 280170 529274 280226
rect 529342 280170 529398 280226
rect 528970 280046 529026 280102
rect 529094 280046 529150 280102
rect 529218 280046 529274 280102
rect 529342 280046 529398 280102
rect 528970 279922 529026 279978
rect 529094 279922 529150 279978
rect 529218 279922 529274 279978
rect 529342 279922 529398 279978
rect 528970 262294 529026 262350
rect 529094 262294 529150 262350
rect 529218 262294 529274 262350
rect 529342 262294 529398 262350
rect 528970 262170 529026 262226
rect 529094 262170 529150 262226
rect 529218 262170 529274 262226
rect 529342 262170 529398 262226
rect 528970 262046 529026 262102
rect 529094 262046 529150 262102
rect 529218 262046 529274 262102
rect 529342 262046 529398 262102
rect 528970 261922 529026 261978
rect 529094 261922 529150 261978
rect 529218 261922 529274 261978
rect 529342 261922 529398 261978
rect 528970 244294 529026 244350
rect 529094 244294 529150 244350
rect 529218 244294 529274 244350
rect 529342 244294 529398 244350
rect 528970 244170 529026 244226
rect 529094 244170 529150 244226
rect 529218 244170 529274 244226
rect 529342 244170 529398 244226
rect 528970 244046 529026 244102
rect 529094 244046 529150 244102
rect 529218 244046 529274 244102
rect 529342 244046 529398 244102
rect 528970 243922 529026 243978
rect 529094 243922 529150 243978
rect 529218 243922 529274 243978
rect 529342 243922 529398 243978
rect 528970 226294 529026 226350
rect 529094 226294 529150 226350
rect 529218 226294 529274 226350
rect 529342 226294 529398 226350
rect 528970 226170 529026 226226
rect 529094 226170 529150 226226
rect 529218 226170 529274 226226
rect 529342 226170 529398 226226
rect 528970 226046 529026 226102
rect 529094 226046 529150 226102
rect 529218 226046 529274 226102
rect 529342 226046 529398 226102
rect 528970 225922 529026 225978
rect 529094 225922 529150 225978
rect 529218 225922 529274 225978
rect 529342 225922 529398 225978
rect 528970 208294 529026 208350
rect 529094 208294 529150 208350
rect 529218 208294 529274 208350
rect 529342 208294 529398 208350
rect 528970 208170 529026 208226
rect 529094 208170 529150 208226
rect 529218 208170 529274 208226
rect 529342 208170 529398 208226
rect 528970 208046 529026 208102
rect 529094 208046 529150 208102
rect 529218 208046 529274 208102
rect 529342 208046 529398 208102
rect 528970 207922 529026 207978
rect 529094 207922 529150 207978
rect 529218 207922 529274 207978
rect 529342 207922 529398 207978
rect 528970 190294 529026 190350
rect 529094 190294 529150 190350
rect 529218 190294 529274 190350
rect 529342 190294 529398 190350
rect 528970 190170 529026 190226
rect 529094 190170 529150 190226
rect 529218 190170 529274 190226
rect 529342 190170 529398 190226
rect 528970 190046 529026 190102
rect 529094 190046 529150 190102
rect 529218 190046 529274 190102
rect 529342 190046 529398 190102
rect 528970 189922 529026 189978
rect 529094 189922 529150 189978
rect 529218 189922 529274 189978
rect 529342 189922 529398 189978
rect 528970 172294 529026 172350
rect 529094 172294 529150 172350
rect 529218 172294 529274 172350
rect 529342 172294 529398 172350
rect 528970 172170 529026 172226
rect 529094 172170 529150 172226
rect 529218 172170 529274 172226
rect 529342 172170 529398 172226
rect 528970 172046 529026 172102
rect 529094 172046 529150 172102
rect 529218 172046 529274 172102
rect 529342 172046 529398 172102
rect 528970 171922 529026 171978
rect 529094 171922 529150 171978
rect 529218 171922 529274 171978
rect 529342 171922 529398 171978
rect 528970 154294 529026 154350
rect 529094 154294 529150 154350
rect 529218 154294 529274 154350
rect 529342 154294 529398 154350
rect 528970 154170 529026 154226
rect 529094 154170 529150 154226
rect 529218 154170 529274 154226
rect 529342 154170 529398 154226
rect 528970 154046 529026 154102
rect 529094 154046 529150 154102
rect 529218 154046 529274 154102
rect 529342 154046 529398 154102
rect 528970 153922 529026 153978
rect 529094 153922 529150 153978
rect 529218 153922 529274 153978
rect 529342 153922 529398 153978
rect 528970 136294 529026 136350
rect 529094 136294 529150 136350
rect 529218 136294 529274 136350
rect 529342 136294 529398 136350
rect 528970 136170 529026 136226
rect 529094 136170 529150 136226
rect 529218 136170 529274 136226
rect 529342 136170 529398 136226
rect 528970 136046 529026 136102
rect 529094 136046 529150 136102
rect 529218 136046 529274 136102
rect 529342 136046 529398 136102
rect 528970 135922 529026 135978
rect 529094 135922 529150 135978
rect 529218 135922 529274 135978
rect 529342 135922 529398 135978
rect 528970 118294 529026 118350
rect 529094 118294 529150 118350
rect 529218 118294 529274 118350
rect 529342 118294 529398 118350
rect 528970 118170 529026 118226
rect 529094 118170 529150 118226
rect 529218 118170 529274 118226
rect 529342 118170 529398 118226
rect 528970 118046 529026 118102
rect 529094 118046 529150 118102
rect 529218 118046 529274 118102
rect 529342 118046 529398 118102
rect 528970 117922 529026 117978
rect 529094 117922 529150 117978
rect 529218 117922 529274 117978
rect 529342 117922 529398 117978
rect 528970 100294 529026 100350
rect 529094 100294 529150 100350
rect 529218 100294 529274 100350
rect 529342 100294 529398 100350
rect 528970 100170 529026 100226
rect 529094 100170 529150 100226
rect 529218 100170 529274 100226
rect 529342 100170 529398 100226
rect 528970 100046 529026 100102
rect 529094 100046 529150 100102
rect 529218 100046 529274 100102
rect 529342 100046 529398 100102
rect 528970 99922 529026 99978
rect 529094 99922 529150 99978
rect 529218 99922 529274 99978
rect 529342 99922 529398 99978
rect 528970 82294 529026 82350
rect 529094 82294 529150 82350
rect 529218 82294 529274 82350
rect 529342 82294 529398 82350
rect 528970 82170 529026 82226
rect 529094 82170 529150 82226
rect 529218 82170 529274 82226
rect 529342 82170 529398 82226
rect 528970 82046 529026 82102
rect 529094 82046 529150 82102
rect 529218 82046 529274 82102
rect 529342 82046 529398 82102
rect 528970 81922 529026 81978
rect 529094 81922 529150 81978
rect 529218 81922 529274 81978
rect 529342 81922 529398 81978
rect 528970 64294 529026 64350
rect 529094 64294 529150 64350
rect 529218 64294 529274 64350
rect 529342 64294 529398 64350
rect 528970 64170 529026 64226
rect 529094 64170 529150 64226
rect 529218 64170 529274 64226
rect 529342 64170 529398 64226
rect 528970 64046 529026 64102
rect 529094 64046 529150 64102
rect 529218 64046 529274 64102
rect 529342 64046 529398 64102
rect 528970 63922 529026 63978
rect 529094 63922 529150 63978
rect 529218 63922 529274 63978
rect 529342 63922 529398 63978
rect 528970 46294 529026 46350
rect 529094 46294 529150 46350
rect 529218 46294 529274 46350
rect 529342 46294 529398 46350
rect 528970 46170 529026 46226
rect 529094 46170 529150 46226
rect 529218 46170 529274 46226
rect 529342 46170 529398 46226
rect 528970 46046 529026 46102
rect 529094 46046 529150 46102
rect 529218 46046 529274 46102
rect 529342 46046 529398 46102
rect 528970 45922 529026 45978
rect 529094 45922 529150 45978
rect 529218 45922 529274 45978
rect 529342 45922 529398 45978
rect 528970 28294 529026 28350
rect 529094 28294 529150 28350
rect 529218 28294 529274 28350
rect 529342 28294 529398 28350
rect 528970 28170 529026 28226
rect 529094 28170 529150 28226
rect 529218 28170 529274 28226
rect 529342 28170 529398 28226
rect 528970 28046 529026 28102
rect 529094 28046 529150 28102
rect 529218 28046 529274 28102
rect 529342 28046 529398 28102
rect 528970 27922 529026 27978
rect 529094 27922 529150 27978
rect 529218 27922 529274 27978
rect 529342 27922 529398 27978
rect 528970 10294 529026 10350
rect 529094 10294 529150 10350
rect 529218 10294 529274 10350
rect 529342 10294 529398 10350
rect 528970 10170 529026 10226
rect 529094 10170 529150 10226
rect 529218 10170 529274 10226
rect 529342 10170 529398 10226
rect 528970 10046 529026 10102
rect 529094 10046 529150 10102
rect 529218 10046 529274 10102
rect 529342 10046 529398 10102
rect 528970 9922 529026 9978
rect 529094 9922 529150 9978
rect 529218 9922 529274 9978
rect 529342 9922 529398 9978
rect 528970 -1176 529026 -1120
rect 529094 -1176 529150 -1120
rect 529218 -1176 529274 -1120
rect 529342 -1176 529398 -1120
rect 528970 -1300 529026 -1244
rect 529094 -1300 529150 -1244
rect 529218 -1300 529274 -1244
rect 529342 -1300 529398 -1244
rect 528970 -1424 529026 -1368
rect 529094 -1424 529150 -1368
rect 529218 -1424 529274 -1368
rect 529342 -1424 529398 -1368
rect 528970 -1548 529026 -1492
rect 529094 -1548 529150 -1492
rect 529218 -1548 529274 -1492
rect 529342 -1548 529398 -1492
rect 543250 597156 543306 597212
rect 543374 597156 543430 597212
rect 543498 597156 543554 597212
rect 543622 597156 543678 597212
rect 543250 597032 543306 597088
rect 543374 597032 543430 597088
rect 543498 597032 543554 597088
rect 543622 597032 543678 597088
rect 543250 596908 543306 596964
rect 543374 596908 543430 596964
rect 543498 596908 543554 596964
rect 543622 596908 543678 596964
rect 543250 596784 543306 596840
rect 543374 596784 543430 596840
rect 543498 596784 543554 596840
rect 543622 596784 543678 596840
rect 543250 580294 543306 580350
rect 543374 580294 543430 580350
rect 543498 580294 543554 580350
rect 543622 580294 543678 580350
rect 543250 580170 543306 580226
rect 543374 580170 543430 580226
rect 543498 580170 543554 580226
rect 543622 580170 543678 580226
rect 543250 580046 543306 580102
rect 543374 580046 543430 580102
rect 543498 580046 543554 580102
rect 543622 580046 543678 580102
rect 543250 579922 543306 579978
rect 543374 579922 543430 579978
rect 543498 579922 543554 579978
rect 543622 579922 543678 579978
rect 543250 562294 543306 562350
rect 543374 562294 543430 562350
rect 543498 562294 543554 562350
rect 543622 562294 543678 562350
rect 543250 562170 543306 562226
rect 543374 562170 543430 562226
rect 543498 562170 543554 562226
rect 543622 562170 543678 562226
rect 543250 562046 543306 562102
rect 543374 562046 543430 562102
rect 543498 562046 543554 562102
rect 543622 562046 543678 562102
rect 543250 561922 543306 561978
rect 543374 561922 543430 561978
rect 543498 561922 543554 561978
rect 543622 561922 543678 561978
rect 543250 544294 543306 544350
rect 543374 544294 543430 544350
rect 543498 544294 543554 544350
rect 543622 544294 543678 544350
rect 543250 544170 543306 544226
rect 543374 544170 543430 544226
rect 543498 544170 543554 544226
rect 543622 544170 543678 544226
rect 543250 544046 543306 544102
rect 543374 544046 543430 544102
rect 543498 544046 543554 544102
rect 543622 544046 543678 544102
rect 543250 543922 543306 543978
rect 543374 543922 543430 543978
rect 543498 543922 543554 543978
rect 543622 543922 543678 543978
rect 543250 526294 543306 526350
rect 543374 526294 543430 526350
rect 543498 526294 543554 526350
rect 543622 526294 543678 526350
rect 543250 526170 543306 526226
rect 543374 526170 543430 526226
rect 543498 526170 543554 526226
rect 543622 526170 543678 526226
rect 543250 526046 543306 526102
rect 543374 526046 543430 526102
rect 543498 526046 543554 526102
rect 543622 526046 543678 526102
rect 543250 525922 543306 525978
rect 543374 525922 543430 525978
rect 543498 525922 543554 525978
rect 543622 525922 543678 525978
rect 543250 508294 543306 508350
rect 543374 508294 543430 508350
rect 543498 508294 543554 508350
rect 543622 508294 543678 508350
rect 543250 508170 543306 508226
rect 543374 508170 543430 508226
rect 543498 508170 543554 508226
rect 543622 508170 543678 508226
rect 543250 508046 543306 508102
rect 543374 508046 543430 508102
rect 543498 508046 543554 508102
rect 543622 508046 543678 508102
rect 543250 507922 543306 507978
rect 543374 507922 543430 507978
rect 543498 507922 543554 507978
rect 543622 507922 543678 507978
rect 543250 490294 543306 490350
rect 543374 490294 543430 490350
rect 543498 490294 543554 490350
rect 543622 490294 543678 490350
rect 543250 490170 543306 490226
rect 543374 490170 543430 490226
rect 543498 490170 543554 490226
rect 543622 490170 543678 490226
rect 543250 490046 543306 490102
rect 543374 490046 543430 490102
rect 543498 490046 543554 490102
rect 543622 490046 543678 490102
rect 543250 489922 543306 489978
rect 543374 489922 543430 489978
rect 543498 489922 543554 489978
rect 543622 489922 543678 489978
rect 543250 472294 543306 472350
rect 543374 472294 543430 472350
rect 543498 472294 543554 472350
rect 543622 472294 543678 472350
rect 543250 472170 543306 472226
rect 543374 472170 543430 472226
rect 543498 472170 543554 472226
rect 543622 472170 543678 472226
rect 543250 472046 543306 472102
rect 543374 472046 543430 472102
rect 543498 472046 543554 472102
rect 543622 472046 543678 472102
rect 543250 471922 543306 471978
rect 543374 471922 543430 471978
rect 543498 471922 543554 471978
rect 543622 471922 543678 471978
rect 543250 454294 543306 454350
rect 543374 454294 543430 454350
rect 543498 454294 543554 454350
rect 543622 454294 543678 454350
rect 543250 454170 543306 454226
rect 543374 454170 543430 454226
rect 543498 454170 543554 454226
rect 543622 454170 543678 454226
rect 543250 454046 543306 454102
rect 543374 454046 543430 454102
rect 543498 454046 543554 454102
rect 543622 454046 543678 454102
rect 543250 453922 543306 453978
rect 543374 453922 543430 453978
rect 543498 453922 543554 453978
rect 543622 453922 543678 453978
rect 543250 436294 543306 436350
rect 543374 436294 543430 436350
rect 543498 436294 543554 436350
rect 543622 436294 543678 436350
rect 543250 436170 543306 436226
rect 543374 436170 543430 436226
rect 543498 436170 543554 436226
rect 543622 436170 543678 436226
rect 543250 436046 543306 436102
rect 543374 436046 543430 436102
rect 543498 436046 543554 436102
rect 543622 436046 543678 436102
rect 543250 435922 543306 435978
rect 543374 435922 543430 435978
rect 543498 435922 543554 435978
rect 543622 435922 543678 435978
rect 543250 418294 543306 418350
rect 543374 418294 543430 418350
rect 543498 418294 543554 418350
rect 543622 418294 543678 418350
rect 543250 418170 543306 418226
rect 543374 418170 543430 418226
rect 543498 418170 543554 418226
rect 543622 418170 543678 418226
rect 543250 418046 543306 418102
rect 543374 418046 543430 418102
rect 543498 418046 543554 418102
rect 543622 418046 543678 418102
rect 543250 417922 543306 417978
rect 543374 417922 543430 417978
rect 543498 417922 543554 417978
rect 543622 417922 543678 417978
rect 543250 400294 543306 400350
rect 543374 400294 543430 400350
rect 543498 400294 543554 400350
rect 543622 400294 543678 400350
rect 543250 400170 543306 400226
rect 543374 400170 543430 400226
rect 543498 400170 543554 400226
rect 543622 400170 543678 400226
rect 543250 400046 543306 400102
rect 543374 400046 543430 400102
rect 543498 400046 543554 400102
rect 543622 400046 543678 400102
rect 543250 399922 543306 399978
rect 543374 399922 543430 399978
rect 543498 399922 543554 399978
rect 543622 399922 543678 399978
rect 543250 382294 543306 382350
rect 543374 382294 543430 382350
rect 543498 382294 543554 382350
rect 543622 382294 543678 382350
rect 543250 382170 543306 382226
rect 543374 382170 543430 382226
rect 543498 382170 543554 382226
rect 543622 382170 543678 382226
rect 543250 382046 543306 382102
rect 543374 382046 543430 382102
rect 543498 382046 543554 382102
rect 543622 382046 543678 382102
rect 543250 381922 543306 381978
rect 543374 381922 543430 381978
rect 543498 381922 543554 381978
rect 543622 381922 543678 381978
rect 543250 364294 543306 364350
rect 543374 364294 543430 364350
rect 543498 364294 543554 364350
rect 543622 364294 543678 364350
rect 543250 364170 543306 364226
rect 543374 364170 543430 364226
rect 543498 364170 543554 364226
rect 543622 364170 543678 364226
rect 543250 364046 543306 364102
rect 543374 364046 543430 364102
rect 543498 364046 543554 364102
rect 543622 364046 543678 364102
rect 543250 363922 543306 363978
rect 543374 363922 543430 363978
rect 543498 363922 543554 363978
rect 543622 363922 543678 363978
rect 543250 346294 543306 346350
rect 543374 346294 543430 346350
rect 543498 346294 543554 346350
rect 543622 346294 543678 346350
rect 543250 346170 543306 346226
rect 543374 346170 543430 346226
rect 543498 346170 543554 346226
rect 543622 346170 543678 346226
rect 543250 346046 543306 346102
rect 543374 346046 543430 346102
rect 543498 346046 543554 346102
rect 543622 346046 543678 346102
rect 543250 345922 543306 345978
rect 543374 345922 543430 345978
rect 543498 345922 543554 345978
rect 543622 345922 543678 345978
rect 543250 328294 543306 328350
rect 543374 328294 543430 328350
rect 543498 328294 543554 328350
rect 543622 328294 543678 328350
rect 543250 328170 543306 328226
rect 543374 328170 543430 328226
rect 543498 328170 543554 328226
rect 543622 328170 543678 328226
rect 543250 328046 543306 328102
rect 543374 328046 543430 328102
rect 543498 328046 543554 328102
rect 543622 328046 543678 328102
rect 543250 327922 543306 327978
rect 543374 327922 543430 327978
rect 543498 327922 543554 327978
rect 543622 327922 543678 327978
rect 543250 310294 543306 310350
rect 543374 310294 543430 310350
rect 543498 310294 543554 310350
rect 543622 310294 543678 310350
rect 543250 310170 543306 310226
rect 543374 310170 543430 310226
rect 543498 310170 543554 310226
rect 543622 310170 543678 310226
rect 543250 310046 543306 310102
rect 543374 310046 543430 310102
rect 543498 310046 543554 310102
rect 543622 310046 543678 310102
rect 543250 309922 543306 309978
rect 543374 309922 543430 309978
rect 543498 309922 543554 309978
rect 543622 309922 543678 309978
rect 543250 292294 543306 292350
rect 543374 292294 543430 292350
rect 543498 292294 543554 292350
rect 543622 292294 543678 292350
rect 543250 292170 543306 292226
rect 543374 292170 543430 292226
rect 543498 292170 543554 292226
rect 543622 292170 543678 292226
rect 543250 292046 543306 292102
rect 543374 292046 543430 292102
rect 543498 292046 543554 292102
rect 543622 292046 543678 292102
rect 543250 291922 543306 291978
rect 543374 291922 543430 291978
rect 543498 291922 543554 291978
rect 543622 291922 543678 291978
rect 543250 274294 543306 274350
rect 543374 274294 543430 274350
rect 543498 274294 543554 274350
rect 543622 274294 543678 274350
rect 543250 274170 543306 274226
rect 543374 274170 543430 274226
rect 543498 274170 543554 274226
rect 543622 274170 543678 274226
rect 543250 274046 543306 274102
rect 543374 274046 543430 274102
rect 543498 274046 543554 274102
rect 543622 274046 543678 274102
rect 543250 273922 543306 273978
rect 543374 273922 543430 273978
rect 543498 273922 543554 273978
rect 543622 273922 543678 273978
rect 543250 256294 543306 256350
rect 543374 256294 543430 256350
rect 543498 256294 543554 256350
rect 543622 256294 543678 256350
rect 543250 256170 543306 256226
rect 543374 256170 543430 256226
rect 543498 256170 543554 256226
rect 543622 256170 543678 256226
rect 543250 256046 543306 256102
rect 543374 256046 543430 256102
rect 543498 256046 543554 256102
rect 543622 256046 543678 256102
rect 543250 255922 543306 255978
rect 543374 255922 543430 255978
rect 543498 255922 543554 255978
rect 543622 255922 543678 255978
rect 543250 238294 543306 238350
rect 543374 238294 543430 238350
rect 543498 238294 543554 238350
rect 543622 238294 543678 238350
rect 543250 238170 543306 238226
rect 543374 238170 543430 238226
rect 543498 238170 543554 238226
rect 543622 238170 543678 238226
rect 543250 238046 543306 238102
rect 543374 238046 543430 238102
rect 543498 238046 543554 238102
rect 543622 238046 543678 238102
rect 543250 237922 543306 237978
rect 543374 237922 543430 237978
rect 543498 237922 543554 237978
rect 543622 237922 543678 237978
rect 543250 220294 543306 220350
rect 543374 220294 543430 220350
rect 543498 220294 543554 220350
rect 543622 220294 543678 220350
rect 543250 220170 543306 220226
rect 543374 220170 543430 220226
rect 543498 220170 543554 220226
rect 543622 220170 543678 220226
rect 543250 220046 543306 220102
rect 543374 220046 543430 220102
rect 543498 220046 543554 220102
rect 543622 220046 543678 220102
rect 543250 219922 543306 219978
rect 543374 219922 543430 219978
rect 543498 219922 543554 219978
rect 543622 219922 543678 219978
rect 543250 202294 543306 202350
rect 543374 202294 543430 202350
rect 543498 202294 543554 202350
rect 543622 202294 543678 202350
rect 543250 202170 543306 202226
rect 543374 202170 543430 202226
rect 543498 202170 543554 202226
rect 543622 202170 543678 202226
rect 543250 202046 543306 202102
rect 543374 202046 543430 202102
rect 543498 202046 543554 202102
rect 543622 202046 543678 202102
rect 543250 201922 543306 201978
rect 543374 201922 543430 201978
rect 543498 201922 543554 201978
rect 543622 201922 543678 201978
rect 543250 184294 543306 184350
rect 543374 184294 543430 184350
rect 543498 184294 543554 184350
rect 543622 184294 543678 184350
rect 543250 184170 543306 184226
rect 543374 184170 543430 184226
rect 543498 184170 543554 184226
rect 543622 184170 543678 184226
rect 543250 184046 543306 184102
rect 543374 184046 543430 184102
rect 543498 184046 543554 184102
rect 543622 184046 543678 184102
rect 543250 183922 543306 183978
rect 543374 183922 543430 183978
rect 543498 183922 543554 183978
rect 543622 183922 543678 183978
rect 543250 166294 543306 166350
rect 543374 166294 543430 166350
rect 543498 166294 543554 166350
rect 543622 166294 543678 166350
rect 543250 166170 543306 166226
rect 543374 166170 543430 166226
rect 543498 166170 543554 166226
rect 543622 166170 543678 166226
rect 543250 166046 543306 166102
rect 543374 166046 543430 166102
rect 543498 166046 543554 166102
rect 543622 166046 543678 166102
rect 543250 165922 543306 165978
rect 543374 165922 543430 165978
rect 543498 165922 543554 165978
rect 543622 165922 543678 165978
rect 543250 148294 543306 148350
rect 543374 148294 543430 148350
rect 543498 148294 543554 148350
rect 543622 148294 543678 148350
rect 543250 148170 543306 148226
rect 543374 148170 543430 148226
rect 543498 148170 543554 148226
rect 543622 148170 543678 148226
rect 543250 148046 543306 148102
rect 543374 148046 543430 148102
rect 543498 148046 543554 148102
rect 543622 148046 543678 148102
rect 543250 147922 543306 147978
rect 543374 147922 543430 147978
rect 543498 147922 543554 147978
rect 543622 147922 543678 147978
rect 543250 130294 543306 130350
rect 543374 130294 543430 130350
rect 543498 130294 543554 130350
rect 543622 130294 543678 130350
rect 543250 130170 543306 130226
rect 543374 130170 543430 130226
rect 543498 130170 543554 130226
rect 543622 130170 543678 130226
rect 543250 130046 543306 130102
rect 543374 130046 543430 130102
rect 543498 130046 543554 130102
rect 543622 130046 543678 130102
rect 543250 129922 543306 129978
rect 543374 129922 543430 129978
rect 543498 129922 543554 129978
rect 543622 129922 543678 129978
rect 543250 112294 543306 112350
rect 543374 112294 543430 112350
rect 543498 112294 543554 112350
rect 543622 112294 543678 112350
rect 543250 112170 543306 112226
rect 543374 112170 543430 112226
rect 543498 112170 543554 112226
rect 543622 112170 543678 112226
rect 543250 112046 543306 112102
rect 543374 112046 543430 112102
rect 543498 112046 543554 112102
rect 543622 112046 543678 112102
rect 543250 111922 543306 111978
rect 543374 111922 543430 111978
rect 543498 111922 543554 111978
rect 543622 111922 543678 111978
rect 543250 94294 543306 94350
rect 543374 94294 543430 94350
rect 543498 94294 543554 94350
rect 543622 94294 543678 94350
rect 543250 94170 543306 94226
rect 543374 94170 543430 94226
rect 543498 94170 543554 94226
rect 543622 94170 543678 94226
rect 543250 94046 543306 94102
rect 543374 94046 543430 94102
rect 543498 94046 543554 94102
rect 543622 94046 543678 94102
rect 543250 93922 543306 93978
rect 543374 93922 543430 93978
rect 543498 93922 543554 93978
rect 543622 93922 543678 93978
rect 543250 76294 543306 76350
rect 543374 76294 543430 76350
rect 543498 76294 543554 76350
rect 543622 76294 543678 76350
rect 543250 76170 543306 76226
rect 543374 76170 543430 76226
rect 543498 76170 543554 76226
rect 543622 76170 543678 76226
rect 543250 76046 543306 76102
rect 543374 76046 543430 76102
rect 543498 76046 543554 76102
rect 543622 76046 543678 76102
rect 543250 75922 543306 75978
rect 543374 75922 543430 75978
rect 543498 75922 543554 75978
rect 543622 75922 543678 75978
rect 543250 58294 543306 58350
rect 543374 58294 543430 58350
rect 543498 58294 543554 58350
rect 543622 58294 543678 58350
rect 543250 58170 543306 58226
rect 543374 58170 543430 58226
rect 543498 58170 543554 58226
rect 543622 58170 543678 58226
rect 543250 58046 543306 58102
rect 543374 58046 543430 58102
rect 543498 58046 543554 58102
rect 543622 58046 543678 58102
rect 543250 57922 543306 57978
rect 543374 57922 543430 57978
rect 543498 57922 543554 57978
rect 543622 57922 543678 57978
rect 543250 40294 543306 40350
rect 543374 40294 543430 40350
rect 543498 40294 543554 40350
rect 543622 40294 543678 40350
rect 543250 40170 543306 40226
rect 543374 40170 543430 40226
rect 543498 40170 543554 40226
rect 543622 40170 543678 40226
rect 543250 40046 543306 40102
rect 543374 40046 543430 40102
rect 543498 40046 543554 40102
rect 543622 40046 543678 40102
rect 543250 39922 543306 39978
rect 543374 39922 543430 39978
rect 543498 39922 543554 39978
rect 543622 39922 543678 39978
rect 543250 22294 543306 22350
rect 543374 22294 543430 22350
rect 543498 22294 543554 22350
rect 543622 22294 543678 22350
rect 543250 22170 543306 22226
rect 543374 22170 543430 22226
rect 543498 22170 543554 22226
rect 543622 22170 543678 22226
rect 543250 22046 543306 22102
rect 543374 22046 543430 22102
rect 543498 22046 543554 22102
rect 543622 22046 543678 22102
rect 543250 21922 543306 21978
rect 543374 21922 543430 21978
rect 543498 21922 543554 21978
rect 543622 21922 543678 21978
rect 543250 4294 543306 4350
rect 543374 4294 543430 4350
rect 543498 4294 543554 4350
rect 543622 4294 543678 4350
rect 543250 4170 543306 4226
rect 543374 4170 543430 4226
rect 543498 4170 543554 4226
rect 543622 4170 543678 4226
rect 543250 4046 543306 4102
rect 543374 4046 543430 4102
rect 543498 4046 543554 4102
rect 543622 4046 543678 4102
rect 543250 3922 543306 3978
rect 543374 3922 543430 3978
rect 543498 3922 543554 3978
rect 543622 3922 543678 3978
rect 543250 -216 543306 -160
rect 543374 -216 543430 -160
rect 543498 -216 543554 -160
rect 543622 -216 543678 -160
rect 543250 -340 543306 -284
rect 543374 -340 543430 -284
rect 543498 -340 543554 -284
rect 543622 -340 543678 -284
rect 543250 -464 543306 -408
rect 543374 -464 543430 -408
rect 543498 -464 543554 -408
rect 543622 -464 543678 -408
rect 543250 -588 543306 -532
rect 543374 -588 543430 -532
rect 543498 -588 543554 -532
rect 543622 -588 543678 -532
rect 546970 598116 547026 598172
rect 547094 598116 547150 598172
rect 547218 598116 547274 598172
rect 547342 598116 547398 598172
rect 546970 597992 547026 598048
rect 547094 597992 547150 598048
rect 547218 597992 547274 598048
rect 547342 597992 547398 598048
rect 546970 597868 547026 597924
rect 547094 597868 547150 597924
rect 547218 597868 547274 597924
rect 547342 597868 547398 597924
rect 546970 597744 547026 597800
rect 547094 597744 547150 597800
rect 547218 597744 547274 597800
rect 547342 597744 547398 597800
rect 546970 586294 547026 586350
rect 547094 586294 547150 586350
rect 547218 586294 547274 586350
rect 547342 586294 547398 586350
rect 546970 586170 547026 586226
rect 547094 586170 547150 586226
rect 547218 586170 547274 586226
rect 547342 586170 547398 586226
rect 546970 586046 547026 586102
rect 547094 586046 547150 586102
rect 547218 586046 547274 586102
rect 547342 586046 547398 586102
rect 546970 585922 547026 585978
rect 547094 585922 547150 585978
rect 547218 585922 547274 585978
rect 547342 585922 547398 585978
rect 546970 568294 547026 568350
rect 547094 568294 547150 568350
rect 547218 568294 547274 568350
rect 547342 568294 547398 568350
rect 546970 568170 547026 568226
rect 547094 568170 547150 568226
rect 547218 568170 547274 568226
rect 547342 568170 547398 568226
rect 546970 568046 547026 568102
rect 547094 568046 547150 568102
rect 547218 568046 547274 568102
rect 547342 568046 547398 568102
rect 546970 567922 547026 567978
rect 547094 567922 547150 567978
rect 547218 567922 547274 567978
rect 547342 567922 547398 567978
rect 546970 550294 547026 550350
rect 547094 550294 547150 550350
rect 547218 550294 547274 550350
rect 547342 550294 547398 550350
rect 546970 550170 547026 550226
rect 547094 550170 547150 550226
rect 547218 550170 547274 550226
rect 547342 550170 547398 550226
rect 546970 550046 547026 550102
rect 547094 550046 547150 550102
rect 547218 550046 547274 550102
rect 547342 550046 547398 550102
rect 546970 549922 547026 549978
rect 547094 549922 547150 549978
rect 547218 549922 547274 549978
rect 547342 549922 547398 549978
rect 546970 532294 547026 532350
rect 547094 532294 547150 532350
rect 547218 532294 547274 532350
rect 547342 532294 547398 532350
rect 546970 532170 547026 532226
rect 547094 532170 547150 532226
rect 547218 532170 547274 532226
rect 547342 532170 547398 532226
rect 546970 532046 547026 532102
rect 547094 532046 547150 532102
rect 547218 532046 547274 532102
rect 547342 532046 547398 532102
rect 546970 531922 547026 531978
rect 547094 531922 547150 531978
rect 547218 531922 547274 531978
rect 547342 531922 547398 531978
rect 546970 514294 547026 514350
rect 547094 514294 547150 514350
rect 547218 514294 547274 514350
rect 547342 514294 547398 514350
rect 546970 514170 547026 514226
rect 547094 514170 547150 514226
rect 547218 514170 547274 514226
rect 547342 514170 547398 514226
rect 546970 514046 547026 514102
rect 547094 514046 547150 514102
rect 547218 514046 547274 514102
rect 547342 514046 547398 514102
rect 546970 513922 547026 513978
rect 547094 513922 547150 513978
rect 547218 513922 547274 513978
rect 547342 513922 547398 513978
rect 546970 496294 547026 496350
rect 547094 496294 547150 496350
rect 547218 496294 547274 496350
rect 547342 496294 547398 496350
rect 546970 496170 547026 496226
rect 547094 496170 547150 496226
rect 547218 496170 547274 496226
rect 547342 496170 547398 496226
rect 546970 496046 547026 496102
rect 547094 496046 547150 496102
rect 547218 496046 547274 496102
rect 547342 496046 547398 496102
rect 546970 495922 547026 495978
rect 547094 495922 547150 495978
rect 547218 495922 547274 495978
rect 547342 495922 547398 495978
rect 546970 478294 547026 478350
rect 547094 478294 547150 478350
rect 547218 478294 547274 478350
rect 547342 478294 547398 478350
rect 546970 478170 547026 478226
rect 547094 478170 547150 478226
rect 547218 478170 547274 478226
rect 547342 478170 547398 478226
rect 546970 478046 547026 478102
rect 547094 478046 547150 478102
rect 547218 478046 547274 478102
rect 547342 478046 547398 478102
rect 546970 477922 547026 477978
rect 547094 477922 547150 477978
rect 547218 477922 547274 477978
rect 547342 477922 547398 477978
rect 546970 460294 547026 460350
rect 547094 460294 547150 460350
rect 547218 460294 547274 460350
rect 547342 460294 547398 460350
rect 546970 460170 547026 460226
rect 547094 460170 547150 460226
rect 547218 460170 547274 460226
rect 547342 460170 547398 460226
rect 546970 460046 547026 460102
rect 547094 460046 547150 460102
rect 547218 460046 547274 460102
rect 547342 460046 547398 460102
rect 546970 459922 547026 459978
rect 547094 459922 547150 459978
rect 547218 459922 547274 459978
rect 547342 459922 547398 459978
rect 546970 442294 547026 442350
rect 547094 442294 547150 442350
rect 547218 442294 547274 442350
rect 547342 442294 547398 442350
rect 546970 442170 547026 442226
rect 547094 442170 547150 442226
rect 547218 442170 547274 442226
rect 547342 442170 547398 442226
rect 546970 442046 547026 442102
rect 547094 442046 547150 442102
rect 547218 442046 547274 442102
rect 547342 442046 547398 442102
rect 546970 441922 547026 441978
rect 547094 441922 547150 441978
rect 547218 441922 547274 441978
rect 547342 441922 547398 441978
rect 546970 424294 547026 424350
rect 547094 424294 547150 424350
rect 547218 424294 547274 424350
rect 547342 424294 547398 424350
rect 546970 424170 547026 424226
rect 547094 424170 547150 424226
rect 547218 424170 547274 424226
rect 547342 424170 547398 424226
rect 546970 424046 547026 424102
rect 547094 424046 547150 424102
rect 547218 424046 547274 424102
rect 547342 424046 547398 424102
rect 546970 423922 547026 423978
rect 547094 423922 547150 423978
rect 547218 423922 547274 423978
rect 547342 423922 547398 423978
rect 546970 406294 547026 406350
rect 547094 406294 547150 406350
rect 547218 406294 547274 406350
rect 547342 406294 547398 406350
rect 546970 406170 547026 406226
rect 547094 406170 547150 406226
rect 547218 406170 547274 406226
rect 547342 406170 547398 406226
rect 546970 406046 547026 406102
rect 547094 406046 547150 406102
rect 547218 406046 547274 406102
rect 547342 406046 547398 406102
rect 546970 405922 547026 405978
rect 547094 405922 547150 405978
rect 547218 405922 547274 405978
rect 547342 405922 547398 405978
rect 546970 388294 547026 388350
rect 547094 388294 547150 388350
rect 547218 388294 547274 388350
rect 547342 388294 547398 388350
rect 546970 388170 547026 388226
rect 547094 388170 547150 388226
rect 547218 388170 547274 388226
rect 547342 388170 547398 388226
rect 546970 388046 547026 388102
rect 547094 388046 547150 388102
rect 547218 388046 547274 388102
rect 547342 388046 547398 388102
rect 546970 387922 547026 387978
rect 547094 387922 547150 387978
rect 547218 387922 547274 387978
rect 547342 387922 547398 387978
rect 546970 370294 547026 370350
rect 547094 370294 547150 370350
rect 547218 370294 547274 370350
rect 547342 370294 547398 370350
rect 546970 370170 547026 370226
rect 547094 370170 547150 370226
rect 547218 370170 547274 370226
rect 547342 370170 547398 370226
rect 546970 370046 547026 370102
rect 547094 370046 547150 370102
rect 547218 370046 547274 370102
rect 547342 370046 547398 370102
rect 546970 369922 547026 369978
rect 547094 369922 547150 369978
rect 547218 369922 547274 369978
rect 547342 369922 547398 369978
rect 546970 352294 547026 352350
rect 547094 352294 547150 352350
rect 547218 352294 547274 352350
rect 547342 352294 547398 352350
rect 546970 352170 547026 352226
rect 547094 352170 547150 352226
rect 547218 352170 547274 352226
rect 547342 352170 547398 352226
rect 546970 352046 547026 352102
rect 547094 352046 547150 352102
rect 547218 352046 547274 352102
rect 547342 352046 547398 352102
rect 546970 351922 547026 351978
rect 547094 351922 547150 351978
rect 547218 351922 547274 351978
rect 547342 351922 547398 351978
rect 546970 334294 547026 334350
rect 547094 334294 547150 334350
rect 547218 334294 547274 334350
rect 547342 334294 547398 334350
rect 546970 334170 547026 334226
rect 547094 334170 547150 334226
rect 547218 334170 547274 334226
rect 547342 334170 547398 334226
rect 546970 334046 547026 334102
rect 547094 334046 547150 334102
rect 547218 334046 547274 334102
rect 547342 334046 547398 334102
rect 546970 333922 547026 333978
rect 547094 333922 547150 333978
rect 547218 333922 547274 333978
rect 547342 333922 547398 333978
rect 546970 316294 547026 316350
rect 547094 316294 547150 316350
rect 547218 316294 547274 316350
rect 547342 316294 547398 316350
rect 546970 316170 547026 316226
rect 547094 316170 547150 316226
rect 547218 316170 547274 316226
rect 547342 316170 547398 316226
rect 546970 316046 547026 316102
rect 547094 316046 547150 316102
rect 547218 316046 547274 316102
rect 547342 316046 547398 316102
rect 546970 315922 547026 315978
rect 547094 315922 547150 315978
rect 547218 315922 547274 315978
rect 547342 315922 547398 315978
rect 546970 298294 547026 298350
rect 547094 298294 547150 298350
rect 547218 298294 547274 298350
rect 547342 298294 547398 298350
rect 546970 298170 547026 298226
rect 547094 298170 547150 298226
rect 547218 298170 547274 298226
rect 547342 298170 547398 298226
rect 546970 298046 547026 298102
rect 547094 298046 547150 298102
rect 547218 298046 547274 298102
rect 547342 298046 547398 298102
rect 546970 297922 547026 297978
rect 547094 297922 547150 297978
rect 547218 297922 547274 297978
rect 547342 297922 547398 297978
rect 546970 280294 547026 280350
rect 547094 280294 547150 280350
rect 547218 280294 547274 280350
rect 547342 280294 547398 280350
rect 546970 280170 547026 280226
rect 547094 280170 547150 280226
rect 547218 280170 547274 280226
rect 547342 280170 547398 280226
rect 546970 280046 547026 280102
rect 547094 280046 547150 280102
rect 547218 280046 547274 280102
rect 547342 280046 547398 280102
rect 546970 279922 547026 279978
rect 547094 279922 547150 279978
rect 547218 279922 547274 279978
rect 547342 279922 547398 279978
rect 546970 262294 547026 262350
rect 547094 262294 547150 262350
rect 547218 262294 547274 262350
rect 547342 262294 547398 262350
rect 546970 262170 547026 262226
rect 547094 262170 547150 262226
rect 547218 262170 547274 262226
rect 547342 262170 547398 262226
rect 546970 262046 547026 262102
rect 547094 262046 547150 262102
rect 547218 262046 547274 262102
rect 547342 262046 547398 262102
rect 546970 261922 547026 261978
rect 547094 261922 547150 261978
rect 547218 261922 547274 261978
rect 547342 261922 547398 261978
rect 546970 244294 547026 244350
rect 547094 244294 547150 244350
rect 547218 244294 547274 244350
rect 547342 244294 547398 244350
rect 546970 244170 547026 244226
rect 547094 244170 547150 244226
rect 547218 244170 547274 244226
rect 547342 244170 547398 244226
rect 546970 244046 547026 244102
rect 547094 244046 547150 244102
rect 547218 244046 547274 244102
rect 547342 244046 547398 244102
rect 546970 243922 547026 243978
rect 547094 243922 547150 243978
rect 547218 243922 547274 243978
rect 547342 243922 547398 243978
rect 546970 226294 547026 226350
rect 547094 226294 547150 226350
rect 547218 226294 547274 226350
rect 547342 226294 547398 226350
rect 546970 226170 547026 226226
rect 547094 226170 547150 226226
rect 547218 226170 547274 226226
rect 547342 226170 547398 226226
rect 546970 226046 547026 226102
rect 547094 226046 547150 226102
rect 547218 226046 547274 226102
rect 547342 226046 547398 226102
rect 546970 225922 547026 225978
rect 547094 225922 547150 225978
rect 547218 225922 547274 225978
rect 547342 225922 547398 225978
rect 546970 208294 547026 208350
rect 547094 208294 547150 208350
rect 547218 208294 547274 208350
rect 547342 208294 547398 208350
rect 546970 208170 547026 208226
rect 547094 208170 547150 208226
rect 547218 208170 547274 208226
rect 547342 208170 547398 208226
rect 546970 208046 547026 208102
rect 547094 208046 547150 208102
rect 547218 208046 547274 208102
rect 547342 208046 547398 208102
rect 546970 207922 547026 207978
rect 547094 207922 547150 207978
rect 547218 207922 547274 207978
rect 547342 207922 547398 207978
rect 546970 190294 547026 190350
rect 547094 190294 547150 190350
rect 547218 190294 547274 190350
rect 547342 190294 547398 190350
rect 546970 190170 547026 190226
rect 547094 190170 547150 190226
rect 547218 190170 547274 190226
rect 547342 190170 547398 190226
rect 546970 190046 547026 190102
rect 547094 190046 547150 190102
rect 547218 190046 547274 190102
rect 547342 190046 547398 190102
rect 546970 189922 547026 189978
rect 547094 189922 547150 189978
rect 547218 189922 547274 189978
rect 547342 189922 547398 189978
rect 546970 172294 547026 172350
rect 547094 172294 547150 172350
rect 547218 172294 547274 172350
rect 547342 172294 547398 172350
rect 546970 172170 547026 172226
rect 547094 172170 547150 172226
rect 547218 172170 547274 172226
rect 547342 172170 547398 172226
rect 546970 172046 547026 172102
rect 547094 172046 547150 172102
rect 547218 172046 547274 172102
rect 547342 172046 547398 172102
rect 546970 171922 547026 171978
rect 547094 171922 547150 171978
rect 547218 171922 547274 171978
rect 547342 171922 547398 171978
rect 546970 154294 547026 154350
rect 547094 154294 547150 154350
rect 547218 154294 547274 154350
rect 547342 154294 547398 154350
rect 546970 154170 547026 154226
rect 547094 154170 547150 154226
rect 547218 154170 547274 154226
rect 547342 154170 547398 154226
rect 546970 154046 547026 154102
rect 547094 154046 547150 154102
rect 547218 154046 547274 154102
rect 547342 154046 547398 154102
rect 546970 153922 547026 153978
rect 547094 153922 547150 153978
rect 547218 153922 547274 153978
rect 547342 153922 547398 153978
rect 546970 136294 547026 136350
rect 547094 136294 547150 136350
rect 547218 136294 547274 136350
rect 547342 136294 547398 136350
rect 546970 136170 547026 136226
rect 547094 136170 547150 136226
rect 547218 136170 547274 136226
rect 547342 136170 547398 136226
rect 546970 136046 547026 136102
rect 547094 136046 547150 136102
rect 547218 136046 547274 136102
rect 547342 136046 547398 136102
rect 546970 135922 547026 135978
rect 547094 135922 547150 135978
rect 547218 135922 547274 135978
rect 547342 135922 547398 135978
rect 546970 118294 547026 118350
rect 547094 118294 547150 118350
rect 547218 118294 547274 118350
rect 547342 118294 547398 118350
rect 546970 118170 547026 118226
rect 547094 118170 547150 118226
rect 547218 118170 547274 118226
rect 547342 118170 547398 118226
rect 546970 118046 547026 118102
rect 547094 118046 547150 118102
rect 547218 118046 547274 118102
rect 547342 118046 547398 118102
rect 546970 117922 547026 117978
rect 547094 117922 547150 117978
rect 547218 117922 547274 117978
rect 547342 117922 547398 117978
rect 546970 100294 547026 100350
rect 547094 100294 547150 100350
rect 547218 100294 547274 100350
rect 547342 100294 547398 100350
rect 546970 100170 547026 100226
rect 547094 100170 547150 100226
rect 547218 100170 547274 100226
rect 547342 100170 547398 100226
rect 546970 100046 547026 100102
rect 547094 100046 547150 100102
rect 547218 100046 547274 100102
rect 547342 100046 547398 100102
rect 546970 99922 547026 99978
rect 547094 99922 547150 99978
rect 547218 99922 547274 99978
rect 547342 99922 547398 99978
rect 546970 82294 547026 82350
rect 547094 82294 547150 82350
rect 547218 82294 547274 82350
rect 547342 82294 547398 82350
rect 546970 82170 547026 82226
rect 547094 82170 547150 82226
rect 547218 82170 547274 82226
rect 547342 82170 547398 82226
rect 546970 82046 547026 82102
rect 547094 82046 547150 82102
rect 547218 82046 547274 82102
rect 547342 82046 547398 82102
rect 546970 81922 547026 81978
rect 547094 81922 547150 81978
rect 547218 81922 547274 81978
rect 547342 81922 547398 81978
rect 546970 64294 547026 64350
rect 547094 64294 547150 64350
rect 547218 64294 547274 64350
rect 547342 64294 547398 64350
rect 546970 64170 547026 64226
rect 547094 64170 547150 64226
rect 547218 64170 547274 64226
rect 547342 64170 547398 64226
rect 546970 64046 547026 64102
rect 547094 64046 547150 64102
rect 547218 64046 547274 64102
rect 547342 64046 547398 64102
rect 546970 63922 547026 63978
rect 547094 63922 547150 63978
rect 547218 63922 547274 63978
rect 547342 63922 547398 63978
rect 546970 46294 547026 46350
rect 547094 46294 547150 46350
rect 547218 46294 547274 46350
rect 547342 46294 547398 46350
rect 546970 46170 547026 46226
rect 547094 46170 547150 46226
rect 547218 46170 547274 46226
rect 547342 46170 547398 46226
rect 546970 46046 547026 46102
rect 547094 46046 547150 46102
rect 547218 46046 547274 46102
rect 547342 46046 547398 46102
rect 546970 45922 547026 45978
rect 547094 45922 547150 45978
rect 547218 45922 547274 45978
rect 547342 45922 547398 45978
rect 546970 28294 547026 28350
rect 547094 28294 547150 28350
rect 547218 28294 547274 28350
rect 547342 28294 547398 28350
rect 546970 28170 547026 28226
rect 547094 28170 547150 28226
rect 547218 28170 547274 28226
rect 547342 28170 547398 28226
rect 546970 28046 547026 28102
rect 547094 28046 547150 28102
rect 547218 28046 547274 28102
rect 547342 28046 547398 28102
rect 546970 27922 547026 27978
rect 547094 27922 547150 27978
rect 547218 27922 547274 27978
rect 547342 27922 547398 27978
rect 546970 10294 547026 10350
rect 547094 10294 547150 10350
rect 547218 10294 547274 10350
rect 547342 10294 547398 10350
rect 546970 10170 547026 10226
rect 547094 10170 547150 10226
rect 547218 10170 547274 10226
rect 547342 10170 547398 10226
rect 546970 10046 547026 10102
rect 547094 10046 547150 10102
rect 547218 10046 547274 10102
rect 547342 10046 547398 10102
rect 546970 9922 547026 9978
rect 547094 9922 547150 9978
rect 547218 9922 547274 9978
rect 547342 9922 547398 9978
rect 546970 -1176 547026 -1120
rect 547094 -1176 547150 -1120
rect 547218 -1176 547274 -1120
rect 547342 -1176 547398 -1120
rect 546970 -1300 547026 -1244
rect 547094 -1300 547150 -1244
rect 547218 -1300 547274 -1244
rect 547342 -1300 547398 -1244
rect 546970 -1424 547026 -1368
rect 547094 -1424 547150 -1368
rect 547218 -1424 547274 -1368
rect 547342 -1424 547398 -1368
rect 546970 -1548 547026 -1492
rect 547094 -1548 547150 -1492
rect 547218 -1548 547274 -1492
rect 547342 -1548 547398 -1492
rect 561250 597156 561306 597212
rect 561374 597156 561430 597212
rect 561498 597156 561554 597212
rect 561622 597156 561678 597212
rect 561250 597032 561306 597088
rect 561374 597032 561430 597088
rect 561498 597032 561554 597088
rect 561622 597032 561678 597088
rect 561250 596908 561306 596964
rect 561374 596908 561430 596964
rect 561498 596908 561554 596964
rect 561622 596908 561678 596964
rect 561250 596784 561306 596840
rect 561374 596784 561430 596840
rect 561498 596784 561554 596840
rect 561622 596784 561678 596840
rect 561250 580294 561306 580350
rect 561374 580294 561430 580350
rect 561498 580294 561554 580350
rect 561622 580294 561678 580350
rect 561250 580170 561306 580226
rect 561374 580170 561430 580226
rect 561498 580170 561554 580226
rect 561622 580170 561678 580226
rect 561250 580046 561306 580102
rect 561374 580046 561430 580102
rect 561498 580046 561554 580102
rect 561622 580046 561678 580102
rect 561250 579922 561306 579978
rect 561374 579922 561430 579978
rect 561498 579922 561554 579978
rect 561622 579922 561678 579978
rect 561250 562294 561306 562350
rect 561374 562294 561430 562350
rect 561498 562294 561554 562350
rect 561622 562294 561678 562350
rect 561250 562170 561306 562226
rect 561374 562170 561430 562226
rect 561498 562170 561554 562226
rect 561622 562170 561678 562226
rect 561250 562046 561306 562102
rect 561374 562046 561430 562102
rect 561498 562046 561554 562102
rect 561622 562046 561678 562102
rect 561250 561922 561306 561978
rect 561374 561922 561430 561978
rect 561498 561922 561554 561978
rect 561622 561922 561678 561978
rect 561250 544294 561306 544350
rect 561374 544294 561430 544350
rect 561498 544294 561554 544350
rect 561622 544294 561678 544350
rect 561250 544170 561306 544226
rect 561374 544170 561430 544226
rect 561498 544170 561554 544226
rect 561622 544170 561678 544226
rect 561250 544046 561306 544102
rect 561374 544046 561430 544102
rect 561498 544046 561554 544102
rect 561622 544046 561678 544102
rect 561250 543922 561306 543978
rect 561374 543922 561430 543978
rect 561498 543922 561554 543978
rect 561622 543922 561678 543978
rect 561250 526294 561306 526350
rect 561374 526294 561430 526350
rect 561498 526294 561554 526350
rect 561622 526294 561678 526350
rect 561250 526170 561306 526226
rect 561374 526170 561430 526226
rect 561498 526170 561554 526226
rect 561622 526170 561678 526226
rect 561250 526046 561306 526102
rect 561374 526046 561430 526102
rect 561498 526046 561554 526102
rect 561622 526046 561678 526102
rect 561250 525922 561306 525978
rect 561374 525922 561430 525978
rect 561498 525922 561554 525978
rect 561622 525922 561678 525978
rect 561250 508294 561306 508350
rect 561374 508294 561430 508350
rect 561498 508294 561554 508350
rect 561622 508294 561678 508350
rect 561250 508170 561306 508226
rect 561374 508170 561430 508226
rect 561498 508170 561554 508226
rect 561622 508170 561678 508226
rect 561250 508046 561306 508102
rect 561374 508046 561430 508102
rect 561498 508046 561554 508102
rect 561622 508046 561678 508102
rect 561250 507922 561306 507978
rect 561374 507922 561430 507978
rect 561498 507922 561554 507978
rect 561622 507922 561678 507978
rect 561250 490294 561306 490350
rect 561374 490294 561430 490350
rect 561498 490294 561554 490350
rect 561622 490294 561678 490350
rect 561250 490170 561306 490226
rect 561374 490170 561430 490226
rect 561498 490170 561554 490226
rect 561622 490170 561678 490226
rect 561250 490046 561306 490102
rect 561374 490046 561430 490102
rect 561498 490046 561554 490102
rect 561622 490046 561678 490102
rect 561250 489922 561306 489978
rect 561374 489922 561430 489978
rect 561498 489922 561554 489978
rect 561622 489922 561678 489978
rect 561250 472294 561306 472350
rect 561374 472294 561430 472350
rect 561498 472294 561554 472350
rect 561622 472294 561678 472350
rect 561250 472170 561306 472226
rect 561374 472170 561430 472226
rect 561498 472170 561554 472226
rect 561622 472170 561678 472226
rect 561250 472046 561306 472102
rect 561374 472046 561430 472102
rect 561498 472046 561554 472102
rect 561622 472046 561678 472102
rect 561250 471922 561306 471978
rect 561374 471922 561430 471978
rect 561498 471922 561554 471978
rect 561622 471922 561678 471978
rect 561250 454294 561306 454350
rect 561374 454294 561430 454350
rect 561498 454294 561554 454350
rect 561622 454294 561678 454350
rect 561250 454170 561306 454226
rect 561374 454170 561430 454226
rect 561498 454170 561554 454226
rect 561622 454170 561678 454226
rect 561250 454046 561306 454102
rect 561374 454046 561430 454102
rect 561498 454046 561554 454102
rect 561622 454046 561678 454102
rect 561250 453922 561306 453978
rect 561374 453922 561430 453978
rect 561498 453922 561554 453978
rect 561622 453922 561678 453978
rect 561250 436294 561306 436350
rect 561374 436294 561430 436350
rect 561498 436294 561554 436350
rect 561622 436294 561678 436350
rect 561250 436170 561306 436226
rect 561374 436170 561430 436226
rect 561498 436170 561554 436226
rect 561622 436170 561678 436226
rect 561250 436046 561306 436102
rect 561374 436046 561430 436102
rect 561498 436046 561554 436102
rect 561622 436046 561678 436102
rect 561250 435922 561306 435978
rect 561374 435922 561430 435978
rect 561498 435922 561554 435978
rect 561622 435922 561678 435978
rect 561250 418294 561306 418350
rect 561374 418294 561430 418350
rect 561498 418294 561554 418350
rect 561622 418294 561678 418350
rect 561250 418170 561306 418226
rect 561374 418170 561430 418226
rect 561498 418170 561554 418226
rect 561622 418170 561678 418226
rect 561250 418046 561306 418102
rect 561374 418046 561430 418102
rect 561498 418046 561554 418102
rect 561622 418046 561678 418102
rect 561250 417922 561306 417978
rect 561374 417922 561430 417978
rect 561498 417922 561554 417978
rect 561622 417922 561678 417978
rect 561250 400294 561306 400350
rect 561374 400294 561430 400350
rect 561498 400294 561554 400350
rect 561622 400294 561678 400350
rect 561250 400170 561306 400226
rect 561374 400170 561430 400226
rect 561498 400170 561554 400226
rect 561622 400170 561678 400226
rect 561250 400046 561306 400102
rect 561374 400046 561430 400102
rect 561498 400046 561554 400102
rect 561622 400046 561678 400102
rect 561250 399922 561306 399978
rect 561374 399922 561430 399978
rect 561498 399922 561554 399978
rect 561622 399922 561678 399978
rect 561250 382294 561306 382350
rect 561374 382294 561430 382350
rect 561498 382294 561554 382350
rect 561622 382294 561678 382350
rect 561250 382170 561306 382226
rect 561374 382170 561430 382226
rect 561498 382170 561554 382226
rect 561622 382170 561678 382226
rect 561250 382046 561306 382102
rect 561374 382046 561430 382102
rect 561498 382046 561554 382102
rect 561622 382046 561678 382102
rect 561250 381922 561306 381978
rect 561374 381922 561430 381978
rect 561498 381922 561554 381978
rect 561622 381922 561678 381978
rect 561250 364294 561306 364350
rect 561374 364294 561430 364350
rect 561498 364294 561554 364350
rect 561622 364294 561678 364350
rect 561250 364170 561306 364226
rect 561374 364170 561430 364226
rect 561498 364170 561554 364226
rect 561622 364170 561678 364226
rect 561250 364046 561306 364102
rect 561374 364046 561430 364102
rect 561498 364046 561554 364102
rect 561622 364046 561678 364102
rect 561250 363922 561306 363978
rect 561374 363922 561430 363978
rect 561498 363922 561554 363978
rect 561622 363922 561678 363978
rect 561250 346294 561306 346350
rect 561374 346294 561430 346350
rect 561498 346294 561554 346350
rect 561622 346294 561678 346350
rect 561250 346170 561306 346226
rect 561374 346170 561430 346226
rect 561498 346170 561554 346226
rect 561622 346170 561678 346226
rect 561250 346046 561306 346102
rect 561374 346046 561430 346102
rect 561498 346046 561554 346102
rect 561622 346046 561678 346102
rect 561250 345922 561306 345978
rect 561374 345922 561430 345978
rect 561498 345922 561554 345978
rect 561622 345922 561678 345978
rect 561250 328294 561306 328350
rect 561374 328294 561430 328350
rect 561498 328294 561554 328350
rect 561622 328294 561678 328350
rect 561250 328170 561306 328226
rect 561374 328170 561430 328226
rect 561498 328170 561554 328226
rect 561622 328170 561678 328226
rect 561250 328046 561306 328102
rect 561374 328046 561430 328102
rect 561498 328046 561554 328102
rect 561622 328046 561678 328102
rect 561250 327922 561306 327978
rect 561374 327922 561430 327978
rect 561498 327922 561554 327978
rect 561622 327922 561678 327978
rect 561250 310294 561306 310350
rect 561374 310294 561430 310350
rect 561498 310294 561554 310350
rect 561622 310294 561678 310350
rect 561250 310170 561306 310226
rect 561374 310170 561430 310226
rect 561498 310170 561554 310226
rect 561622 310170 561678 310226
rect 561250 310046 561306 310102
rect 561374 310046 561430 310102
rect 561498 310046 561554 310102
rect 561622 310046 561678 310102
rect 561250 309922 561306 309978
rect 561374 309922 561430 309978
rect 561498 309922 561554 309978
rect 561622 309922 561678 309978
rect 561250 292294 561306 292350
rect 561374 292294 561430 292350
rect 561498 292294 561554 292350
rect 561622 292294 561678 292350
rect 561250 292170 561306 292226
rect 561374 292170 561430 292226
rect 561498 292170 561554 292226
rect 561622 292170 561678 292226
rect 561250 292046 561306 292102
rect 561374 292046 561430 292102
rect 561498 292046 561554 292102
rect 561622 292046 561678 292102
rect 561250 291922 561306 291978
rect 561374 291922 561430 291978
rect 561498 291922 561554 291978
rect 561622 291922 561678 291978
rect 561250 274294 561306 274350
rect 561374 274294 561430 274350
rect 561498 274294 561554 274350
rect 561622 274294 561678 274350
rect 561250 274170 561306 274226
rect 561374 274170 561430 274226
rect 561498 274170 561554 274226
rect 561622 274170 561678 274226
rect 561250 274046 561306 274102
rect 561374 274046 561430 274102
rect 561498 274046 561554 274102
rect 561622 274046 561678 274102
rect 561250 273922 561306 273978
rect 561374 273922 561430 273978
rect 561498 273922 561554 273978
rect 561622 273922 561678 273978
rect 561250 256294 561306 256350
rect 561374 256294 561430 256350
rect 561498 256294 561554 256350
rect 561622 256294 561678 256350
rect 561250 256170 561306 256226
rect 561374 256170 561430 256226
rect 561498 256170 561554 256226
rect 561622 256170 561678 256226
rect 561250 256046 561306 256102
rect 561374 256046 561430 256102
rect 561498 256046 561554 256102
rect 561622 256046 561678 256102
rect 561250 255922 561306 255978
rect 561374 255922 561430 255978
rect 561498 255922 561554 255978
rect 561622 255922 561678 255978
rect 561250 238294 561306 238350
rect 561374 238294 561430 238350
rect 561498 238294 561554 238350
rect 561622 238294 561678 238350
rect 561250 238170 561306 238226
rect 561374 238170 561430 238226
rect 561498 238170 561554 238226
rect 561622 238170 561678 238226
rect 561250 238046 561306 238102
rect 561374 238046 561430 238102
rect 561498 238046 561554 238102
rect 561622 238046 561678 238102
rect 561250 237922 561306 237978
rect 561374 237922 561430 237978
rect 561498 237922 561554 237978
rect 561622 237922 561678 237978
rect 561250 220294 561306 220350
rect 561374 220294 561430 220350
rect 561498 220294 561554 220350
rect 561622 220294 561678 220350
rect 561250 220170 561306 220226
rect 561374 220170 561430 220226
rect 561498 220170 561554 220226
rect 561622 220170 561678 220226
rect 561250 220046 561306 220102
rect 561374 220046 561430 220102
rect 561498 220046 561554 220102
rect 561622 220046 561678 220102
rect 561250 219922 561306 219978
rect 561374 219922 561430 219978
rect 561498 219922 561554 219978
rect 561622 219922 561678 219978
rect 561250 202294 561306 202350
rect 561374 202294 561430 202350
rect 561498 202294 561554 202350
rect 561622 202294 561678 202350
rect 561250 202170 561306 202226
rect 561374 202170 561430 202226
rect 561498 202170 561554 202226
rect 561622 202170 561678 202226
rect 561250 202046 561306 202102
rect 561374 202046 561430 202102
rect 561498 202046 561554 202102
rect 561622 202046 561678 202102
rect 561250 201922 561306 201978
rect 561374 201922 561430 201978
rect 561498 201922 561554 201978
rect 561622 201922 561678 201978
rect 561250 184294 561306 184350
rect 561374 184294 561430 184350
rect 561498 184294 561554 184350
rect 561622 184294 561678 184350
rect 561250 184170 561306 184226
rect 561374 184170 561430 184226
rect 561498 184170 561554 184226
rect 561622 184170 561678 184226
rect 561250 184046 561306 184102
rect 561374 184046 561430 184102
rect 561498 184046 561554 184102
rect 561622 184046 561678 184102
rect 561250 183922 561306 183978
rect 561374 183922 561430 183978
rect 561498 183922 561554 183978
rect 561622 183922 561678 183978
rect 561250 166294 561306 166350
rect 561374 166294 561430 166350
rect 561498 166294 561554 166350
rect 561622 166294 561678 166350
rect 561250 166170 561306 166226
rect 561374 166170 561430 166226
rect 561498 166170 561554 166226
rect 561622 166170 561678 166226
rect 561250 166046 561306 166102
rect 561374 166046 561430 166102
rect 561498 166046 561554 166102
rect 561622 166046 561678 166102
rect 561250 165922 561306 165978
rect 561374 165922 561430 165978
rect 561498 165922 561554 165978
rect 561622 165922 561678 165978
rect 561250 148294 561306 148350
rect 561374 148294 561430 148350
rect 561498 148294 561554 148350
rect 561622 148294 561678 148350
rect 561250 148170 561306 148226
rect 561374 148170 561430 148226
rect 561498 148170 561554 148226
rect 561622 148170 561678 148226
rect 561250 148046 561306 148102
rect 561374 148046 561430 148102
rect 561498 148046 561554 148102
rect 561622 148046 561678 148102
rect 561250 147922 561306 147978
rect 561374 147922 561430 147978
rect 561498 147922 561554 147978
rect 561622 147922 561678 147978
rect 561250 130294 561306 130350
rect 561374 130294 561430 130350
rect 561498 130294 561554 130350
rect 561622 130294 561678 130350
rect 561250 130170 561306 130226
rect 561374 130170 561430 130226
rect 561498 130170 561554 130226
rect 561622 130170 561678 130226
rect 561250 130046 561306 130102
rect 561374 130046 561430 130102
rect 561498 130046 561554 130102
rect 561622 130046 561678 130102
rect 561250 129922 561306 129978
rect 561374 129922 561430 129978
rect 561498 129922 561554 129978
rect 561622 129922 561678 129978
rect 561250 112294 561306 112350
rect 561374 112294 561430 112350
rect 561498 112294 561554 112350
rect 561622 112294 561678 112350
rect 561250 112170 561306 112226
rect 561374 112170 561430 112226
rect 561498 112170 561554 112226
rect 561622 112170 561678 112226
rect 561250 112046 561306 112102
rect 561374 112046 561430 112102
rect 561498 112046 561554 112102
rect 561622 112046 561678 112102
rect 561250 111922 561306 111978
rect 561374 111922 561430 111978
rect 561498 111922 561554 111978
rect 561622 111922 561678 111978
rect 561250 94294 561306 94350
rect 561374 94294 561430 94350
rect 561498 94294 561554 94350
rect 561622 94294 561678 94350
rect 561250 94170 561306 94226
rect 561374 94170 561430 94226
rect 561498 94170 561554 94226
rect 561622 94170 561678 94226
rect 561250 94046 561306 94102
rect 561374 94046 561430 94102
rect 561498 94046 561554 94102
rect 561622 94046 561678 94102
rect 561250 93922 561306 93978
rect 561374 93922 561430 93978
rect 561498 93922 561554 93978
rect 561622 93922 561678 93978
rect 561250 76294 561306 76350
rect 561374 76294 561430 76350
rect 561498 76294 561554 76350
rect 561622 76294 561678 76350
rect 561250 76170 561306 76226
rect 561374 76170 561430 76226
rect 561498 76170 561554 76226
rect 561622 76170 561678 76226
rect 561250 76046 561306 76102
rect 561374 76046 561430 76102
rect 561498 76046 561554 76102
rect 561622 76046 561678 76102
rect 561250 75922 561306 75978
rect 561374 75922 561430 75978
rect 561498 75922 561554 75978
rect 561622 75922 561678 75978
rect 561250 58294 561306 58350
rect 561374 58294 561430 58350
rect 561498 58294 561554 58350
rect 561622 58294 561678 58350
rect 561250 58170 561306 58226
rect 561374 58170 561430 58226
rect 561498 58170 561554 58226
rect 561622 58170 561678 58226
rect 561250 58046 561306 58102
rect 561374 58046 561430 58102
rect 561498 58046 561554 58102
rect 561622 58046 561678 58102
rect 561250 57922 561306 57978
rect 561374 57922 561430 57978
rect 561498 57922 561554 57978
rect 561622 57922 561678 57978
rect 561250 40294 561306 40350
rect 561374 40294 561430 40350
rect 561498 40294 561554 40350
rect 561622 40294 561678 40350
rect 561250 40170 561306 40226
rect 561374 40170 561430 40226
rect 561498 40170 561554 40226
rect 561622 40170 561678 40226
rect 561250 40046 561306 40102
rect 561374 40046 561430 40102
rect 561498 40046 561554 40102
rect 561622 40046 561678 40102
rect 561250 39922 561306 39978
rect 561374 39922 561430 39978
rect 561498 39922 561554 39978
rect 561622 39922 561678 39978
rect 561250 22294 561306 22350
rect 561374 22294 561430 22350
rect 561498 22294 561554 22350
rect 561622 22294 561678 22350
rect 561250 22170 561306 22226
rect 561374 22170 561430 22226
rect 561498 22170 561554 22226
rect 561622 22170 561678 22226
rect 561250 22046 561306 22102
rect 561374 22046 561430 22102
rect 561498 22046 561554 22102
rect 561622 22046 561678 22102
rect 561250 21922 561306 21978
rect 561374 21922 561430 21978
rect 561498 21922 561554 21978
rect 561622 21922 561678 21978
rect 561250 4294 561306 4350
rect 561374 4294 561430 4350
rect 561498 4294 561554 4350
rect 561622 4294 561678 4350
rect 561250 4170 561306 4226
rect 561374 4170 561430 4226
rect 561498 4170 561554 4226
rect 561622 4170 561678 4226
rect 561250 4046 561306 4102
rect 561374 4046 561430 4102
rect 561498 4046 561554 4102
rect 561622 4046 561678 4102
rect 561250 3922 561306 3978
rect 561374 3922 561430 3978
rect 561498 3922 561554 3978
rect 561622 3922 561678 3978
rect 561250 -216 561306 -160
rect 561374 -216 561430 -160
rect 561498 -216 561554 -160
rect 561622 -216 561678 -160
rect 561250 -340 561306 -284
rect 561374 -340 561430 -284
rect 561498 -340 561554 -284
rect 561622 -340 561678 -284
rect 561250 -464 561306 -408
rect 561374 -464 561430 -408
rect 561498 -464 561554 -408
rect 561622 -464 561678 -408
rect 561250 -588 561306 -532
rect 561374 -588 561430 -532
rect 561498 -588 561554 -532
rect 561622 -588 561678 -532
rect 564970 598116 565026 598172
rect 565094 598116 565150 598172
rect 565218 598116 565274 598172
rect 565342 598116 565398 598172
rect 564970 597992 565026 598048
rect 565094 597992 565150 598048
rect 565218 597992 565274 598048
rect 565342 597992 565398 598048
rect 564970 597868 565026 597924
rect 565094 597868 565150 597924
rect 565218 597868 565274 597924
rect 565342 597868 565398 597924
rect 564970 597744 565026 597800
rect 565094 597744 565150 597800
rect 565218 597744 565274 597800
rect 565342 597744 565398 597800
rect 564970 586294 565026 586350
rect 565094 586294 565150 586350
rect 565218 586294 565274 586350
rect 565342 586294 565398 586350
rect 564970 586170 565026 586226
rect 565094 586170 565150 586226
rect 565218 586170 565274 586226
rect 565342 586170 565398 586226
rect 564970 586046 565026 586102
rect 565094 586046 565150 586102
rect 565218 586046 565274 586102
rect 565342 586046 565398 586102
rect 564970 585922 565026 585978
rect 565094 585922 565150 585978
rect 565218 585922 565274 585978
rect 565342 585922 565398 585978
rect 564970 568294 565026 568350
rect 565094 568294 565150 568350
rect 565218 568294 565274 568350
rect 565342 568294 565398 568350
rect 564970 568170 565026 568226
rect 565094 568170 565150 568226
rect 565218 568170 565274 568226
rect 565342 568170 565398 568226
rect 564970 568046 565026 568102
rect 565094 568046 565150 568102
rect 565218 568046 565274 568102
rect 565342 568046 565398 568102
rect 564970 567922 565026 567978
rect 565094 567922 565150 567978
rect 565218 567922 565274 567978
rect 565342 567922 565398 567978
rect 564970 550294 565026 550350
rect 565094 550294 565150 550350
rect 565218 550294 565274 550350
rect 565342 550294 565398 550350
rect 564970 550170 565026 550226
rect 565094 550170 565150 550226
rect 565218 550170 565274 550226
rect 565342 550170 565398 550226
rect 564970 550046 565026 550102
rect 565094 550046 565150 550102
rect 565218 550046 565274 550102
rect 565342 550046 565398 550102
rect 564970 549922 565026 549978
rect 565094 549922 565150 549978
rect 565218 549922 565274 549978
rect 565342 549922 565398 549978
rect 564970 532294 565026 532350
rect 565094 532294 565150 532350
rect 565218 532294 565274 532350
rect 565342 532294 565398 532350
rect 564970 532170 565026 532226
rect 565094 532170 565150 532226
rect 565218 532170 565274 532226
rect 565342 532170 565398 532226
rect 564970 532046 565026 532102
rect 565094 532046 565150 532102
rect 565218 532046 565274 532102
rect 565342 532046 565398 532102
rect 564970 531922 565026 531978
rect 565094 531922 565150 531978
rect 565218 531922 565274 531978
rect 565342 531922 565398 531978
rect 564970 514294 565026 514350
rect 565094 514294 565150 514350
rect 565218 514294 565274 514350
rect 565342 514294 565398 514350
rect 564970 514170 565026 514226
rect 565094 514170 565150 514226
rect 565218 514170 565274 514226
rect 565342 514170 565398 514226
rect 564970 514046 565026 514102
rect 565094 514046 565150 514102
rect 565218 514046 565274 514102
rect 565342 514046 565398 514102
rect 564970 513922 565026 513978
rect 565094 513922 565150 513978
rect 565218 513922 565274 513978
rect 565342 513922 565398 513978
rect 564970 496294 565026 496350
rect 565094 496294 565150 496350
rect 565218 496294 565274 496350
rect 565342 496294 565398 496350
rect 564970 496170 565026 496226
rect 565094 496170 565150 496226
rect 565218 496170 565274 496226
rect 565342 496170 565398 496226
rect 564970 496046 565026 496102
rect 565094 496046 565150 496102
rect 565218 496046 565274 496102
rect 565342 496046 565398 496102
rect 564970 495922 565026 495978
rect 565094 495922 565150 495978
rect 565218 495922 565274 495978
rect 565342 495922 565398 495978
rect 564970 478294 565026 478350
rect 565094 478294 565150 478350
rect 565218 478294 565274 478350
rect 565342 478294 565398 478350
rect 564970 478170 565026 478226
rect 565094 478170 565150 478226
rect 565218 478170 565274 478226
rect 565342 478170 565398 478226
rect 564970 478046 565026 478102
rect 565094 478046 565150 478102
rect 565218 478046 565274 478102
rect 565342 478046 565398 478102
rect 564970 477922 565026 477978
rect 565094 477922 565150 477978
rect 565218 477922 565274 477978
rect 565342 477922 565398 477978
rect 564970 460294 565026 460350
rect 565094 460294 565150 460350
rect 565218 460294 565274 460350
rect 565342 460294 565398 460350
rect 564970 460170 565026 460226
rect 565094 460170 565150 460226
rect 565218 460170 565274 460226
rect 565342 460170 565398 460226
rect 564970 460046 565026 460102
rect 565094 460046 565150 460102
rect 565218 460046 565274 460102
rect 565342 460046 565398 460102
rect 564970 459922 565026 459978
rect 565094 459922 565150 459978
rect 565218 459922 565274 459978
rect 565342 459922 565398 459978
rect 564970 442294 565026 442350
rect 565094 442294 565150 442350
rect 565218 442294 565274 442350
rect 565342 442294 565398 442350
rect 564970 442170 565026 442226
rect 565094 442170 565150 442226
rect 565218 442170 565274 442226
rect 565342 442170 565398 442226
rect 564970 442046 565026 442102
rect 565094 442046 565150 442102
rect 565218 442046 565274 442102
rect 565342 442046 565398 442102
rect 564970 441922 565026 441978
rect 565094 441922 565150 441978
rect 565218 441922 565274 441978
rect 565342 441922 565398 441978
rect 564970 424294 565026 424350
rect 565094 424294 565150 424350
rect 565218 424294 565274 424350
rect 565342 424294 565398 424350
rect 564970 424170 565026 424226
rect 565094 424170 565150 424226
rect 565218 424170 565274 424226
rect 565342 424170 565398 424226
rect 564970 424046 565026 424102
rect 565094 424046 565150 424102
rect 565218 424046 565274 424102
rect 565342 424046 565398 424102
rect 564970 423922 565026 423978
rect 565094 423922 565150 423978
rect 565218 423922 565274 423978
rect 565342 423922 565398 423978
rect 564970 406294 565026 406350
rect 565094 406294 565150 406350
rect 565218 406294 565274 406350
rect 565342 406294 565398 406350
rect 564970 406170 565026 406226
rect 565094 406170 565150 406226
rect 565218 406170 565274 406226
rect 565342 406170 565398 406226
rect 564970 406046 565026 406102
rect 565094 406046 565150 406102
rect 565218 406046 565274 406102
rect 565342 406046 565398 406102
rect 564970 405922 565026 405978
rect 565094 405922 565150 405978
rect 565218 405922 565274 405978
rect 565342 405922 565398 405978
rect 564970 388294 565026 388350
rect 565094 388294 565150 388350
rect 565218 388294 565274 388350
rect 565342 388294 565398 388350
rect 564970 388170 565026 388226
rect 565094 388170 565150 388226
rect 565218 388170 565274 388226
rect 565342 388170 565398 388226
rect 564970 388046 565026 388102
rect 565094 388046 565150 388102
rect 565218 388046 565274 388102
rect 565342 388046 565398 388102
rect 564970 387922 565026 387978
rect 565094 387922 565150 387978
rect 565218 387922 565274 387978
rect 565342 387922 565398 387978
rect 564970 370294 565026 370350
rect 565094 370294 565150 370350
rect 565218 370294 565274 370350
rect 565342 370294 565398 370350
rect 564970 370170 565026 370226
rect 565094 370170 565150 370226
rect 565218 370170 565274 370226
rect 565342 370170 565398 370226
rect 564970 370046 565026 370102
rect 565094 370046 565150 370102
rect 565218 370046 565274 370102
rect 565342 370046 565398 370102
rect 564970 369922 565026 369978
rect 565094 369922 565150 369978
rect 565218 369922 565274 369978
rect 565342 369922 565398 369978
rect 564970 352294 565026 352350
rect 565094 352294 565150 352350
rect 565218 352294 565274 352350
rect 565342 352294 565398 352350
rect 564970 352170 565026 352226
rect 565094 352170 565150 352226
rect 565218 352170 565274 352226
rect 565342 352170 565398 352226
rect 564970 352046 565026 352102
rect 565094 352046 565150 352102
rect 565218 352046 565274 352102
rect 565342 352046 565398 352102
rect 564970 351922 565026 351978
rect 565094 351922 565150 351978
rect 565218 351922 565274 351978
rect 565342 351922 565398 351978
rect 564970 334294 565026 334350
rect 565094 334294 565150 334350
rect 565218 334294 565274 334350
rect 565342 334294 565398 334350
rect 564970 334170 565026 334226
rect 565094 334170 565150 334226
rect 565218 334170 565274 334226
rect 565342 334170 565398 334226
rect 564970 334046 565026 334102
rect 565094 334046 565150 334102
rect 565218 334046 565274 334102
rect 565342 334046 565398 334102
rect 564970 333922 565026 333978
rect 565094 333922 565150 333978
rect 565218 333922 565274 333978
rect 565342 333922 565398 333978
rect 564970 316294 565026 316350
rect 565094 316294 565150 316350
rect 565218 316294 565274 316350
rect 565342 316294 565398 316350
rect 564970 316170 565026 316226
rect 565094 316170 565150 316226
rect 565218 316170 565274 316226
rect 565342 316170 565398 316226
rect 564970 316046 565026 316102
rect 565094 316046 565150 316102
rect 565218 316046 565274 316102
rect 565342 316046 565398 316102
rect 564970 315922 565026 315978
rect 565094 315922 565150 315978
rect 565218 315922 565274 315978
rect 565342 315922 565398 315978
rect 564970 298294 565026 298350
rect 565094 298294 565150 298350
rect 565218 298294 565274 298350
rect 565342 298294 565398 298350
rect 564970 298170 565026 298226
rect 565094 298170 565150 298226
rect 565218 298170 565274 298226
rect 565342 298170 565398 298226
rect 564970 298046 565026 298102
rect 565094 298046 565150 298102
rect 565218 298046 565274 298102
rect 565342 298046 565398 298102
rect 564970 297922 565026 297978
rect 565094 297922 565150 297978
rect 565218 297922 565274 297978
rect 565342 297922 565398 297978
rect 564970 280294 565026 280350
rect 565094 280294 565150 280350
rect 565218 280294 565274 280350
rect 565342 280294 565398 280350
rect 564970 280170 565026 280226
rect 565094 280170 565150 280226
rect 565218 280170 565274 280226
rect 565342 280170 565398 280226
rect 564970 280046 565026 280102
rect 565094 280046 565150 280102
rect 565218 280046 565274 280102
rect 565342 280046 565398 280102
rect 564970 279922 565026 279978
rect 565094 279922 565150 279978
rect 565218 279922 565274 279978
rect 565342 279922 565398 279978
rect 564970 262294 565026 262350
rect 565094 262294 565150 262350
rect 565218 262294 565274 262350
rect 565342 262294 565398 262350
rect 564970 262170 565026 262226
rect 565094 262170 565150 262226
rect 565218 262170 565274 262226
rect 565342 262170 565398 262226
rect 564970 262046 565026 262102
rect 565094 262046 565150 262102
rect 565218 262046 565274 262102
rect 565342 262046 565398 262102
rect 564970 261922 565026 261978
rect 565094 261922 565150 261978
rect 565218 261922 565274 261978
rect 565342 261922 565398 261978
rect 564970 244294 565026 244350
rect 565094 244294 565150 244350
rect 565218 244294 565274 244350
rect 565342 244294 565398 244350
rect 564970 244170 565026 244226
rect 565094 244170 565150 244226
rect 565218 244170 565274 244226
rect 565342 244170 565398 244226
rect 564970 244046 565026 244102
rect 565094 244046 565150 244102
rect 565218 244046 565274 244102
rect 565342 244046 565398 244102
rect 564970 243922 565026 243978
rect 565094 243922 565150 243978
rect 565218 243922 565274 243978
rect 565342 243922 565398 243978
rect 564970 226294 565026 226350
rect 565094 226294 565150 226350
rect 565218 226294 565274 226350
rect 565342 226294 565398 226350
rect 564970 226170 565026 226226
rect 565094 226170 565150 226226
rect 565218 226170 565274 226226
rect 565342 226170 565398 226226
rect 564970 226046 565026 226102
rect 565094 226046 565150 226102
rect 565218 226046 565274 226102
rect 565342 226046 565398 226102
rect 564970 225922 565026 225978
rect 565094 225922 565150 225978
rect 565218 225922 565274 225978
rect 565342 225922 565398 225978
rect 564970 208294 565026 208350
rect 565094 208294 565150 208350
rect 565218 208294 565274 208350
rect 565342 208294 565398 208350
rect 564970 208170 565026 208226
rect 565094 208170 565150 208226
rect 565218 208170 565274 208226
rect 565342 208170 565398 208226
rect 564970 208046 565026 208102
rect 565094 208046 565150 208102
rect 565218 208046 565274 208102
rect 565342 208046 565398 208102
rect 564970 207922 565026 207978
rect 565094 207922 565150 207978
rect 565218 207922 565274 207978
rect 565342 207922 565398 207978
rect 564970 190294 565026 190350
rect 565094 190294 565150 190350
rect 565218 190294 565274 190350
rect 565342 190294 565398 190350
rect 564970 190170 565026 190226
rect 565094 190170 565150 190226
rect 565218 190170 565274 190226
rect 565342 190170 565398 190226
rect 564970 190046 565026 190102
rect 565094 190046 565150 190102
rect 565218 190046 565274 190102
rect 565342 190046 565398 190102
rect 564970 189922 565026 189978
rect 565094 189922 565150 189978
rect 565218 189922 565274 189978
rect 565342 189922 565398 189978
rect 564970 172294 565026 172350
rect 565094 172294 565150 172350
rect 565218 172294 565274 172350
rect 565342 172294 565398 172350
rect 564970 172170 565026 172226
rect 565094 172170 565150 172226
rect 565218 172170 565274 172226
rect 565342 172170 565398 172226
rect 564970 172046 565026 172102
rect 565094 172046 565150 172102
rect 565218 172046 565274 172102
rect 565342 172046 565398 172102
rect 564970 171922 565026 171978
rect 565094 171922 565150 171978
rect 565218 171922 565274 171978
rect 565342 171922 565398 171978
rect 564970 154294 565026 154350
rect 565094 154294 565150 154350
rect 565218 154294 565274 154350
rect 565342 154294 565398 154350
rect 564970 154170 565026 154226
rect 565094 154170 565150 154226
rect 565218 154170 565274 154226
rect 565342 154170 565398 154226
rect 564970 154046 565026 154102
rect 565094 154046 565150 154102
rect 565218 154046 565274 154102
rect 565342 154046 565398 154102
rect 564970 153922 565026 153978
rect 565094 153922 565150 153978
rect 565218 153922 565274 153978
rect 565342 153922 565398 153978
rect 564970 136294 565026 136350
rect 565094 136294 565150 136350
rect 565218 136294 565274 136350
rect 565342 136294 565398 136350
rect 564970 136170 565026 136226
rect 565094 136170 565150 136226
rect 565218 136170 565274 136226
rect 565342 136170 565398 136226
rect 564970 136046 565026 136102
rect 565094 136046 565150 136102
rect 565218 136046 565274 136102
rect 565342 136046 565398 136102
rect 564970 135922 565026 135978
rect 565094 135922 565150 135978
rect 565218 135922 565274 135978
rect 565342 135922 565398 135978
rect 564970 118294 565026 118350
rect 565094 118294 565150 118350
rect 565218 118294 565274 118350
rect 565342 118294 565398 118350
rect 564970 118170 565026 118226
rect 565094 118170 565150 118226
rect 565218 118170 565274 118226
rect 565342 118170 565398 118226
rect 564970 118046 565026 118102
rect 565094 118046 565150 118102
rect 565218 118046 565274 118102
rect 565342 118046 565398 118102
rect 564970 117922 565026 117978
rect 565094 117922 565150 117978
rect 565218 117922 565274 117978
rect 565342 117922 565398 117978
rect 564970 100294 565026 100350
rect 565094 100294 565150 100350
rect 565218 100294 565274 100350
rect 565342 100294 565398 100350
rect 564970 100170 565026 100226
rect 565094 100170 565150 100226
rect 565218 100170 565274 100226
rect 565342 100170 565398 100226
rect 564970 100046 565026 100102
rect 565094 100046 565150 100102
rect 565218 100046 565274 100102
rect 565342 100046 565398 100102
rect 564970 99922 565026 99978
rect 565094 99922 565150 99978
rect 565218 99922 565274 99978
rect 565342 99922 565398 99978
rect 564970 82294 565026 82350
rect 565094 82294 565150 82350
rect 565218 82294 565274 82350
rect 565342 82294 565398 82350
rect 564970 82170 565026 82226
rect 565094 82170 565150 82226
rect 565218 82170 565274 82226
rect 565342 82170 565398 82226
rect 564970 82046 565026 82102
rect 565094 82046 565150 82102
rect 565218 82046 565274 82102
rect 565342 82046 565398 82102
rect 564970 81922 565026 81978
rect 565094 81922 565150 81978
rect 565218 81922 565274 81978
rect 565342 81922 565398 81978
rect 564970 64294 565026 64350
rect 565094 64294 565150 64350
rect 565218 64294 565274 64350
rect 565342 64294 565398 64350
rect 564970 64170 565026 64226
rect 565094 64170 565150 64226
rect 565218 64170 565274 64226
rect 565342 64170 565398 64226
rect 564970 64046 565026 64102
rect 565094 64046 565150 64102
rect 565218 64046 565274 64102
rect 565342 64046 565398 64102
rect 564970 63922 565026 63978
rect 565094 63922 565150 63978
rect 565218 63922 565274 63978
rect 565342 63922 565398 63978
rect 564970 46294 565026 46350
rect 565094 46294 565150 46350
rect 565218 46294 565274 46350
rect 565342 46294 565398 46350
rect 564970 46170 565026 46226
rect 565094 46170 565150 46226
rect 565218 46170 565274 46226
rect 565342 46170 565398 46226
rect 564970 46046 565026 46102
rect 565094 46046 565150 46102
rect 565218 46046 565274 46102
rect 565342 46046 565398 46102
rect 564970 45922 565026 45978
rect 565094 45922 565150 45978
rect 565218 45922 565274 45978
rect 565342 45922 565398 45978
rect 564970 28294 565026 28350
rect 565094 28294 565150 28350
rect 565218 28294 565274 28350
rect 565342 28294 565398 28350
rect 564970 28170 565026 28226
rect 565094 28170 565150 28226
rect 565218 28170 565274 28226
rect 565342 28170 565398 28226
rect 564970 28046 565026 28102
rect 565094 28046 565150 28102
rect 565218 28046 565274 28102
rect 565342 28046 565398 28102
rect 564970 27922 565026 27978
rect 565094 27922 565150 27978
rect 565218 27922 565274 27978
rect 565342 27922 565398 27978
rect 564970 10294 565026 10350
rect 565094 10294 565150 10350
rect 565218 10294 565274 10350
rect 565342 10294 565398 10350
rect 564970 10170 565026 10226
rect 565094 10170 565150 10226
rect 565218 10170 565274 10226
rect 565342 10170 565398 10226
rect 564970 10046 565026 10102
rect 565094 10046 565150 10102
rect 565218 10046 565274 10102
rect 565342 10046 565398 10102
rect 564970 9922 565026 9978
rect 565094 9922 565150 9978
rect 565218 9922 565274 9978
rect 565342 9922 565398 9978
rect 564970 -1176 565026 -1120
rect 565094 -1176 565150 -1120
rect 565218 -1176 565274 -1120
rect 565342 -1176 565398 -1120
rect 564970 -1300 565026 -1244
rect 565094 -1300 565150 -1244
rect 565218 -1300 565274 -1244
rect 565342 -1300 565398 -1244
rect 564970 -1424 565026 -1368
rect 565094 -1424 565150 -1368
rect 565218 -1424 565274 -1368
rect 565342 -1424 565398 -1368
rect 564970 -1548 565026 -1492
rect 565094 -1548 565150 -1492
rect 565218 -1548 565274 -1492
rect 565342 -1548 565398 -1492
rect 579250 597156 579306 597212
rect 579374 597156 579430 597212
rect 579498 597156 579554 597212
rect 579622 597156 579678 597212
rect 579250 597032 579306 597088
rect 579374 597032 579430 597088
rect 579498 597032 579554 597088
rect 579622 597032 579678 597088
rect 579250 596908 579306 596964
rect 579374 596908 579430 596964
rect 579498 596908 579554 596964
rect 579622 596908 579678 596964
rect 579250 596784 579306 596840
rect 579374 596784 579430 596840
rect 579498 596784 579554 596840
rect 579622 596784 579678 596840
rect 579250 580294 579306 580350
rect 579374 580294 579430 580350
rect 579498 580294 579554 580350
rect 579622 580294 579678 580350
rect 579250 580170 579306 580226
rect 579374 580170 579430 580226
rect 579498 580170 579554 580226
rect 579622 580170 579678 580226
rect 579250 580046 579306 580102
rect 579374 580046 579430 580102
rect 579498 580046 579554 580102
rect 579622 580046 579678 580102
rect 579250 579922 579306 579978
rect 579374 579922 579430 579978
rect 579498 579922 579554 579978
rect 579622 579922 579678 579978
rect 579250 562294 579306 562350
rect 579374 562294 579430 562350
rect 579498 562294 579554 562350
rect 579622 562294 579678 562350
rect 579250 562170 579306 562226
rect 579374 562170 579430 562226
rect 579498 562170 579554 562226
rect 579622 562170 579678 562226
rect 579250 562046 579306 562102
rect 579374 562046 579430 562102
rect 579498 562046 579554 562102
rect 579622 562046 579678 562102
rect 579250 561922 579306 561978
rect 579374 561922 579430 561978
rect 579498 561922 579554 561978
rect 579622 561922 579678 561978
rect 579250 544294 579306 544350
rect 579374 544294 579430 544350
rect 579498 544294 579554 544350
rect 579622 544294 579678 544350
rect 579250 544170 579306 544226
rect 579374 544170 579430 544226
rect 579498 544170 579554 544226
rect 579622 544170 579678 544226
rect 579250 544046 579306 544102
rect 579374 544046 579430 544102
rect 579498 544046 579554 544102
rect 579622 544046 579678 544102
rect 579250 543922 579306 543978
rect 579374 543922 579430 543978
rect 579498 543922 579554 543978
rect 579622 543922 579678 543978
rect 579250 526294 579306 526350
rect 579374 526294 579430 526350
rect 579498 526294 579554 526350
rect 579622 526294 579678 526350
rect 579250 526170 579306 526226
rect 579374 526170 579430 526226
rect 579498 526170 579554 526226
rect 579622 526170 579678 526226
rect 579250 526046 579306 526102
rect 579374 526046 579430 526102
rect 579498 526046 579554 526102
rect 579622 526046 579678 526102
rect 579250 525922 579306 525978
rect 579374 525922 579430 525978
rect 579498 525922 579554 525978
rect 579622 525922 579678 525978
rect 579250 508294 579306 508350
rect 579374 508294 579430 508350
rect 579498 508294 579554 508350
rect 579622 508294 579678 508350
rect 579250 508170 579306 508226
rect 579374 508170 579430 508226
rect 579498 508170 579554 508226
rect 579622 508170 579678 508226
rect 579250 508046 579306 508102
rect 579374 508046 579430 508102
rect 579498 508046 579554 508102
rect 579622 508046 579678 508102
rect 579250 507922 579306 507978
rect 579374 507922 579430 507978
rect 579498 507922 579554 507978
rect 579622 507922 579678 507978
rect 579250 490294 579306 490350
rect 579374 490294 579430 490350
rect 579498 490294 579554 490350
rect 579622 490294 579678 490350
rect 579250 490170 579306 490226
rect 579374 490170 579430 490226
rect 579498 490170 579554 490226
rect 579622 490170 579678 490226
rect 579250 490046 579306 490102
rect 579374 490046 579430 490102
rect 579498 490046 579554 490102
rect 579622 490046 579678 490102
rect 579250 489922 579306 489978
rect 579374 489922 579430 489978
rect 579498 489922 579554 489978
rect 579622 489922 579678 489978
rect 579250 472294 579306 472350
rect 579374 472294 579430 472350
rect 579498 472294 579554 472350
rect 579622 472294 579678 472350
rect 579250 472170 579306 472226
rect 579374 472170 579430 472226
rect 579498 472170 579554 472226
rect 579622 472170 579678 472226
rect 579250 472046 579306 472102
rect 579374 472046 579430 472102
rect 579498 472046 579554 472102
rect 579622 472046 579678 472102
rect 579250 471922 579306 471978
rect 579374 471922 579430 471978
rect 579498 471922 579554 471978
rect 579622 471922 579678 471978
rect 579250 454294 579306 454350
rect 579374 454294 579430 454350
rect 579498 454294 579554 454350
rect 579622 454294 579678 454350
rect 579250 454170 579306 454226
rect 579374 454170 579430 454226
rect 579498 454170 579554 454226
rect 579622 454170 579678 454226
rect 579250 454046 579306 454102
rect 579374 454046 579430 454102
rect 579498 454046 579554 454102
rect 579622 454046 579678 454102
rect 579250 453922 579306 453978
rect 579374 453922 579430 453978
rect 579498 453922 579554 453978
rect 579622 453922 579678 453978
rect 579250 436294 579306 436350
rect 579374 436294 579430 436350
rect 579498 436294 579554 436350
rect 579622 436294 579678 436350
rect 579250 436170 579306 436226
rect 579374 436170 579430 436226
rect 579498 436170 579554 436226
rect 579622 436170 579678 436226
rect 579250 436046 579306 436102
rect 579374 436046 579430 436102
rect 579498 436046 579554 436102
rect 579622 436046 579678 436102
rect 579250 435922 579306 435978
rect 579374 435922 579430 435978
rect 579498 435922 579554 435978
rect 579622 435922 579678 435978
rect 579250 418294 579306 418350
rect 579374 418294 579430 418350
rect 579498 418294 579554 418350
rect 579622 418294 579678 418350
rect 579250 418170 579306 418226
rect 579374 418170 579430 418226
rect 579498 418170 579554 418226
rect 579622 418170 579678 418226
rect 579250 418046 579306 418102
rect 579374 418046 579430 418102
rect 579498 418046 579554 418102
rect 579622 418046 579678 418102
rect 579250 417922 579306 417978
rect 579374 417922 579430 417978
rect 579498 417922 579554 417978
rect 579622 417922 579678 417978
rect 579250 400294 579306 400350
rect 579374 400294 579430 400350
rect 579498 400294 579554 400350
rect 579622 400294 579678 400350
rect 579250 400170 579306 400226
rect 579374 400170 579430 400226
rect 579498 400170 579554 400226
rect 579622 400170 579678 400226
rect 579250 400046 579306 400102
rect 579374 400046 579430 400102
rect 579498 400046 579554 400102
rect 579622 400046 579678 400102
rect 579250 399922 579306 399978
rect 579374 399922 579430 399978
rect 579498 399922 579554 399978
rect 579622 399922 579678 399978
rect 579250 382294 579306 382350
rect 579374 382294 579430 382350
rect 579498 382294 579554 382350
rect 579622 382294 579678 382350
rect 579250 382170 579306 382226
rect 579374 382170 579430 382226
rect 579498 382170 579554 382226
rect 579622 382170 579678 382226
rect 579250 382046 579306 382102
rect 579374 382046 579430 382102
rect 579498 382046 579554 382102
rect 579622 382046 579678 382102
rect 579250 381922 579306 381978
rect 579374 381922 579430 381978
rect 579498 381922 579554 381978
rect 579622 381922 579678 381978
rect 579250 364294 579306 364350
rect 579374 364294 579430 364350
rect 579498 364294 579554 364350
rect 579622 364294 579678 364350
rect 579250 364170 579306 364226
rect 579374 364170 579430 364226
rect 579498 364170 579554 364226
rect 579622 364170 579678 364226
rect 579250 364046 579306 364102
rect 579374 364046 579430 364102
rect 579498 364046 579554 364102
rect 579622 364046 579678 364102
rect 579250 363922 579306 363978
rect 579374 363922 579430 363978
rect 579498 363922 579554 363978
rect 579622 363922 579678 363978
rect 579250 346294 579306 346350
rect 579374 346294 579430 346350
rect 579498 346294 579554 346350
rect 579622 346294 579678 346350
rect 579250 346170 579306 346226
rect 579374 346170 579430 346226
rect 579498 346170 579554 346226
rect 579622 346170 579678 346226
rect 579250 346046 579306 346102
rect 579374 346046 579430 346102
rect 579498 346046 579554 346102
rect 579622 346046 579678 346102
rect 579250 345922 579306 345978
rect 579374 345922 579430 345978
rect 579498 345922 579554 345978
rect 579622 345922 579678 345978
rect 579250 328294 579306 328350
rect 579374 328294 579430 328350
rect 579498 328294 579554 328350
rect 579622 328294 579678 328350
rect 579250 328170 579306 328226
rect 579374 328170 579430 328226
rect 579498 328170 579554 328226
rect 579622 328170 579678 328226
rect 579250 328046 579306 328102
rect 579374 328046 579430 328102
rect 579498 328046 579554 328102
rect 579622 328046 579678 328102
rect 579250 327922 579306 327978
rect 579374 327922 579430 327978
rect 579498 327922 579554 327978
rect 579622 327922 579678 327978
rect 579250 310294 579306 310350
rect 579374 310294 579430 310350
rect 579498 310294 579554 310350
rect 579622 310294 579678 310350
rect 579250 310170 579306 310226
rect 579374 310170 579430 310226
rect 579498 310170 579554 310226
rect 579622 310170 579678 310226
rect 579250 310046 579306 310102
rect 579374 310046 579430 310102
rect 579498 310046 579554 310102
rect 579622 310046 579678 310102
rect 579250 309922 579306 309978
rect 579374 309922 579430 309978
rect 579498 309922 579554 309978
rect 579622 309922 579678 309978
rect 579250 292294 579306 292350
rect 579374 292294 579430 292350
rect 579498 292294 579554 292350
rect 579622 292294 579678 292350
rect 579250 292170 579306 292226
rect 579374 292170 579430 292226
rect 579498 292170 579554 292226
rect 579622 292170 579678 292226
rect 579250 292046 579306 292102
rect 579374 292046 579430 292102
rect 579498 292046 579554 292102
rect 579622 292046 579678 292102
rect 579250 291922 579306 291978
rect 579374 291922 579430 291978
rect 579498 291922 579554 291978
rect 579622 291922 579678 291978
rect 579250 274294 579306 274350
rect 579374 274294 579430 274350
rect 579498 274294 579554 274350
rect 579622 274294 579678 274350
rect 579250 274170 579306 274226
rect 579374 274170 579430 274226
rect 579498 274170 579554 274226
rect 579622 274170 579678 274226
rect 579250 274046 579306 274102
rect 579374 274046 579430 274102
rect 579498 274046 579554 274102
rect 579622 274046 579678 274102
rect 579250 273922 579306 273978
rect 579374 273922 579430 273978
rect 579498 273922 579554 273978
rect 579622 273922 579678 273978
rect 579250 256294 579306 256350
rect 579374 256294 579430 256350
rect 579498 256294 579554 256350
rect 579622 256294 579678 256350
rect 579250 256170 579306 256226
rect 579374 256170 579430 256226
rect 579498 256170 579554 256226
rect 579622 256170 579678 256226
rect 579250 256046 579306 256102
rect 579374 256046 579430 256102
rect 579498 256046 579554 256102
rect 579622 256046 579678 256102
rect 579250 255922 579306 255978
rect 579374 255922 579430 255978
rect 579498 255922 579554 255978
rect 579622 255922 579678 255978
rect 579250 238294 579306 238350
rect 579374 238294 579430 238350
rect 579498 238294 579554 238350
rect 579622 238294 579678 238350
rect 579250 238170 579306 238226
rect 579374 238170 579430 238226
rect 579498 238170 579554 238226
rect 579622 238170 579678 238226
rect 579250 238046 579306 238102
rect 579374 238046 579430 238102
rect 579498 238046 579554 238102
rect 579622 238046 579678 238102
rect 579250 237922 579306 237978
rect 579374 237922 579430 237978
rect 579498 237922 579554 237978
rect 579622 237922 579678 237978
rect 579250 220294 579306 220350
rect 579374 220294 579430 220350
rect 579498 220294 579554 220350
rect 579622 220294 579678 220350
rect 579250 220170 579306 220226
rect 579374 220170 579430 220226
rect 579498 220170 579554 220226
rect 579622 220170 579678 220226
rect 579250 220046 579306 220102
rect 579374 220046 579430 220102
rect 579498 220046 579554 220102
rect 579622 220046 579678 220102
rect 579250 219922 579306 219978
rect 579374 219922 579430 219978
rect 579498 219922 579554 219978
rect 579622 219922 579678 219978
rect 579250 202294 579306 202350
rect 579374 202294 579430 202350
rect 579498 202294 579554 202350
rect 579622 202294 579678 202350
rect 579250 202170 579306 202226
rect 579374 202170 579430 202226
rect 579498 202170 579554 202226
rect 579622 202170 579678 202226
rect 579250 202046 579306 202102
rect 579374 202046 579430 202102
rect 579498 202046 579554 202102
rect 579622 202046 579678 202102
rect 579250 201922 579306 201978
rect 579374 201922 579430 201978
rect 579498 201922 579554 201978
rect 579622 201922 579678 201978
rect 579250 184294 579306 184350
rect 579374 184294 579430 184350
rect 579498 184294 579554 184350
rect 579622 184294 579678 184350
rect 579250 184170 579306 184226
rect 579374 184170 579430 184226
rect 579498 184170 579554 184226
rect 579622 184170 579678 184226
rect 579250 184046 579306 184102
rect 579374 184046 579430 184102
rect 579498 184046 579554 184102
rect 579622 184046 579678 184102
rect 579250 183922 579306 183978
rect 579374 183922 579430 183978
rect 579498 183922 579554 183978
rect 579622 183922 579678 183978
rect 579250 166294 579306 166350
rect 579374 166294 579430 166350
rect 579498 166294 579554 166350
rect 579622 166294 579678 166350
rect 579250 166170 579306 166226
rect 579374 166170 579430 166226
rect 579498 166170 579554 166226
rect 579622 166170 579678 166226
rect 579250 166046 579306 166102
rect 579374 166046 579430 166102
rect 579498 166046 579554 166102
rect 579622 166046 579678 166102
rect 579250 165922 579306 165978
rect 579374 165922 579430 165978
rect 579498 165922 579554 165978
rect 579622 165922 579678 165978
rect 579250 148294 579306 148350
rect 579374 148294 579430 148350
rect 579498 148294 579554 148350
rect 579622 148294 579678 148350
rect 579250 148170 579306 148226
rect 579374 148170 579430 148226
rect 579498 148170 579554 148226
rect 579622 148170 579678 148226
rect 579250 148046 579306 148102
rect 579374 148046 579430 148102
rect 579498 148046 579554 148102
rect 579622 148046 579678 148102
rect 579250 147922 579306 147978
rect 579374 147922 579430 147978
rect 579498 147922 579554 147978
rect 579622 147922 579678 147978
rect 579250 130294 579306 130350
rect 579374 130294 579430 130350
rect 579498 130294 579554 130350
rect 579622 130294 579678 130350
rect 579250 130170 579306 130226
rect 579374 130170 579430 130226
rect 579498 130170 579554 130226
rect 579622 130170 579678 130226
rect 579250 130046 579306 130102
rect 579374 130046 579430 130102
rect 579498 130046 579554 130102
rect 579622 130046 579678 130102
rect 579250 129922 579306 129978
rect 579374 129922 579430 129978
rect 579498 129922 579554 129978
rect 579622 129922 579678 129978
rect 579250 112294 579306 112350
rect 579374 112294 579430 112350
rect 579498 112294 579554 112350
rect 579622 112294 579678 112350
rect 579250 112170 579306 112226
rect 579374 112170 579430 112226
rect 579498 112170 579554 112226
rect 579622 112170 579678 112226
rect 579250 112046 579306 112102
rect 579374 112046 579430 112102
rect 579498 112046 579554 112102
rect 579622 112046 579678 112102
rect 579250 111922 579306 111978
rect 579374 111922 579430 111978
rect 579498 111922 579554 111978
rect 579622 111922 579678 111978
rect 579250 94294 579306 94350
rect 579374 94294 579430 94350
rect 579498 94294 579554 94350
rect 579622 94294 579678 94350
rect 579250 94170 579306 94226
rect 579374 94170 579430 94226
rect 579498 94170 579554 94226
rect 579622 94170 579678 94226
rect 579250 94046 579306 94102
rect 579374 94046 579430 94102
rect 579498 94046 579554 94102
rect 579622 94046 579678 94102
rect 579250 93922 579306 93978
rect 579374 93922 579430 93978
rect 579498 93922 579554 93978
rect 579622 93922 579678 93978
rect 579250 76294 579306 76350
rect 579374 76294 579430 76350
rect 579498 76294 579554 76350
rect 579622 76294 579678 76350
rect 579250 76170 579306 76226
rect 579374 76170 579430 76226
rect 579498 76170 579554 76226
rect 579622 76170 579678 76226
rect 579250 76046 579306 76102
rect 579374 76046 579430 76102
rect 579498 76046 579554 76102
rect 579622 76046 579678 76102
rect 579250 75922 579306 75978
rect 579374 75922 579430 75978
rect 579498 75922 579554 75978
rect 579622 75922 579678 75978
rect 579250 58294 579306 58350
rect 579374 58294 579430 58350
rect 579498 58294 579554 58350
rect 579622 58294 579678 58350
rect 579250 58170 579306 58226
rect 579374 58170 579430 58226
rect 579498 58170 579554 58226
rect 579622 58170 579678 58226
rect 579250 58046 579306 58102
rect 579374 58046 579430 58102
rect 579498 58046 579554 58102
rect 579622 58046 579678 58102
rect 579250 57922 579306 57978
rect 579374 57922 579430 57978
rect 579498 57922 579554 57978
rect 579622 57922 579678 57978
rect 579250 40294 579306 40350
rect 579374 40294 579430 40350
rect 579498 40294 579554 40350
rect 579622 40294 579678 40350
rect 579250 40170 579306 40226
rect 579374 40170 579430 40226
rect 579498 40170 579554 40226
rect 579622 40170 579678 40226
rect 579250 40046 579306 40102
rect 579374 40046 579430 40102
rect 579498 40046 579554 40102
rect 579622 40046 579678 40102
rect 579250 39922 579306 39978
rect 579374 39922 579430 39978
rect 579498 39922 579554 39978
rect 579622 39922 579678 39978
rect 579250 22294 579306 22350
rect 579374 22294 579430 22350
rect 579498 22294 579554 22350
rect 579622 22294 579678 22350
rect 579250 22170 579306 22226
rect 579374 22170 579430 22226
rect 579498 22170 579554 22226
rect 579622 22170 579678 22226
rect 579250 22046 579306 22102
rect 579374 22046 579430 22102
rect 579498 22046 579554 22102
rect 579622 22046 579678 22102
rect 579250 21922 579306 21978
rect 579374 21922 579430 21978
rect 579498 21922 579554 21978
rect 579622 21922 579678 21978
rect 579250 4294 579306 4350
rect 579374 4294 579430 4350
rect 579498 4294 579554 4350
rect 579622 4294 579678 4350
rect 579250 4170 579306 4226
rect 579374 4170 579430 4226
rect 579498 4170 579554 4226
rect 579622 4170 579678 4226
rect 579250 4046 579306 4102
rect 579374 4046 579430 4102
rect 579498 4046 579554 4102
rect 579622 4046 579678 4102
rect 579250 3922 579306 3978
rect 579374 3922 579430 3978
rect 579498 3922 579554 3978
rect 579622 3922 579678 3978
rect 579250 -216 579306 -160
rect 579374 -216 579430 -160
rect 579498 -216 579554 -160
rect 579622 -216 579678 -160
rect 579250 -340 579306 -284
rect 579374 -340 579430 -284
rect 579498 -340 579554 -284
rect 579622 -340 579678 -284
rect 579250 -464 579306 -408
rect 579374 -464 579430 -408
rect 579498 -464 579554 -408
rect 579622 -464 579678 -408
rect 579250 -588 579306 -532
rect 579374 -588 579430 -532
rect 579498 -588 579554 -532
rect 579622 -588 579678 -532
rect 582970 598116 583026 598172
rect 583094 598116 583150 598172
rect 583218 598116 583274 598172
rect 583342 598116 583398 598172
rect 582970 597992 583026 598048
rect 583094 597992 583150 598048
rect 583218 597992 583274 598048
rect 583342 597992 583398 598048
rect 582970 597868 583026 597924
rect 583094 597868 583150 597924
rect 583218 597868 583274 597924
rect 583342 597868 583398 597924
rect 582970 597744 583026 597800
rect 583094 597744 583150 597800
rect 583218 597744 583274 597800
rect 583342 597744 583398 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 582970 586294 583026 586350
rect 583094 586294 583150 586350
rect 583218 586294 583274 586350
rect 583342 586294 583398 586350
rect 582970 586170 583026 586226
rect 583094 586170 583150 586226
rect 583218 586170 583274 586226
rect 583342 586170 583398 586226
rect 582970 586046 583026 586102
rect 583094 586046 583150 586102
rect 583218 586046 583274 586102
rect 583342 586046 583398 586102
rect 582970 585922 583026 585978
rect 583094 585922 583150 585978
rect 583218 585922 583274 585978
rect 583342 585922 583398 585978
rect 582970 568294 583026 568350
rect 583094 568294 583150 568350
rect 583218 568294 583274 568350
rect 583342 568294 583398 568350
rect 582970 568170 583026 568226
rect 583094 568170 583150 568226
rect 583218 568170 583274 568226
rect 583342 568170 583398 568226
rect 582970 568046 583026 568102
rect 583094 568046 583150 568102
rect 583218 568046 583274 568102
rect 583342 568046 583398 568102
rect 582970 567922 583026 567978
rect 583094 567922 583150 567978
rect 583218 567922 583274 567978
rect 583342 567922 583398 567978
rect 582970 550294 583026 550350
rect 583094 550294 583150 550350
rect 583218 550294 583274 550350
rect 583342 550294 583398 550350
rect 582970 550170 583026 550226
rect 583094 550170 583150 550226
rect 583218 550170 583274 550226
rect 583342 550170 583398 550226
rect 582970 550046 583026 550102
rect 583094 550046 583150 550102
rect 583218 550046 583274 550102
rect 583342 550046 583398 550102
rect 582970 549922 583026 549978
rect 583094 549922 583150 549978
rect 583218 549922 583274 549978
rect 583342 549922 583398 549978
rect 582970 532294 583026 532350
rect 583094 532294 583150 532350
rect 583218 532294 583274 532350
rect 583342 532294 583398 532350
rect 582970 532170 583026 532226
rect 583094 532170 583150 532226
rect 583218 532170 583274 532226
rect 583342 532170 583398 532226
rect 582970 532046 583026 532102
rect 583094 532046 583150 532102
rect 583218 532046 583274 532102
rect 583342 532046 583398 532102
rect 582970 531922 583026 531978
rect 583094 531922 583150 531978
rect 583218 531922 583274 531978
rect 583342 531922 583398 531978
rect 582970 514294 583026 514350
rect 583094 514294 583150 514350
rect 583218 514294 583274 514350
rect 583342 514294 583398 514350
rect 582970 514170 583026 514226
rect 583094 514170 583150 514226
rect 583218 514170 583274 514226
rect 583342 514170 583398 514226
rect 582970 514046 583026 514102
rect 583094 514046 583150 514102
rect 583218 514046 583274 514102
rect 583342 514046 583398 514102
rect 582970 513922 583026 513978
rect 583094 513922 583150 513978
rect 583218 513922 583274 513978
rect 583342 513922 583398 513978
rect 582970 496294 583026 496350
rect 583094 496294 583150 496350
rect 583218 496294 583274 496350
rect 583342 496294 583398 496350
rect 582970 496170 583026 496226
rect 583094 496170 583150 496226
rect 583218 496170 583274 496226
rect 583342 496170 583398 496226
rect 582970 496046 583026 496102
rect 583094 496046 583150 496102
rect 583218 496046 583274 496102
rect 583342 496046 583398 496102
rect 582970 495922 583026 495978
rect 583094 495922 583150 495978
rect 583218 495922 583274 495978
rect 583342 495922 583398 495978
rect 582970 478294 583026 478350
rect 583094 478294 583150 478350
rect 583218 478294 583274 478350
rect 583342 478294 583398 478350
rect 582970 478170 583026 478226
rect 583094 478170 583150 478226
rect 583218 478170 583274 478226
rect 583342 478170 583398 478226
rect 582970 478046 583026 478102
rect 583094 478046 583150 478102
rect 583218 478046 583274 478102
rect 583342 478046 583398 478102
rect 582970 477922 583026 477978
rect 583094 477922 583150 477978
rect 583218 477922 583274 477978
rect 583342 477922 583398 477978
rect 582970 460294 583026 460350
rect 583094 460294 583150 460350
rect 583218 460294 583274 460350
rect 583342 460294 583398 460350
rect 582970 460170 583026 460226
rect 583094 460170 583150 460226
rect 583218 460170 583274 460226
rect 583342 460170 583398 460226
rect 582970 460046 583026 460102
rect 583094 460046 583150 460102
rect 583218 460046 583274 460102
rect 583342 460046 583398 460102
rect 582970 459922 583026 459978
rect 583094 459922 583150 459978
rect 583218 459922 583274 459978
rect 583342 459922 583398 459978
rect 582970 442294 583026 442350
rect 583094 442294 583150 442350
rect 583218 442294 583274 442350
rect 583342 442294 583398 442350
rect 582970 442170 583026 442226
rect 583094 442170 583150 442226
rect 583218 442170 583274 442226
rect 583342 442170 583398 442226
rect 582970 442046 583026 442102
rect 583094 442046 583150 442102
rect 583218 442046 583274 442102
rect 583342 442046 583398 442102
rect 582970 441922 583026 441978
rect 583094 441922 583150 441978
rect 583218 441922 583274 441978
rect 583342 441922 583398 441978
rect 582970 424294 583026 424350
rect 583094 424294 583150 424350
rect 583218 424294 583274 424350
rect 583342 424294 583398 424350
rect 582970 424170 583026 424226
rect 583094 424170 583150 424226
rect 583218 424170 583274 424226
rect 583342 424170 583398 424226
rect 582970 424046 583026 424102
rect 583094 424046 583150 424102
rect 583218 424046 583274 424102
rect 583342 424046 583398 424102
rect 582970 423922 583026 423978
rect 583094 423922 583150 423978
rect 583218 423922 583274 423978
rect 583342 423922 583398 423978
rect 582970 406294 583026 406350
rect 583094 406294 583150 406350
rect 583218 406294 583274 406350
rect 583342 406294 583398 406350
rect 582970 406170 583026 406226
rect 583094 406170 583150 406226
rect 583218 406170 583274 406226
rect 583342 406170 583398 406226
rect 582970 406046 583026 406102
rect 583094 406046 583150 406102
rect 583218 406046 583274 406102
rect 583342 406046 583398 406102
rect 582970 405922 583026 405978
rect 583094 405922 583150 405978
rect 583218 405922 583274 405978
rect 583342 405922 583398 405978
rect 582970 388294 583026 388350
rect 583094 388294 583150 388350
rect 583218 388294 583274 388350
rect 583342 388294 583398 388350
rect 582970 388170 583026 388226
rect 583094 388170 583150 388226
rect 583218 388170 583274 388226
rect 583342 388170 583398 388226
rect 582970 388046 583026 388102
rect 583094 388046 583150 388102
rect 583218 388046 583274 388102
rect 583342 388046 583398 388102
rect 582970 387922 583026 387978
rect 583094 387922 583150 387978
rect 583218 387922 583274 387978
rect 583342 387922 583398 387978
rect 582970 370294 583026 370350
rect 583094 370294 583150 370350
rect 583218 370294 583274 370350
rect 583342 370294 583398 370350
rect 582970 370170 583026 370226
rect 583094 370170 583150 370226
rect 583218 370170 583274 370226
rect 583342 370170 583398 370226
rect 582970 370046 583026 370102
rect 583094 370046 583150 370102
rect 583218 370046 583274 370102
rect 583342 370046 583398 370102
rect 582970 369922 583026 369978
rect 583094 369922 583150 369978
rect 583218 369922 583274 369978
rect 583342 369922 583398 369978
rect 582970 352294 583026 352350
rect 583094 352294 583150 352350
rect 583218 352294 583274 352350
rect 583342 352294 583398 352350
rect 582970 352170 583026 352226
rect 583094 352170 583150 352226
rect 583218 352170 583274 352226
rect 583342 352170 583398 352226
rect 582970 352046 583026 352102
rect 583094 352046 583150 352102
rect 583218 352046 583274 352102
rect 583342 352046 583398 352102
rect 582970 351922 583026 351978
rect 583094 351922 583150 351978
rect 583218 351922 583274 351978
rect 583342 351922 583398 351978
rect 582970 334294 583026 334350
rect 583094 334294 583150 334350
rect 583218 334294 583274 334350
rect 583342 334294 583398 334350
rect 582970 334170 583026 334226
rect 583094 334170 583150 334226
rect 583218 334170 583274 334226
rect 583342 334170 583398 334226
rect 582970 334046 583026 334102
rect 583094 334046 583150 334102
rect 583218 334046 583274 334102
rect 583342 334046 583398 334102
rect 582970 333922 583026 333978
rect 583094 333922 583150 333978
rect 583218 333922 583274 333978
rect 583342 333922 583398 333978
rect 582970 316294 583026 316350
rect 583094 316294 583150 316350
rect 583218 316294 583274 316350
rect 583342 316294 583398 316350
rect 582970 316170 583026 316226
rect 583094 316170 583150 316226
rect 583218 316170 583274 316226
rect 583342 316170 583398 316226
rect 582970 316046 583026 316102
rect 583094 316046 583150 316102
rect 583218 316046 583274 316102
rect 583342 316046 583398 316102
rect 582970 315922 583026 315978
rect 583094 315922 583150 315978
rect 583218 315922 583274 315978
rect 583342 315922 583398 315978
rect 582970 298294 583026 298350
rect 583094 298294 583150 298350
rect 583218 298294 583274 298350
rect 583342 298294 583398 298350
rect 582970 298170 583026 298226
rect 583094 298170 583150 298226
rect 583218 298170 583274 298226
rect 583342 298170 583398 298226
rect 582970 298046 583026 298102
rect 583094 298046 583150 298102
rect 583218 298046 583274 298102
rect 583342 298046 583398 298102
rect 582970 297922 583026 297978
rect 583094 297922 583150 297978
rect 583218 297922 583274 297978
rect 583342 297922 583398 297978
rect 582970 280294 583026 280350
rect 583094 280294 583150 280350
rect 583218 280294 583274 280350
rect 583342 280294 583398 280350
rect 582970 280170 583026 280226
rect 583094 280170 583150 280226
rect 583218 280170 583274 280226
rect 583342 280170 583398 280226
rect 582970 280046 583026 280102
rect 583094 280046 583150 280102
rect 583218 280046 583274 280102
rect 583342 280046 583398 280102
rect 582970 279922 583026 279978
rect 583094 279922 583150 279978
rect 583218 279922 583274 279978
rect 583342 279922 583398 279978
rect 582970 262294 583026 262350
rect 583094 262294 583150 262350
rect 583218 262294 583274 262350
rect 583342 262294 583398 262350
rect 582970 262170 583026 262226
rect 583094 262170 583150 262226
rect 583218 262170 583274 262226
rect 583342 262170 583398 262226
rect 582970 262046 583026 262102
rect 583094 262046 583150 262102
rect 583218 262046 583274 262102
rect 583342 262046 583398 262102
rect 582970 261922 583026 261978
rect 583094 261922 583150 261978
rect 583218 261922 583274 261978
rect 583342 261922 583398 261978
rect 582970 244294 583026 244350
rect 583094 244294 583150 244350
rect 583218 244294 583274 244350
rect 583342 244294 583398 244350
rect 582970 244170 583026 244226
rect 583094 244170 583150 244226
rect 583218 244170 583274 244226
rect 583342 244170 583398 244226
rect 582970 244046 583026 244102
rect 583094 244046 583150 244102
rect 583218 244046 583274 244102
rect 583342 244046 583398 244102
rect 582970 243922 583026 243978
rect 583094 243922 583150 243978
rect 583218 243922 583274 243978
rect 583342 243922 583398 243978
rect 582970 226294 583026 226350
rect 583094 226294 583150 226350
rect 583218 226294 583274 226350
rect 583342 226294 583398 226350
rect 582970 226170 583026 226226
rect 583094 226170 583150 226226
rect 583218 226170 583274 226226
rect 583342 226170 583398 226226
rect 582970 226046 583026 226102
rect 583094 226046 583150 226102
rect 583218 226046 583274 226102
rect 583342 226046 583398 226102
rect 582970 225922 583026 225978
rect 583094 225922 583150 225978
rect 583218 225922 583274 225978
rect 583342 225922 583398 225978
rect 582970 208294 583026 208350
rect 583094 208294 583150 208350
rect 583218 208294 583274 208350
rect 583342 208294 583398 208350
rect 582970 208170 583026 208226
rect 583094 208170 583150 208226
rect 583218 208170 583274 208226
rect 583342 208170 583398 208226
rect 582970 208046 583026 208102
rect 583094 208046 583150 208102
rect 583218 208046 583274 208102
rect 583342 208046 583398 208102
rect 582970 207922 583026 207978
rect 583094 207922 583150 207978
rect 583218 207922 583274 207978
rect 583342 207922 583398 207978
rect 582970 190294 583026 190350
rect 583094 190294 583150 190350
rect 583218 190294 583274 190350
rect 583342 190294 583398 190350
rect 582970 190170 583026 190226
rect 583094 190170 583150 190226
rect 583218 190170 583274 190226
rect 583342 190170 583398 190226
rect 582970 190046 583026 190102
rect 583094 190046 583150 190102
rect 583218 190046 583274 190102
rect 583342 190046 583398 190102
rect 582970 189922 583026 189978
rect 583094 189922 583150 189978
rect 583218 189922 583274 189978
rect 583342 189922 583398 189978
rect 582970 172294 583026 172350
rect 583094 172294 583150 172350
rect 583218 172294 583274 172350
rect 583342 172294 583398 172350
rect 582970 172170 583026 172226
rect 583094 172170 583150 172226
rect 583218 172170 583274 172226
rect 583342 172170 583398 172226
rect 582970 172046 583026 172102
rect 583094 172046 583150 172102
rect 583218 172046 583274 172102
rect 583342 172046 583398 172102
rect 582970 171922 583026 171978
rect 583094 171922 583150 171978
rect 583218 171922 583274 171978
rect 583342 171922 583398 171978
rect 582970 154294 583026 154350
rect 583094 154294 583150 154350
rect 583218 154294 583274 154350
rect 583342 154294 583398 154350
rect 582970 154170 583026 154226
rect 583094 154170 583150 154226
rect 583218 154170 583274 154226
rect 583342 154170 583398 154226
rect 582970 154046 583026 154102
rect 583094 154046 583150 154102
rect 583218 154046 583274 154102
rect 583342 154046 583398 154102
rect 582970 153922 583026 153978
rect 583094 153922 583150 153978
rect 583218 153922 583274 153978
rect 583342 153922 583398 153978
rect 582970 136294 583026 136350
rect 583094 136294 583150 136350
rect 583218 136294 583274 136350
rect 583342 136294 583398 136350
rect 582970 136170 583026 136226
rect 583094 136170 583150 136226
rect 583218 136170 583274 136226
rect 583342 136170 583398 136226
rect 582970 136046 583026 136102
rect 583094 136046 583150 136102
rect 583218 136046 583274 136102
rect 583342 136046 583398 136102
rect 582970 135922 583026 135978
rect 583094 135922 583150 135978
rect 583218 135922 583274 135978
rect 583342 135922 583398 135978
rect 582970 118294 583026 118350
rect 583094 118294 583150 118350
rect 583218 118294 583274 118350
rect 583342 118294 583398 118350
rect 582970 118170 583026 118226
rect 583094 118170 583150 118226
rect 583218 118170 583274 118226
rect 583342 118170 583398 118226
rect 582970 118046 583026 118102
rect 583094 118046 583150 118102
rect 583218 118046 583274 118102
rect 583342 118046 583398 118102
rect 582970 117922 583026 117978
rect 583094 117922 583150 117978
rect 583218 117922 583274 117978
rect 583342 117922 583398 117978
rect 582970 100294 583026 100350
rect 583094 100294 583150 100350
rect 583218 100294 583274 100350
rect 583342 100294 583398 100350
rect 582970 100170 583026 100226
rect 583094 100170 583150 100226
rect 583218 100170 583274 100226
rect 583342 100170 583398 100226
rect 582970 100046 583026 100102
rect 583094 100046 583150 100102
rect 583218 100046 583274 100102
rect 583342 100046 583398 100102
rect 582970 99922 583026 99978
rect 583094 99922 583150 99978
rect 583218 99922 583274 99978
rect 583342 99922 583398 99978
rect 582970 82294 583026 82350
rect 583094 82294 583150 82350
rect 583218 82294 583274 82350
rect 583342 82294 583398 82350
rect 582970 82170 583026 82226
rect 583094 82170 583150 82226
rect 583218 82170 583274 82226
rect 583342 82170 583398 82226
rect 582970 82046 583026 82102
rect 583094 82046 583150 82102
rect 583218 82046 583274 82102
rect 583342 82046 583398 82102
rect 582970 81922 583026 81978
rect 583094 81922 583150 81978
rect 583218 81922 583274 81978
rect 583342 81922 583398 81978
rect 582970 64294 583026 64350
rect 583094 64294 583150 64350
rect 583218 64294 583274 64350
rect 583342 64294 583398 64350
rect 582970 64170 583026 64226
rect 583094 64170 583150 64226
rect 583218 64170 583274 64226
rect 583342 64170 583398 64226
rect 582970 64046 583026 64102
rect 583094 64046 583150 64102
rect 583218 64046 583274 64102
rect 583342 64046 583398 64102
rect 582970 63922 583026 63978
rect 583094 63922 583150 63978
rect 583218 63922 583274 63978
rect 583342 63922 583398 63978
rect 582970 46294 583026 46350
rect 583094 46294 583150 46350
rect 583218 46294 583274 46350
rect 583342 46294 583398 46350
rect 582970 46170 583026 46226
rect 583094 46170 583150 46226
rect 583218 46170 583274 46226
rect 583342 46170 583398 46226
rect 582970 46046 583026 46102
rect 583094 46046 583150 46102
rect 583218 46046 583274 46102
rect 583342 46046 583398 46102
rect 582970 45922 583026 45978
rect 583094 45922 583150 45978
rect 583218 45922 583274 45978
rect 583342 45922 583398 45978
rect 582970 28294 583026 28350
rect 583094 28294 583150 28350
rect 583218 28294 583274 28350
rect 583342 28294 583398 28350
rect 582970 28170 583026 28226
rect 583094 28170 583150 28226
rect 583218 28170 583274 28226
rect 583342 28170 583398 28226
rect 582970 28046 583026 28102
rect 583094 28046 583150 28102
rect 583218 28046 583274 28102
rect 583342 28046 583398 28102
rect 582970 27922 583026 27978
rect 583094 27922 583150 27978
rect 583218 27922 583274 27978
rect 583342 27922 583398 27978
rect 582970 10294 583026 10350
rect 583094 10294 583150 10350
rect 583218 10294 583274 10350
rect 583342 10294 583398 10350
rect 582970 10170 583026 10226
rect 583094 10170 583150 10226
rect 583218 10170 583274 10226
rect 583342 10170 583398 10226
rect 582970 10046 583026 10102
rect 583094 10046 583150 10102
rect 583218 10046 583274 10102
rect 583342 10046 583398 10102
rect 582970 9922 583026 9978
rect 583094 9922 583150 9978
rect 583218 9922 583274 9978
rect 583342 9922 583398 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 582970 -1176 583026 -1120
rect 583094 -1176 583150 -1120
rect 583218 -1176 583274 -1120
rect 583342 -1176 583398 -1120
rect 582970 -1300 583026 -1244
rect 583094 -1300 583150 -1244
rect 583218 -1300 583274 -1244
rect 583342 -1300 583398 -1244
rect 582970 -1424 583026 -1368
rect 583094 -1424 583150 -1368
rect 583218 -1424 583274 -1368
rect 583342 -1424 583398 -1368
rect 582970 -1548 583026 -1492
rect 583094 -1548 583150 -1492
rect 583218 -1548 583274 -1492
rect 583342 -1548 583398 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 6970 598172
rect 7026 598116 7094 598172
rect 7150 598116 7218 598172
rect 7274 598116 7342 598172
rect 7398 598116 24970 598172
rect 25026 598116 25094 598172
rect 25150 598116 25218 598172
rect 25274 598116 25342 598172
rect 25398 598116 42970 598172
rect 43026 598116 43094 598172
rect 43150 598116 43218 598172
rect 43274 598116 43342 598172
rect 43398 598116 60970 598172
rect 61026 598116 61094 598172
rect 61150 598116 61218 598172
rect 61274 598116 61342 598172
rect 61398 598116 78970 598172
rect 79026 598116 79094 598172
rect 79150 598116 79218 598172
rect 79274 598116 79342 598172
rect 79398 598116 96970 598172
rect 97026 598116 97094 598172
rect 97150 598116 97218 598172
rect 97274 598116 97342 598172
rect 97398 598116 114970 598172
rect 115026 598116 115094 598172
rect 115150 598116 115218 598172
rect 115274 598116 115342 598172
rect 115398 598116 132970 598172
rect 133026 598116 133094 598172
rect 133150 598116 133218 598172
rect 133274 598116 133342 598172
rect 133398 598116 150970 598172
rect 151026 598116 151094 598172
rect 151150 598116 151218 598172
rect 151274 598116 151342 598172
rect 151398 598116 168970 598172
rect 169026 598116 169094 598172
rect 169150 598116 169218 598172
rect 169274 598116 169342 598172
rect 169398 598116 186970 598172
rect 187026 598116 187094 598172
rect 187150 598116 187218 598172
rect 187274 598116 187342 598172
rect 187398 598116 204970 598172
rect 205026 598116 205094 598172
rect 205150 598116 205218 598172
rect 205274 598116 205342 598172
rect 205398 598116 222970 598172
rect 223026 598116 223094 598172
rect 223150 598116 223218 598172
rect 223274 598116 223342 598172
rect 223398 598116 240970 598172
rect 241026 598116 241094 598172
rect 241150 598116 241218 598172
rect 241274 598116 241342 598172
rect 241398 598116 258970 598172
rect 259026 598116 259094 598172
rect 259150 598116 259218 598172
rect 259274 598116 259342 598172
rect 259398 598116 276970 598172
rect 277026 598116 277094 598172
rect 277150 598116 277218 598172
rect 277274 598116 277342 598172
rect 277398 598116 294970 598172
rect 295026 598116 295094 598172
rect 295150 598116 295218 598172
rect 295274 598116 295342 598172
rect 295398 598116 312970 598172
rect 313026 598116 313094 598172
rect 313150 598116 313218 598172
rect 313274 598116 313342 598172
rect 313398 598116 330970 598172
rect 331026 598116 331094 598172
rect 331150 598116 331218 598172
rect 331274 598116 331342 598172
rect 331398 598116 348970 598172
rect 349026 598116 349094 598172
rect 349150 598116 349218 598172
rect 349274 598116 349342 598172
rect 349398 598116 366970 598172
rect 367026 598116 367094 598172
rect 367150 598116 367218 598172
rect 367274 598116 367342 598172
rect 367398 598116 384970 598172
rect 385026 598116 385094 598172
rect 385150 598116 385218 598172
rect 385274 598116 385342 598172
rect 385398 598116 402970 598172
rect 403026 598116 403094 598172
rect 403150 598116 403218 598172
rect 403274 598116 403342 598172
rect 403398 598116 420970 598172
rect 421026 598116 421094 598172
rect 421150 598116 421218 598172
rect 421274 598116 421342 598172
rect 421398 598116 438970 598172
rect 439026 598116 439094 598172
rect 439150 598116 439218 598172
rect 439274 598116 439342 598172
rect 439398 598116 456970 598172
rect 457026 598116 457094 598172
rect 457150 598116 457218 598172
rect 457274 598116 457342 598172
rect 457398 598116 474970 598172
rect 475026 598116 475094 598172
rect 475150 598116 475218 598172
rect 475274 598116 475342 598172
rect 475398 598116 492970 598172
rect 493026 598116 493094 598172
rect 493150 598116 493218 598172
rect 493274 598116 493342 598172
rect 493398 598116 510970 598172
rect 511026 598116 511094 598172
rect 511150 598116 511218 598172
rect 511274 598116 511342 598172
rect 511398 598116 528970 598172
rect 529026 598116 529094 598172
rect 529150 598116 529218 598172
rect 529274 598116 529342 598172
rect 529398 598116 546970 598172
rect 547026 598116 547094 598172
rect 547150 598116 547218 598172
rect 547274 598116 547342 598172
rect 547398 598116 564970 598172
rect 565026 598116 565094 598172
rect 565150 598116 565218 598172
rect 565274 598116 565342 598172
rect 565398 598116 582970 598172
rect 583026 598116 583094 598172
rect 583150 598116 583218 598172
rect 583274 598116 583342 598172
rect 583398 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 6970 598048
rect 7026 597992 7094 598048
rect 7150 597992 7218 598048
rect 7274 597992 7342 598048
rect 7398 597992 24970 598048
rect 25026 597992 25094 598048
rect 25150 597992 25218 598048
rect 25274 597992 25342 598048
rect 25398 597992 42970 598048
rect 43026 597992 43094 598048
rect 43150 597992 43218 598048
rect 43274 597992 43342 598048
rect 43398 597992 60970 598048
rect 61026 597992 61094 598048
rect 61150 597992 61218 598048
rect 61274 597992 61342 598048
rect 61398 597992 78970 598048
rect 79026 597992 79094 598048
rect 79150 597992 79218 598048
rect 79274 597992 79342 598048
rect 79398 597992 96970 598048
rect 97026 597992 97094 598048
rect 97150 597992 97218 598048
rect 97274 597992 97342 598048
rect 97398 597992 114970 598048
rect 115026 597992 115094 598048
rect 115150 597992 115218 598048
rect 115274 597992 115342 598048
rect 115398 597992 132970 598048
rect 133026 597992 133094 598048
rect 133150 597992 133218 598048
rect 133274 597992 133342 598048
rect 133398 597992 150970 598048
rect 151026 597992 151094 598048
rect 151150 597992 151218 598048
rect 151274 597992 151342 598048
rect 151398 597992 168970 598048
rect 169026 597992 169094 598048
rect 169150 597992 169218 598048
rect 169274 597992 169342 598048
rect 169398 597992 186970 598048
rect 187026 597992 187094 598048
rect 187150 597992 187218 598048
rect 187274 597992 187342 598048
rect 187398 597992 204970 598048
rect 205026 597992 205094 598048
rect 205150 597992 205218 598048
rect 205274 597992 205342 598048
rect 205398 597992 222970 598048
rect 223026 597992 223094 598048
rect 223150 597992 223218 598048
rect 223274 597992 223342 598048
rect 223398 597992 240970 598048
rect 241026 597992 241094 598048
rect 241150 597992 241218 598048
rect 241274 597992 241342 598048
rect 241398 597992 258970 598048
rect 259026 597992 259094 598048
rect 259150 597992 259218 598048
rect 259274 597992 259342 598048
rect 259398 597992 276970 598048
rect 277026 597992 277094 598048
rect 277150 597992 277218 598048
rect 277274 597992 277342 598048
rect 277398 597992 294970 598048
rect 295026 597992 295094 598048
rect 295150 597992 295218 598048
rect 295274 597992 295342 598048
rect 295398 597992 312970 598048
rect 313026 597992 313094 598048
rect 313150 597992 313218 598048
rect 313274 597992 313342 598048
rect 313398 597992 330970 598048
rect 331026 597992 331094 598048
rect 331150 597992 331218 598048
rect 331274 597992 331342 598048
rect 331398 597992 348970 598048
rect 349026 597992 349094 598048
rect 349150 597992 349218 598048
rect 349274 597992 349342 598048
rect 349398 597992 366970 598048
rect 367026 597992 367094 598048
rect 367150 597992 367218 598048
rect 367274 597992 367342 598048
rect 367398 597992 384970 598048
rect 385026 597992 385094 598048
rect 385150 597992 385218 598048
rect 385274 597992 385342 598048
rect 385398 597992 402970 598048
rect 403026 597992 403094 598048
rect 403150 597992 403218 598048
rect 403274 597992 403342 598048
rect 403398 597992 420970 598048
rect 421026 597992 421094 598048
rect 421150 597992 421218 598048
rect 421274 597992 421342 598048
rect 421398 597992 438970 598048
rect 439026 597992 439094 598048
rect 439150 597992 439218 598048
rect 439274 597992 439342 598048
rect 439398 597992 456970 598048
rect 457026 597992 457094 598048
rect 457150 597992 457218 598048
rect 457274 597992 457342 598048
rect 457398 597992 474970 598048
rect 475026 597992 475094 598048
rect 475150 597992 475218 598048
rect 475274 597992 475342 598048
rect 475398 597992 492970 598048
rect 493026 597992 493094 598048
rect 493150 597992 493218 598048
rect 493274 597992 493342 598048
rect 493398 597992 510970 598048
rect 511026 597992 511094 598048
rect 511150 597992 511218 598048
rect 511274 597992 511342 598048
rect 511398 597992 528970 598048
rect 529026 597992 529094 598048
rect 529150 597992 529218 598048
rect 529274 597992 529342 598048
rect 529398 597992 546970 598048
rect 547026 597992 547094 598048
rect 547150 597992 547218 598048
rect 547274 597992 547342 598048
rect 547398 597992 564970 598048
rect 565026 597992 565094 598048
rect 565150 597992 565218 598048
rect 565274 597992 565342 598048
rect 565398 597992 582970 598048
rect 583026 597992 583094 598048
rect 583150 597992 583218 598048
rect 583274 597992 583342 598048
rect 583398 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 6970 597924
rect 7026 597868 7094 597924
rect 7150 597868 7218 597924
rect 7274 597868 7342 597924
rect 7398 597868 24970 597924
rect 25026 597868 25094 597924
rect 25150 597868 25218 597924
rect 25274 597868 25342 597924
rect 25398 597868 42970 597924
rect 43026 597868 43094 597924
rect 43150 597868 43218 597924
rect 43274 597868 43342 597924
rect 43398 597868 60970 597924
rect 61026 597868 61094 597924
rect 61150 597868 61218 597924
rect 61274 597868 61342 597924
rect 61398 597868 78970 597924
rect 79026 597868 79094 597924
rect 79150 597868 79218 597924
rect 79274 597868 79342 597924
rect 79398 597868 96970 597924
rect 97026 597868 97094 597924
rect 97150 597868 97218 597924
rect 97274 597868 97342 597924
rect 97398 597868 114970 597924
rect 115026 597868 115094 597924
rect 115150 597868 115218 597924
rect 115274 597868 115342 597924
rect 115398 597868 132970 597924
rect 133026 597868 133094 597924
rect 133150 597868 133218 597924
rect 133274 597868 133342 597924
rect 133398 597868 150970 597924
rect 151026 597868 151094 597924
rect 151150 597868 151218 597924
rect 151274 597868 151342 597924
rect 151398 597868 168970 597924
rect 169026 597868 169094 597924
rect 169150 597868 169218 597924
rect 169274 597868 169342 597924
rect 169398 597868 186970 597924
rect 187026 597868 187094 597924
rect 187150 597868 187218 597924
rect 187274 597868 187342 597924
rect 187398 597868 204970 597924
rect 205026 597868 205094 597924
rect 205150 597868 205218 597924
rect 205274 597868 205342 597924
rect 205398 597868 222970 597924
rect 223026 597868 223094 597924
rect 223150 597868 223218 597924
rect 223274 597868 223342 597924
rect 223398 597868 240970 597924
rect 241026 597868 241094 597924
rect 241150 597868 241218 597924
rect 241274 597868 241342 597924
rect 241398 597868 258970 597924
rect 259026 597868 259094 597924
rect 259150 597868 259218 597924
rect 259274 597868 259342 597924
rect 259398 597868 276970 597924
rect 277026 597868 277094 597924
rect 277150 597868 277218 597924
rect 277274 597868 277342 597924
rect 277398 597868 294970 597924
rect 295026 597868 295094 597924
rect 295150 597868 295218 597924
rect 295274 597868 295342 597924
rect 295398 597868 312970 597924
rect 313026 597868 313094 597924
rect 313150 597868 313218 597924
rect 313274 597868 313342 597924
rect 313398 597868 330970 597924
rect 331026 597868 331094 597924
rect 331150 597868 331218 597924
rect 331274 597868 331342 597924
rect 331398 597868 348970 597924
rect 349026 597868 349094 597924
rect 349150 597868 349218 597924
rect 349274 597868 349342 597924
rect 349398 597868 366970 597924
rect 367026 597868 367094 597924
rect 367150 597868 367218 597924
rect 367274 597868 367342 597924
rect 367398 597868 384970 597924
rect 385026 597868 385094 597924
rect 385150 597868 385218 597924
rect 385274 597868 385342 597924
rect 385398 597868 402970 597924
rect 403026 597868 403094 597924
rect 403150 597868 403218 597924
rect 403274 597868 403342 597924
rect 403398 597868 420970 597924
rect 421026 597868 421094 597924
rect 421150 597868 421218 597924
rect 421274 597868 421342 597924
rect 421398 597868 438970 597924
rect 439026 597868 439094 597924
rect 439150 597868 439218 597924
rect 439274 597868 439342 597924
rect 439398 597868 456970 597924
rect 457026 597868 457094 597924
rect 457150 597868 457218 597924
rect 457274 597868 457342 597924
rect 457398 597868 474970 597924
rect 475026 597868 475094 597924
rect 475150 597868 475218 597924
rect 475274 597868 475342 597924
rect 475398 597868 492970 597924
rect 493026 597868 493094 597924
rect 493150 597868 493218 597924
rect 493274 597868 493342 597924
rect 493398 597868 510970 597924
rect 511026 597868 511094 597924
rect 511150 597868 511218 597924
rect 511274 597868 511342 597924
rect 511398 597868 528970 597924
rect 529026 597868 529094 597924
rect 529150 597868 529218 597924
rect 529274 597868 529342 597924
rect 529398 597868 546970 597924
rect 547026 597868 547094 597924
rect 547150 597868 547218 597924
rect 547274 597868 547342 597924
rect 547398 597868 564970 597924
rect 565026 597868 565094 597924
rect 565150 597868 565218 597924
rect 565274 597868 565342 597924
rect 565398 597868 582970 597924
rect 583026 597868 583094 597924
rect 583150 597868 583218 597924
rect 583274 597868 583342 597924
rect 583398 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 6970 597800
rect 7026 597744 7094 597800
rect 7150 597744 7218 597800
rect 7274 597744 7342 597800
rect 7398 597744 24970 597800
rect 25026 597744 25094 597800
rect 25150 597744 25218 597800
rect 25274 597744 25342 597800
rect 25398 597744 42970 597800
rect 43026 597744 43094 597800
rect 43150 597744 43218 597800
rect 43274 597744 43342 597800
rect 43398 597744 60970 597800
rect 61026 597744 61094 597800
rect 61150 597744 61218 597800
rect 61274 597744 61342 597800
rect 61398 597744 78970 597800
rect 79026 597744 79094 597800
rect 79150 597744 79218 597800
rect 79274 597744 79342 597800
rect 79398 597744 96970 597800
rect 97026 597744 97094 597800
rect 97150 597744 97218 597800
rect 97274 597744 97342 597800
rect 97398 597744 114970 597800
rect 115026 597744 115094 597800
rect 115150 597744 115218 597800
rect 115274 597744 115342 597800
rect 115398 597744 132970 597800
rect 133026 597744 133094 597800
rect 133150 597744 133218 597800
rect 133274 597744 133342 597800
rect 133398 597744 150970 597800
rect 151026 597744 151094 597800
rect 151150 597744 151218 597800
rect 151274 597744 151342 597800
rect 151398 597744 168970 597800
rect 169026 597744 169094 597800
rect 169150 597744 169218 597800
rect 169274 597744 169342 597800
rect 169398 597744 186970 597800
rect 187026 597744 187094 597800
rect 187150 597744 187218 597800
rect 187274 597744 187342 597800
rect 187398 597744 204970 597800
rect 205026 597744 205094 597800
rect 205150 597744 205218 597800
rect 205274 597744 205342 597800
rect 205398 597744 222970 597800
rect 223026 597744 223094 597800
rect 223150 597744 223218 597800
rect 223274 597744 223342 597800
rect 223398 597744 240970 597800
rect 241026 597744 241094 597800
rect 241150 597744 241218 597800
rect 241274 597744 241342 597800
rect 241398 597744 258970 597800
rect 259026 597744 259094 597800
rect 259150 597744 259218 597800
rect 259274 597744 259342 597800
rect 259398 597744 276970 597800
rect 277026 597744 277094 597800
rect 277150 597744 277218 597800
rect 277274 597744 277342 597800
rect 277398 597744 294970 597800
rect 295026 597744 295094 597800
rect 295150 597744 295218 597800
rect 295274 597744 295342 597800
rect 295398 597744 312970 597800
rect 313026 597744 313094 597800
rect 313150 597744 313218 597800
rect 313274 597744 313342 597800
rect 313398 597744 330970 597800
rect 331026 597744 331094 597800
rect 331150 597744 331218 597800
rect 331274 597744 331342 597800
rect 331398 597744 348970 597800
rect 349026 597744 349094 597800
rect 349150 597744 349218 597800
rect 349274 597744 349342 597800
rect 349398 597744 366970 597800
rect 367026 597744 367094 597800
rect 367150 597744 367218 597800
rect 367274 597744 367342 597800
rect 367398 597744 384970 597800
rect 385026 597744 385094 597800
rect 385150 597744 385218 597800
rect 385274 597744 385342 597800
rect 385398 597744 402970 597800
rect 403026 597744 403094 597800
rect 403150 597744 403218 597800
rect 403274 597744 403342 597800
rect 403398 597744 420970 597800
rect 421026 597744 421094 597800
rect 421150 597744 421218 597800
rect 421274 597744 421342 597800
rect 421398 597744 438970 597800
rect 439026 597744 439094 597800
rect 439150 597744 439218 597800
rect 439274 597744 439342 597800
rect 439398 597744 456970 597800
rect 457026 597744 457094 597800
rect 457150 597744 457218 597800
rect 457274 597744 457342 597800
rect 457398 597744 474970 597800
rect 475026 597744 475094 597800
rect 475150 597744 475218 597800
rect 475274 597744 475342 597800
rect 475398 597744 492970 597800
rect 493026 597744 493094 597800
rect 493150 597744 493218 597800
rect 493274 597744 493342 597800
rect 493398 597744 510970 597800
rect 511026 597744 511094 597800
rect 511150 597744 511218 597800
rect 511274 597744 511342 597800
rect 511398 597744 528970 597800
rect 529026 597744 529094 597800
rect 529150 597744 529218 597800
rect 529274 597744 529342 597800
rect 529398 597744 546970 597800
rect 547026 597744 547094 597800
rect 547150 597744 547218 597800
rect 547274 597744 547342 597800
rect 547398 597744 564970 597800
rect 565026 597744 565094 597800
rect 565150 597744 565218 597800
rect 565274 597744 565342 597800
rect 565398 597744 582970 597800
rect 583026 597744 583094 597800
rect 583150 597744 583218 597800
rect 583274 597744 583342 597800
rect 583398 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 3250 597212
rect 3306 597156 3374 597212
rect 3430 597156 3498 597212
rect 3554 597156 3622 597212
rect 3678 597156 21250 597212
rect 21306 597156 21374 597212
rect 21430 597156 21498 597212
rect 21554 597156 21622 597212
rect 21678 597156 39250 597212
rect 39306 597156 39374 597212
rect 39430 597156 39498 597212
rect 39554 597156 39622 597212
rect 39678 597156 57250 597212
rect 57306 597156 57374 597212
rect 57430 597156 57498 597212
rect 57554 597156 57622 597212
rect 57678 597156 75250 597212
rect 75306 597156 75374 597212
rect 75430 597156 75498 597212
rect 75554 597156 75622 597212
rect 75678 597156 93250 597212
rect 93306 597156 93374 597212
rect 93430 597156 93498 597212
rect 93554 597156 93622 597212
rect 93678 597156 111250 597212
rect 111306 597156 111374 597212
rect 111430 597156 111498 597212
rect 111554 597156 111622 597212
rect 111678 597156 129250 597212
rect 129306 597156 129374 597212
rect 129430 597156 129498 597212
rect 129554 597156 129622 597212
rect 129678 597156 147250 597212
rect 147306 597156 147374 597212
rect 147430 597156 147498 597212
rect 147554 597156 147622 597212
rect 147678 597156 165250 597212
rect 165306 597156 165374 597212
rect 165430 597156 165498 597212
rect 165554 597156 165622 597212
rect 165678 597156 183250 597212
rect 183306 597156 183374 597212
rect 183430 597156 183498 597212
rect 183554 597156 183622 597212
rect 183678 597156 201250 597212
rect 201306 597156 201374 597212
rect 201430 597156 201498 597212
rect 201554 597156 201622 597212
rect 201678 597156 219250 597212
rect 219306 597156 219374 597212
rect 219430 597156 219498 597212
rect 219554 597156 219622 597212
rect 219678 597156 237250 597212
rect 237306 597156 237374 597212
rect 237430 597156 237498 597212
rect 237554 597156 237622 597212
rect 237678 597156 255250 597212
rect 255306 597156 255374 597212
rect 255430 597156 255498 597212
rect 255554 597156 255622 597212
rect 255678 597156 273250 597212
rect 273306 597156 273374 597212
rect 273430 597156 273498 597212
rect 273554 597156 273622 597212
rect 273678 597156 291250 597212
rect 291306 597156 291374 597212
rect 291430 597156 291498 597212
rect 291554 597156 291622 597212
rect 291678 597156 309250 597212
rect 309306 597156 309374 597212
rect 309430 597156 309498 597212
rect 309554 597156 309622 597212
rect 309678 597156 327250 597212
rect 327306 597156 327374 597212
rect 327430 597156 327498 597212
rect 327554 597156 327622 597212
rect 327678 597156 345250 597212
rect 345306 597156 345374 597212
rect 345430 597156 345498 597212
rect 345554 597156 345622 597212
rect 345678 597156 363250 597212
rect 363306 597156 363374 597212
rect 363430 597156 363498 597212
rect 363554 597156 363622 597212
rect 363678 597156 381250 597212
rect 381306 597156 381374 597212
rect 381430 597156 381498 597212
rect 381554 597156 381622 597212
rect 381678 597156 399250 597212
rect 399306 597156 399374 597212
rect 399430 597156 399498 597212
rect 399554 597156 399622 597212
rect 399678 597156 417250 597212
rect 417306 597156 417374 597212
rect 417430 597156 417498 597212
rect 417554 597156 417622 597212
rect 417678 597156 435250 597212
rect 435306 597156 435374 597212
rect 435430 597156 435498 597212
rect 435554 597156 435622 597212
rect 435678 597156 453250 597212
rect 453306 597156 453374 597212
rect 453430 597156 453498 597212
rect 453554 597156 453622 597212
rect 453678 597156 471250 597212
rect 471306 597156 471374 597212
rect 471430 597156 471498 597212
rect 471554 597156 471622 597212
rect 471678 597156 489250 597212
rect 489306 597156 489374 597212
rect 489430 597156 489498 597212
rect 489554 597156 489622 597212
rect 489678 597156 507250 597212
rect 507306 597156 507374 597212
rect 507430 597156 507498 597212
rect 507554 597156 507622 597212
rect 507678 597156 525250 597212
rect 525306 597156 525374 597212
rect 525430 597156 525498 597212
rect 525554 597156 525622 597212
rect 525678 597156 543250 597212
rect 543306 597156 543374 597212
rect 543430 597156 543498 597212
rect 543554 597156 543622 597212
rect 543678 597156 561250 597212
rect 561306 597156 561374 597212
rect 561430 597156 561498 597212
rect 561554 597156 561622 597212
rect 561678 597156 579250 597212
rect 579306 597156 579374 597212
rect 579430 597156 579498 597212
rect 579554 597156 579622 597212
rect 579678 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 3250 597088
rect 3306 597032 3374 597088
rect 3430 597032 3498 597088
rect 3554 597032 3622 597088
rect 3678 597032 21250 597088
rect 21306 597032 21374 597088
rect 21430 597032 21498 597088
rect 21554 597032 21622 597088
rect 21678 597032 39250 597088
rect 39306 597032 39374 597088
rect 39430 597032 39498 597088
rect 39554 597032 39622 597088
rect 39678 597032 57250 597088
rect 57306 597032 57374 597088
rect 57430 597032 57498 597088
rect 57554 597032 57622 597088
rect 57678 597032 75250 597088
rect 75306 597032 75374 597088
rect 75430 597032 75498 597088
rect 75554 597032 75622 597088
rect 75678 597032 93250 597088
rect 93306 597032 93374 597088
rect 93430 597032 93498 597088
rect 93554 597032 93622 597088
rect 93678 597032 111250 597088
rect 111306 597032 111374 597088
rect 111430 597032 111498 597088
rect 111554 597032 111622 597088
rect 111678 597032 129250 597088
rect 129306 597032 129374 597088
rect 129430 597032 129498 597088
rect 129554 597032 129622 597088
rect 129678 597032 147250 597088
rect 147306 597032 147374 597088
rect 147430 597032 147498 597088
rect 147554 597032 147622 597088
rect 147678 597032 165250 597088
rect 165306 597032 165374 597088
rect 165430 597032 165498 597088
rect 165554 597032 165622 597088
rect 165678 597032 183250 597088
rect 183306 597032 183374 597088
rect 183430 597032 183498 597088
rect 183554 597032 183622 597088
rect 183678 597032 201250 597088
rect 201306 597032 201374 597088
rect 201430 597032 201498 597088
rect 201554 597032 201622 597088
rect 201678 597032 219250 597088
rect 219306 597032 219374 597088
rect 219430 597032 219498 597088
rect 219554 597032 219622 597088
rect 219678 597032 237250 597088
rect 237306 597032 237374 597088
rect 237430 597032 237498 597088
rect 237554 597032 237622 597088
rect 237678 597032 255250 597088
rect 255306 597032 255374 597088
rect 255430 597032 255498 597088
rect 255554 597032 255622 597088
rect 255678 597032 273250 597088
rect 273306 597032 273374 597088
rect 273430 597032 273498 597088
rect 273554 597032 273622 597088
rect 273678 597032 291250 597088
rect 291306 597032 291374 597088
rect 291430 597032 291498 597088
rect 291554 597032 291622 597088
rect 291678 597032 309250 597088
rect 309306 597032 309374 597088
rect 309430 597032 309498 597088
rect 309554 597032 309622 597088
rect 309678 597032 327250 597088
rect 327306 597032 327374 597088
rect 327430 597032 327498 597088
rect 327554 597032 327622 597088
rect 327678 597032 345250 597088
rect 345306 597032 345374 597088
rect 345430 597032 345498 597088
rect 345554 597032 345622 597088
rect 345678 597032 363250 597088
rect 363306 597032 363374 597088
rect 363430 597032 363498 597088
rect 363554 597032 363622 597088
rect 363678 597032 381250 597088
rect 381306 597032 381374 597088
rect 381430 597032 381498 597088
rect 381554 597032 381622 597088
rect 381678 597032 399250 597088
rect 399306 597032 399374 597088
rect 399430 597032 399498 597088
rect 399554 597032 399622 597088
rect 399678 597032 417250 597088
rect 417306 597032 417374 597088
rect 417430 597032 417498 597088
rect 417554 597032 417622 597088
rect 417678 597032 435250 597088
rect 435306 597032 435374 597088
rect 435430 597032 435498 597088
rect 435554 597032 435622 597088
rect 435678 597032 453250 597088
rect 453306 597032 453374 597088
rect 453430 597032 453498 597088
rect 453554 597032 453622 597088
rect 453678 597032 471250 597088
rect 471306 597032 471374 597088
rect 471430 597032 471498 597088
rect 471554 597032 471622 597088
rect 471678 597032 489250 597088
rect 489306 597032 489374 597088
rect 489430 597032 489498 597088
rect 489554 597032 489622 597088
rect 489678 597032 507250 597088
rect 507306 597032 507374 597088
rect 507430 597032 507498 597088
rect 507554 597032 507622 597088
rect 507678 597032 525250 597088
rect 525306 597032 525374 597088
rect 525430 597032 525498 597088
rect 525554 597032 525622 597088
rect 525678 597032 543250 597088
rect 543306 597032 543374 597088
rect 543430 597032 543498 597088
rect 543554 597032 543622 597088
rect 543678 597032 561250 597088
rect 561306 597032 561374 597088
rect 561430 597032 561498 597088
rect 561554 597032 561622 597088
rect 561678 597032 579250 597088
rect 579306 597032 579374 597088
rect 579430 597032 579498 597088
rect 579554 597032 579622 597088
rect 579678 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 3250 596964
rect 3306 596908 3374 596964
rect 3430 596908 3498 596964
rect 3554 596908 3622 596964
rect 3678 596908 21250 596964
rect 21306 596908 21374 596964
rect 21430 596908 21498 596964
rect 21554 596908 21622 596964
rect 21678 596908 39250 596964
rect 39306 596908 39374 596964
rect 39430 596908 39498 596964
rect 39554 596908 39622 596964
rect 39678 596908 57250 596964
rect 57306 596908 57374 596964
rect 57430 596908 57498 596964
rect 57554 596908 57622 596964
rect 57678 596908 75250 596964
rect 75306 596908 75374 596964
rect 75430 596908 75498 596964
rect 75554 596908 75622 596964
rect 75678 596908 93250 596964
rect 93306 596908 93374 596964
rect 93430 596908 93498 596964
rect 93554 596908 93622 596964
rect 93678 596908 111250 596964
rect 111306 596908 111374 596964
rect 111430 596908 111498 596964
rect 111554 596908 111622 596964
rect 111678 596908 129250 596964
rect 129306 596908 129374 596964
rect 129430 596908 129498 596964
rect 129554 596908 129622 596964
rect 129678 596908 147250 596964
rect 147306 596908 147374 596964
rect 147430 596908 147498 596964
rect 147554 596908 147622 596964
rect 147678 596908 165250 596964
rect 165306 596908 165374 596964
rect 165430 596908 165498 596964
rect 165554 596908 165622 596964
rect 165678 596908 183250 596964
rect 183306 596908 183374 596964
rect 183430 596908 183498 596964
rect 183554 596908 183622 596964
rect 183678 596908 201250 596964
rect 201306 596908 201374 596964
rect 201430 596908 201498 596964
rect 201554 596908 201622 596964
rect 201678 596908 219250 596964
rect 219306 596908 219374 596964
rect 219430 596908 219498 596964
rect 219554 596908 219622 596964
rect 219678 596908 237250 596964
rect 237306 596908 237374 596964
rect 237430 596908 237498 596964
rect 237554 596908 237622 596964
rect 237678 596908 255250 596964
rect 255306 596908 255374 596964
rect 255430 596908 255498 596964
rect 255554 596908 255622 596964
rect 255678 596908 273250 596964
rect 273306 596908 273374 596964
rect 273430 596908 273498 596964
rect 273554 596908 273622 596964
rect 273678 596908 291250 596964
rect 291306 596908 291374 596964
rect 291430 596908 291498 596964
rect 291554 596908 291622 596964
rect 291678 596908 309250 596964
rect 309306 596908 309374 596964
rect 309430 596908 309498 596964
rect 309554 596908 309622 596964
rect 309678 596908 327250 596964
rect 327306 596908 327374 596964
rect 327430 596908 327498 596964
rect 327554 596908 327622 596964
rect 327678 596908 345250 596964
rect 345306 596908 345374 596964
rect 345430 596908 345498 596964
rect 345554 596908 345622 596964
rect 345678 596908 363250 596964
rect 363306 596908 363374 596964
rect 363430 596908 363498 596964
rect 363554 596908 363622 596964
rect 363678 596908 381250 596964
rect 381306 596908 381374 596964
rect 381430 596908 381498 596964
rect 381554 596908 381622 596964
rect 381678 596908 399250 596964
rect 399306 596908 399374 596964
rect 399430 596908 399498 596964
rect 399554 596908 399622 596964
rect 399678 596908 417250 596964
rect 417306 596908 417374 596964
rect 417430 596908 417498 596964
rect 417554 596908 417622 596964
rect 417678 596908 435250 596964
rect 435306 596908 435374 596964
rect 435430 596908 435498 596964
rect 435554 596908 435622 596964
rect 435678 596908 453250 596964
rect 453306 596908 453374 596964
rect 453430 596908 453498 596964
rect 453554 596908 453622 596964
rect 453678 596908 471250 596964
rect 471306 596908 471374 596964
rect 471430 596908 471498 596964
rect 471554 596908 471622 596964
rect 471678 596908 489250 596964
rect 489306 596908 489374 596964
rect 489430 596908 489498 596964
rect 489554 596908 489622 596964
rect 489678 596908 507250 596964
rect 507306 596908 507374 596964
rect 507430 596908 507498 596964
rect 507554 596908 507622 596964
rect 507678 596908 525250 596964
rect 525306 596908 525374 596964
rect 525430 596908 525498 596964
rect 525554 596908 525622 596964
rect 525678 596908 543250 596964
rect 543306 596908 543374 596964
rect 543430 596908 543498 596964
rect 543554 596908 543622 596964
rect 543678 596908 561250 596964
rect 561306 596908 561374 596964
rect 561430 596908 561498 596964
rect 561554 596908 561622 596964
rect 561678 596908 579250 596964
rect 579306 596908 579374 596964
rect 579430 596908 579498 596964
rect 579554 596908 579622 596964
rect 579678 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 3250 596840
rect 3306 596784 3374 596840
rect 3430 596784 3498 596840
rect 3554 596784 3622 596840
rect 3678 596784 21250 596840
rect 21306 596784 21374 596840
rect 21430 596784 21498 596840
rect 21554 596784 21622 596840
rect 21678 596784 39250 596840
rect 39306 596784 39374 596840
rect 39430 596784 39498 596840
rect 39554 596784 39622 596840
rect 39678 596784 57250 596840
rect 57306 596784 57374 596840
rect 57430 596784 57498 596840
rect 57554 596784 57622 596840
rect 57678 596784 75250 596840
rect 75306 596784 75374 596840
rect 75430 596784 75498 596840
rect 75554 596784 75622 596840
rect 75678 596784 93250 596840
rect 93306 596784 93374 596840
rect 93430 596784 93498 596840
rect 93554 596784 93622 596840
rect 93678 596784 111250 596840
rect 111306 596784 111374 596840
rect 111430 596784 111498 596840
rect 111554 596784 111622 596840
rect 111678 596784 129250 596840
rect 129306 596784 129374 596840
rect 129430 596784 129498 596840
rect 129554 596784 129622 596840
rect 129678 596784 147250 596840
rect 147306 596784 147374 596840
rect 147430 596784 147498 596840
rect 147554 596784 147622 596840
rect 147678 596784 165250 596840
rect 165306 596784 165374 596840
rect 165430 596784 165498 596840
rect 165554 596784 165622 596840
rect 165678 596784 183250 596840
rect 183306 596784 183374 596840
rect 183430 596784 183498 596840
rect 183554 596784 183622 596840
rect 183678 596784 201250 596840
rect 201306 596784 201374 596840
rect 201430 596784 201498 596840
rect 201554 596784 201622 596840
rect 201678 596784 219250 596840
rect 219306 596784 219374 596840
rect 219430 596784 219498 596840
rect 219554 596784 219622 596840
rect 219678 596784 237250 596840
rect 237306 596784 237374 596840
rect 237430 596784 237498 596840
rect 237554 596784 237622 596840
rect 237678 596784 255250 596840
rect 255306 596784 255374 596840
rect 255430 596784 255498 596840
rect 255554 596784 255622 596840
rect 255678 596784 273250 596840
rect 273306 596784 273374 596840
rect 273430 596784 273498 596840
rect 273554 596784 273622 596840
rect 273678 596784 291250 596840
rect 291306 596784 291374 596840
rect 291430 596784 291498 596840
rect 291554 596784 291622 596840
rect 291678 596784 309250 596840
rect 309306 596784 309374 596840
rect 309430 596784 309498 596840
rect 309554 596784 309622 596840
rect 309678 596784 327250 596840
rect 327306 596784 327374 596840
rect 327430 596784 327498 596840
rect 327554 596784 327622 596840
rect 327678 596784 345250 596840
rect 345306 596784 345374 596840
rect 345430 596784 345498 596840
rect 345554 596784 345622 596840
rect 345678 596784 363250 596840
rect 363306 596784 363374 596840
rect 363430 596784 363498 596840
rect 363554 596784 363622 596840
rect 363678 596784 381250 596840
rect 381306 596784 381374 596840
rect 381430 596784 381498 596840
rect 381554 596784 381622 596840
rect 381678 596784 399250 596840
rect 399306 596784 399374 596840
rect 399430 596784 399498 596840
rect 399554 596784 399622 596840
rect 399678 596784 417250 596840
rect 417306 596784 417374 596840
rect 417430 596784 417498 596840
rect 417554 596784 417622 596840
rect 417678 596784 435250 596840
rect 435306 596784 435374 596840
rect 435430 596784 435498 596840
rect 435554 596784 435622 596840
rect 435678 596784 453250 596840
rect 453306 596784 453374 596840
rect 453430 596784 453498 596840
rect 453554 596784 453622 596840
rect 453678 596784 471250 596840
rect 471306 596784 471374 596840
rect 471430 596784 471498 596840
rect 471554 596784 471622 596840
rect 471678 596784 489250 596840
rect 489306 596784 489374 596840
rect 489430 596784 489498 596840
rect 489554 596784 489622 596840
rect 489678 596784 507250 596840
rect 507306 596784 507374 596840
rect 507430 596784 507498 596840
rect 507554 596784 507622 596840
rect 507678 596784 525250 596840
rect 525306 596784 525374 596840
rect 525430 596784 525498 596840
rect 525554 596784 525622 596840
rect 525678 596784 543250 596840
rect 543306 596784 543374 596840
rect 543430 596784 543498 596840
rect 543554 596784 543622 596840
rect 543678 596784 561250 596840
rect 561306 596784 561374 596840
rect 561430 596784 561498 596840
rect 561554 596784 561622 596840
rect 561678 596784 579250 596840
rect 579306 596784 579374 596840
rect 579430 596784 579498 596840
rect 579554 596784 579622 596840
rect 579678 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 6970 586350
rect 7026 586294 7094 586350
rect 7150 586294 7218 586350
rect 7274 586294 7342 586350
rect 7398 586294 24970 586350
rect 25026 586294 25094 586350
rect 25150 586294 25218 586350
rect 25274 586294 25342 586350
rect 25398 586294 42970 586350
rect 43026 586294 43094 586350
rect 43150 586294 43218 586350
rect 43274 586294 43342 586350
rect 43398 586294 60970 586350
rect 61026 586294 61094 586350
rect 61150 586294 61218 586350
rect 61274 586294 61342 586350
rect 61398 586294 78970 586350
rect 79026 586294 79094 586350
rect 79150 586294 79218 586350
rect 79274 586294 79342 586350
rect 79398 586294 96970 586350
rect 97026 586294 97094 586350
rect 97150 586294 97218 586350
rect 97274 586294 97342 586350
rect 97398 586294 114970 586350
rect 115026 586294 115094 586350
rect 115150 586294 115218 586350
rect 115274 586294 115342 586350
rect 115398 586294 132970 586350
rect 133026 586294 133094 586350
rect 133150 586294 133218 586350
rect 133274 586294 133342 586350
rect 133398 586294 150970 586350
rect 151026 586294 151094 586350
rect 151150 586294 151218 586350
rect 151274 586294 151342 586350
rect 151398 586294 168970 586350
rect 169026 586294 169094 586350
rect 169150 586294 169218 586350
rect 169274 586294 169342 586350
rect 169398 586294 186970 586350
rect 187026 586294 187094 586350
rect 187150 586294 187218 586350
rect 187274 586294 187342 586350
rect 187398 586294 204970 586350
rect 205026 586294 205094 586350
rect 205150 586294 205218 586350
rect 205274 586294 205342 586350
rect 205398 586294 222970 586350
rect 223026 586294 223094 586350
rect 223150 586294 223218 586350
rect 223274 586294 223342 586350
rect 223398 586294 240970 586350
rect 241026 586294 241094 586350
rect 241150 586294 241218 586350
rect 241274 586294 241342 586350
rect 241398 586294 258970 586350
rect 259026 586294 259094 586350
rect 259150 586294 259218 586350
rect 259274 586294 259342 586350
rect 259398 586294 276970 586350
rect 277026 586294 277094 586350
rect 277150 586294 277218 586350
rect 277274 586294 277342 586350
rect 277398 586294 294970 586350
rect 295026 586294 295094 586350
rect 295150 586294 295218 586350
rect 295274 586294 295342 586350
rect 295398 586294 312970 586350
rect 313026 586294 313094 586350
rect 313150 586294 313218 586350
rect 313274 586294 313342 586350
rect 313398 586294 330970 586350
rect 331026 586294 331094 586350
rect 331150 586294 331218 586350
rect 331274 586294 331342 586350
rect 331398 586294 348970 586350
rect 349026 586294 349094 586350
rect 349150 586294 349218 586350
rect 349274 586294 349342 586350
rect 349398 586294 366970 586350
rect 367026 586294 367094 586350
rect 367150 586294 367218 586350
rect 367274 586294 367342 586350
rect 367398 586294 384970 586350
rect 385026 586294 385094 586350
rect 385150 586294 385218 586350
rect 385274 586294 385342 586350
rect 385398 586294 402970 586350
rect 403026 586294 403094 586350
rect 403150 586294 403218 586350
rect 403274 586294 403342 586350
rect 403398 586294 420970 586350
rect 421026 586294 421094 586350
rect 421150 586294 421218 586350
rect 421274 586294 421342 586350
rect 421398 586294 438970 586350
rect 439026 586294 439094 586350
rect 439150 586294 439218 586350
rect 439274 586294 439342 586350
rect 439398 586294 456970 586350
rect 457026 586294 457094 586350
rect 457150 586294 457218 586350
rect 457274 586294 457342 586350
rect 457398 586294 474970 586350
rect 475026 586294 475094 586350
rect 475150 586294 475218 586350
rect 475274 586294 475342 586350
rect 475398 586294 492970 586350
rect 493026 586294 493094 586350
rect 493150 586294 493218 586350
rect 493274 586294 493342 586350
rect 493398 586294 510970 586350
rect 511026 586294 511094 586350
rect 511150 586294 511218 586350
rect 511274 586294 511342 586350
rect 511398 586294 528970 586350
rect 529026 586294 529094 586350
rect 529150 586294 529218 586350
rect 529274 586294 529342 586350
rect 529398 586294 546970 586350
rect 547026 586294 547094 586350
rect 547150 586294 547218 586350
rect 547274 586294 547342 586350
rect 547398 586294 564970 586350
rect 565026 586294 565094 586350
rect 565150 586294 565218 586350
rect 565274 586294 565342 586350
rect 565398 586294 582970 586350
rect 583026 586294 583094 586350
rect 583150 586294 583218 586350
rect 583274 586294 583342 586350
rect 583398 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 6970 586226
rect 7026 586170 7094 586226
rect 7150 586170 7218 586226
rect 7274 586170 7342 586226
rect 7398 586170 24970 586226
rect 25026 586170 25094 586226
rect 25150 586170 25218 586226
rect 25274 586170 25342 586226
rect 25398 586170 42970 586226
rect 43026 586170 43094 586226
rect 43150 586170 43218 586226
rect 43274 586170 43342 586226
rect 43398 586170 60970 586226
rect 61026 586170 61094 586226
rect 61150 586170 61218 586226
rect 61274 586170 61342 586226
rect 61398 586170 78970 586226
rect 79026 586170 79094 586226
rect 79150 586170 79218 586226
rect 79274 586170 79342 586226
rect 79398 586170 96970 586226
rect 97026 586170 97094 586226
rect 97150 586170 97218 586226
rect 97274 586170 97342 586226
rect 97398 586170 114970 586226
rect 115026 586170 115094 586226
rect 115150 586170 115218 586226
rect 115274 586170 115342 586226
rect 115398 586170 132970 586226
rect 133026 586170 133094 586226
rect 133150 586170 133218 586226
rect 133274 586170 133342 586226
rect 133398 586170 150970 586226
rect 151026 586170 151094 586226
rect 151150 586170 151218 586226
rect 151274 586170 151342 586226
rect 151398 586170 168970 586226
rect 169026 586170 169094 586226
rect 169150 586170 169218 586226
rect 169274 586170 169342 586226
rect 169398 586170 186970 586226
rect 187026 586170 187094 586226
rect 187150 586170 187218 586226
rect 187274 586170 187342 586226
rect 187398 586170 204970 586226
rect 205026 586170 205094 586226
rect 205150 586170 205218 586226
rect 205274 586170 205342 586226
rect 205398 586170 222970 586226
rect 223026 586170 223094 586226
rect 223150 586170 223218 586226
rect 223274 586170 223342 586226
rect 223398 586170 240970 586226
rect 241026 586170 241094 586226
rect 241150 586170 241218 586226
rect 241274 586170 241342 586226
rect 241398 586170 258970 586226
rect 259026 586170 259094 586226
rect 259150 586170 259218 586226
rect 259274 586170 259342 586226
rect 259398 586170 276970 586226
rect 277026 586170 277094 586226
rect 277150 586170 277218 586226
rect 277274 586170 277342 586226
rect 277398 586170 294970 586226
rect 295026 586170 295094 586226
rect 295150 586170 295218 586226
rect 295274 586170 295342 586226
rect 295398 586170 312970 586226
rect 313026 586170 313094 586226
rect 313150 586170 313218 586226
rect 313274 586170 313342 586226
rect 313398 586170 330970 586226
rect 331026 586170 331094 586226
rect 331150 586170 331218 586226
rect 331274 586170 331342 586226
rect 331398 586170 348970 586226
rect 349026 586170 349094 586226
rect 349150 586170 349218 586226
rect 349274 586170 349342 586226
rect 349398 586170 366970 586226
rect 367026 586170 367094 586226
rect 367150 586170 367218 586226
rect 367274 586170 367342 586226
rect 367398 586170 384970 586226
rect 385026 586170 385094 586226
rect 385150 586170 385218 586226
rect 385274 586170 385342 586226
rect 385398 586170 402970 586226
rect 403026 586170 403094 586226
rect 403150 586170 403218 586226
rect 403274 586170 403342 586226
rect 403398 586170 420970 586226
rect 421026 586170 421094 586226
rect 421150 586170 421218 586226
rect 421274 586170 421342 586226
rect 421398 586170 438970 586226
rect 439026 586170 439094 586226
rect 439150 586170 439218 586226
rect 439274 586170 439342 586226
rect 439398 586170 456970 586226
rect 457026 586170 457094 586226
rect 457150 586170 457218 586226
rect 457274 586170 457342 586226
rect 457398 586170 474970 586226
rect 475026 586170 475094 586226
rect 475150 586170 475218 586226
rect 475274 586170 475342 586226
rect 475398 586170 492970 586226
rect 493026 586170 493094 586226
rect 493150 586170 493218 586226
rect 493274 586170 493342 586226
rect 493398 586170 510970 586226
rect 511026 586170 511094 586226
rect 511150 586170 511218 586226
rect 511274 586170 511342 586226
rect 511398 586170 528970 586226
rect 529026 586170 529094 586226
rect 529150 586170 529218 586226
rect 529274 586170 529342 586226
rect 529398 586170 546970 586226
rect 547026 586170 547094 586226
rect 547150 586170 547218 586226
rect 547274 586170 547342 586226
rect 547398 586170 564970 586226
rect 565026 586170 565094 586226
rect 565150 586170 565218 586226
rect 565274 586170 565342 586226
rect 565398 586170 582970 586226
rect 583026 586170 583094 586226
rect 583150 586170 583218 586226
rect 583274 586170 583342 586226
rect 583398 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 6970 586102
rect 7026 586046 7094 586102
rect 7150 586046 7218 586102
rect 7274 586046 7342 586102
rect 7398 586046 24970 586102
rect 25026 586046 25094 586102
rect 25150 586046 25218 586102
rect 25274 586046 25342 586102
rect 25398 586046 42970 586102
rect 43026 586046 43094 586102
rect 43150 586046 43218 586102
rect 43274 586046 43342 586102
rect 43398 586046 60970 586102
rect 61026 586046 61094 586102
rect 61150 586046 61218 586102
rect 61274 586046 61342 586102
rect 61398 586046 78970 586102
rect 79026 586046 79094 586102
rect 79150 586046 79218 586102
rect 79274 586046 79342 586102
rect 79398 586046 96970 586102
rect 97026 586046 97094 586102
rect 97150 586046 97218 586102
rect 97274 586046 97342 586102
rect 97398 586046 114970 586102
rect 115026 586046 115094 586102
rect 115150 586046 115218 586102
rect 115274 586046 115342 586102
rect 115398 586046 132970 586102
rect 133026 586046 133094 586102
rect 133150 586046 133218 586102
rect 133274 586046 133342 586102
rect 133398 586046 150970 586102
rect 151026 586046 151094 586102
rect 151150 586046 151218 586102
rect 151274 586046 151342 586102
rect 151398 586046 168970 586102
rect 169026 586046 169094 586102
rect 169150 586046 169218 586102
rect 169274 586046 169342 586102
rect 169398 586046 186970 586102
rect 187026 586046 187094 586102
rect 187150 586046 187218 586102
rect 187274 586046 187342 586102
rect 187398 586046 204970 586102
rect 205026 586046 205094 586102
rect 205150 586046 205218 586102
rect 205274 586046 205342 586102
rect 205398 586046 222970 586102
rect 223026 586046 223094 586102
rect 223150 586046 223218 586102
rect 223274 586046 223342 586102
rect 223398 586046 240970 586102
rect 241026 586046 241094 586102
rect 241150 586046 241218 586102
rect 241274 586046 241342 586102
rect 241398 586046 258970 586102
rect 259026 586046 259094 586102
rect 259150 586046 259218 586102
rect 259274 586046 259342 586102
rect 259398 586046 276970 586102
rect 277026 586046 277094 586102
rect 277150 586046 277218 586102
rect 277274 586046 277342 586102
rect 277398 586046 294970 586102
rect 295026 586046 295094 586102
rect 295150 586046 295218 586102
rect 295274 586046 295342 586102
rect 295398 586046 312970 586102
rect 313026 586046 313094 586102
rect 313150 586046 313218 586102
rect 313274 586046 313342 586102
rect 313398 586046 330970 586102
rect 331026 586046 331094 586102
rect 331150 586046 331218 586102
rect 331274 586046 331342 586102
rect 331398 586046 348970 586102
rect 349026 586046 349094 586102
rect 349150 586046 349218 586102
rect 349274 586046 349342 586102
rect 349398 586046 366970 586102
rect 367026 586046 367094 586102
rect 367150 586046 367218 586102
rect 367274 586046 367342 586102
rect 367398 586046 384970 586102
rect 385026 586046 385094 586102
rect 385150 586046 385218 586102
rect 385274 586046 385342 586102
rect 385398 586046 402970 586102
rect 403026 586046 403094 586102
rect 403150 586046 403218 586102
rect 403274 586046 403342 586102
rect 403398 586046 420970 586102
rect 421026 586046 421094 586102
rect 421150 586046 421218 586102
rect 421274 586046 421342 586102
rect 421398 586046 438970 586102
rect 439026 586046 439094 586102
rect 439150 586046 439218 586102
rect 439274 586046 439342 586102
rect 439398 586046 456970 586102
rect 457026 586046 457094 586102
rect 457150 586046 457218 586102
rect 457274 586046 457342 586102
rect 457398 586046 474970 586102
rect 475026 586046 475094 586102
rect 475150 586046 475218 586102
rect 475274 586046 475342 586102
rect 475398 586046 492970 586102
rect 493026 586046 493094 586102
rect 493150 586046 493218 586102
rect 493274 586046 493342 586102
rect 493398 586046 510970 586102
rect 511026 586046 511094 586102
rect 511150 586046 511218 586102
rect 511274 586046 511342 586102
rect 511398 586046 528970 586102
rect 529026 586046 529094 586102
rect 529150 586046 529218 586102
rect 529274 586046 529342 586102
rect 529398 586046 546970 586102
rect 547026 586046 547094 586102
rect 547150 586046 547218 586102
rect 547274 586046 547342 586102
rect 547398 586046 564970 586102
rect 565026 586046 565094 586102
rect 565150 586046 565218 586102
rect 565274 586046 565342 586102
rect 565398 586046 582970 586102
rect 583026 586046 583094 586102
rect 583150 586046 583218 586102
rect 583274 586046 583342 586102
rect 583398 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 6970 585978
rect 7026 585922 7094 585978
rect 7150 585922 7218 585978
rect 7274 585922 7342 585978
rect 7398 585922 24970 585978
rect 25026 585922 25094 585978
rect 25150 585922 25218 585978
rect 25274 585922 25342 585978
rect 25398 585922 42970 585978
rect 43026 585922 43094 585978
rect 43150 585922 43218 585978
rect 43274 585922 43342 585978
rect 43398 585922 60970 585978
rect 61026 585922 61094 585978
rect 61150 585922 61218 585978
rect 61274 585922 61342 585978
rect 61398 585922 78970 585978
rect 79026 585922 79094 585978
rect 79150 585922 79218 585978
rect 79274 585922 79342 585978
rect 79398 585922 96970 585978
rect 97026 585922 97094 585978
rect 97150 585922 97218 585978
rect 97274 585922 97342 585978
rect 97398 585922 114970 585978
rect 115026 585922 115094 585978
rect 115150 585922 115218 585978
rect 115274 585922 115342 585978
rect 115398 585922 132970 585978
rect 133026 585922 133094 585978
rect 133150 585922 133218 585978
rect 133274 585922 133342 585978
rect 133398 585922 150970 585978
rect 151026 585922 151094 585978
rect 151150 585922 151218 585978
rect 151274 585922 151342 585978
rect 151398 585922 168970 585978
rect 169026 585922 169094 585978
rect 169150 585922 169218 585978
rect 169274 585922 169342 585978
rect 169398 585922 186970 585978
rect 187026 585922 187094 585978
rect 187150 585922 187218 585978
rect 187274 585922 187342 585978
rect 187398 585922 204970 585978
rect 205026 585922 205094 585978
rect 205150 585922 205218 585978
rect 205274 585922 205342 585978
rect 205398 585922 222970 585978
rect 223026 585922 223094 585978
rect 223150 585922 223218 585978
rect 223274 585922 223342 585978
rect 223398 585922 240970 585978
rect 241026 585922 241094 585978
rect 241150 585922 241218 585978
rect 241274 585922 241342 585978
rect 241398 585922 258970 585978
rect 259026 585922 259094 585978
rect 259150 585922 259218 585978
rect 259274 585922 259342 585978
rect 259398 585922 276970 585978
rect 277026 585922 277094 585978
rect 277150 585922 277218 585978
rect 277274 585922 277342 585978
rect 277398 585922 294970 585978
rect 295026 585922 295094 585978
rect 295150 585922 295218 585978
rect 295274 585922 295342 585978
rect 295398 585922 312970 585978
rect 313026 585922 313094 585978
rect 313150 585922 313218 585978
rect 313274 585922 313342 585978
rect 313398 585922 330970 585978
rect 331026 585922 331094 585978
rect 331150 585922 331218 585978
rect 331274 585922 331342 585978
rect 331398 585922 348970 585978
rect 349026 585922 349094 585978
rect 349150 585922 349218 585978
rect 349274 585922 349342 585978
rect 349398 585922 366970 585978
rect 367026 585922 367094 585978
rect 367150 585922 367218 585978
rect 367274 585922 367342 585978
rect 367398 585922 384970 585978
rect 385026 585922 385094 585978
rect 385150 585922 385218 585978
rect 385274 585922 385342 585978
rect 385398 585922 402970 585978
rect 403026 585922 403094 585978
rect 403150 585922 403218 585978
rect 403274 585922 403342 585978
rect 403398 585922 420970 585978
rect 421026 585922 421094 585978
rect 421150 585922 421218 585978
rect 421274 585922 421342 585978
rect 421398 585922 438970 585978
rect 439026 585922 439094 585978
rect 439150 585922 439218 585978
rect 439274 585922 439342 585978
rect 439398 585922 456970 585978
rect 457026 585922 457094 585978
rect 457150 585922 457218 585978
rect 457274 585922 457342 585978
rect 457398 585922 474970 585978
rect 475026 585922 475094 585978
rect 475150 585922 475218 585978
rect 475274 585922 475342 585978
rect 475398 585922 492970 585978
rect 493026 585922 493094 585978
rect 493150 585922 493218 585978
rect 493274 585922 493342 585978
rect 493398 585922 510970 585978
rect 511026 585922 511094 585978
rect 511150 585922 511218 585978
rect 511274 585922 511342 585978
rect 511398 585922 528970 585978
rect 529026 585922 529094 585978
rect 529150 585922 529218 585978
rect 529274 585922 529342 585978
rect 529398 585922 546970 585978
rect 547026 585922 547094 585978
rect 547150 585922 547218 585978
rect 547274 585922 547342 585978
rect 547398 585922 564970 585978
rect 565026 585922 565094 585978
rect 565150 585922 565218 585978
rect 565274 585922 565342 585978
rect 565398 585922 582970 585978
rect 583026 585922 583094 585978
rect 583150 585922 583218 585978
rect 583274 585922 583342 585978
rect 583398 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 3250 580350
rect 3306 580294 3374 580350
rect 3430 580294 3498 580350
rect 3554 580294 3622 580350
rect 3678 580294 21250 580350
rect 21306 580294 21374 580350
rect 21430 580294 21498 580350
rect 21554 580294 21622 580350
rect 21678 580294 39250 580350
rect 39306 580294 39374 580350
rect 39430 580294 39498 580350
rect 39554 580294 39622 580350
rect 39678 580294 57250 580350
rect 57306 580294 57374 580350
rect 57430 580294 57498 580350
rect 57554 580294 57622 580350
rect 57678 580294 75250 580350
rect 75306 580294 75374 580350
rect 75430 580294 75498 580350
rect 75554 580294 75622 580350
rect 75678 580294 93250 580350
rect 93306 580294 93374 580350
rect 93430 580294 93498 580350
rect 93554 580294 93622 580350
rect 93678 580294 111250 580350
rect 111306 580294 111374 580350
rect 111430 580294 111498 580350
rect 111554 580294 111622 580350
rect 111678 580294 129250 580350
rect 129306 580294 129374 580350
rect 129430 580294 129498 580350
rect 129554 580294 129622 580350
rect 129678 580294 147250 580350
rect 147306 580294 147374 580350
rect 147430 580294 147498 580350
rect 147554 580294 147622 580350
rect 147678 580294 165250 580350
rect 165306 580294 165374 580350
rect 165430 580294 165498 580350
rect 165554 580294 165622 580350
rect 165678 580294 183250 580350
rect 183306 580294 183374 580350
rect 183430 580294 183498 580350
rect 183554 580294 183622 580350
rect 183678 580294 201250 580350
rect 201306 580294 201374 580350
rect 201430 580294 201498 580350
rect 201554 580294 201622 580350
rect 201678 580294 219250 580350
rect 219306 580294 219374 580350
rect 219430 580294 219498 580350
rect 219554 580294 219622 580350
rect 219678 580294 237250 580350
rect 237306 580294 237374 580350
rect 237430 580294 237498 580350
rect 237554 580294 237622 580350
rect 237678 580294 255250 580350
rect 255306 580294 255374 580350
rect 255430 580294 255498 580350
rect 255554 580294 255622 580350
rect 255678 580294 273250 580350
rect 273306 580294 273374 580350
rect 273430 580294 273498 580350
rect 273554 580294 273622 580350
rect 273678 580294 291250 580350
rect 291306 580294 291374 580350
rect 291430 580294 291498 580350
rect 291554 580294 291622 580350
rect 291678 580294 309250 580350
rect 309306 580294 309374 580350
rect 309430 580294 309498 580350
rect 309554 580294 309622 580350
rect 309678 580294 327250 580350
rect 327306 580294 327374 580350
rect 327430 580294 327498 580350
rect 327554 580294 327622 580350
rect 327678 580294 345250 580350
rect 345306 580294 345374 580350
rect 345430 580294 345498 580350
rect 345554 580294 345622 580350
rect 345678 580294 363250 580350
rect 363306 580294 363374 580350
rect 363430 580294 363498 580350
rect 363554 580294 363622 580350
rect 363678 580294 381250 580350
rect 381306 580294 381374 580350
rect 381430 580294 381498 580350
rect 381554 580294 381622 580350
rect 381678 580294 399250 580350
rect 399306 580294 399374 580350
rect 399430 580294 399498 580350
rect 399554 580294 399622 580350
rect 399678 580294 417250 580350
rect 417306 580294 417374 580350
rect 417430 580294 417498 580350
rect 417554 580294 417622 580350
rect 417678 580294 435250 580350
rect 435306 580294 435374 580350
rect 435430 580294 435498 580350
rect 435554 580294 435622 580350
rect 435678 580294 453250 580350
rect 453306 580294 453374 580350
rect 453430 580294 453498 580350
rect 453554 580294 453622 580350
rect 453678 580294 471250 580350
rect 471306 580294 471374 580350
rect 471430 580294 471498 580350
rect 471554 580294 471622 580350
rect 471678 580294 489250 580350
rect 489306 580294 489374 580350
rect 489430 580294 489498 580350
rect 489554 580294 489622 580350
rect 489678 580294 507250 580350
rect 507306 580294 507374 580350
rect 507430 580294 507498 580350
rect 507554 580294 507622 580350
rect 507678 580294 525250 580350
rect 525306 580294 525374 580350
rect 525430 580294 525498 580350
rect 525554 580294 525622 580350
rect 525678 580294 543250 580350
rect 543306 580294 543374 580350
rect 543430 580294 543498 580350
rect 543554 580294 543622 580350
rect 543678 580294 561250 580350
rect 561306 580294 561374 580350
rect 561430 580294 561498 580350
rect 561554 580294 561622 580350
rect 561678 580294 579250 580350
rect 579306 580294 579374 580350
rect 579430 580294 579498 580350
rect 579554 580294 579622 580350
rect 579678 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 3250 580226
rect 3306 580170 3374 580226
rect 3430 580170 3498 580226
rect 3554 580170 3622 580226
rect 3678 580170 21250 580226
rect 21306 580170 21374 580226
rect 21430 580170 21498 580226
rect 21554 580170 21622 580226
rect 21678 580170 39250 580226
rect 39306 580170 39374 580226
rect 39430 580170 39498 580226
rect 39554 580170 39622 580226
rect 39678 580170 57250 580226
rect 57306 580170 57374 580226
rect 57430 580170 57498 580226
rect 57554 580170 57622 580226
rect 57678 580170 75250 580226
rect 75306 580170 75374 580226
rect 75430 580170 75498 580226
rect 75554 580170 75622 580226
rect 75678 580170 93250 580226
rect 93306 580170 93374 580226
rect 93430 580170 93498 580226
rect 93554 580170 93622 580226
rect 93678 580170 111250 580226
rect 111306 580170 111374 580226
rect 111430 580170 111498 580226
rect 111554 580170 111622 580226
rect 111678 580170 129250 580226
rect 129306 580170 129374 580226
rect 129430 580170 129498 580226
rect 129554 580170 129622 580226
rect 129678 580170 147250 580226
rect 147306 580170 147374 580226
rect 147430 580170 147498 580226
rect 147554 580170 147622 580226
rect 147678 580170 165250 580226
rect 165306 580170 165374 580226
rect 165430 580170 165498 580226
rect 165554 580170 165622 580226
rect 165678 580170 183250 580226
rect 183306 580170 183374 580226
rect 183430 580170 183498 580226
rect 183554 580170 183622 580226
rect 183678 580170 201250 580226
rect 201306 580170 201374 580226
rect 201430 580170 201498 580226
rect 201554 580170 201622 580226
rect 201678 580170 219250 580226
rect 219306 580170 219374 580226
rect 219430 580170 219498 580226
rect 219554 580170 219622 580226
rect 219678 580170 237250 580226
rect 237306 580170 237374 580226
rect 237430 580170 237498 580226
rect 237554 580170 237622 580226
rect 237678 580170 255250 580226
rect 255306 580170 255374 580226
rect 255430 580170 255498 580226
rect 255554 580170 255622 580226
rect 255678 580170 273250 580226
rect 273306 580170 273374 580226
rect 273430 580170 273498 580226
rect 273554 580170 273622 580226
rect 273678 580170 291250 580226
rect 291306 580170 291374 580226
rect 291430 580170 291498 580226
rect 291554 580170 291622 580226
rect 291678 580170 309250 580226
rect 309306 580170 309374 580226
rect 309430 580170 309498 580226
rect 309554 580170 309622 580226
rect 309678 580170 327250 580226
rect 327306 580170 327374 580226
rect 327430 580170 327498 580226
rect 327554 580170 327622 580226
rect 327678 580170 345250 580226
rect 345306 580170 345374 580226
rect 345430 580170 345498 580226
rect 345554 580170 345622 580226
rect 345678 580170 363250 580226
rect 363306 580170 363374 580226
rect 363430 580170 363498 580226
rect 363554 580170 363622 580226
rect 363678 580170 381250 580226
rect 381306 580170 381374 580226
rect 381430 580170 381498 580226
rect 381554 580170 381622 580226
rect 381678 580170 399250 580226
rect 399306 580170 399374 580226
rect 399430 580170 399498 580226
rect 399554 580170 399622 580226
rect 399678 580170 417250 580226
rect 417306 580170 417374 580226
rect 417430 580170 417498 580226
rect 417554 580170 417622 580226
rect 417678 580170 435250 580226
rect 435306 580170 435374 580226
rect 435430 580170 435498 580226
rect 435554 580170 435622 580226
rect 435678 580170 453250 580226
rect 453306 580170 453374 580226
rect 453430 580170 453498 580226
rect 453554 580170 453622 580226
rect 453678 580170 471250 580226
rect 471306 580170 471374 580226
rect 471430 580170 471498 580226
rect 471554 580170 471622 580226
rect 471678 580170 489250 580226
rect 489306 580170 489374 580226
rect 489430 580170 489498 580226
rect 489554 580170 489622 580226
rect 489678 580170 507250 580226
rect 507306 580170 507374 580226
rect 507430 580170 507498 580226
rect 507554 580170 507622 580226
rect 507678 580170 525250 580226
rect 525306 580170 525374 580226
rect 525430 580170 525498 580226
rect 525554 580170 525622 580226
rect 525678 580170 543250 580226
rect 543306 580170 543374 580226
rect 543430 580170 543498 580226
rect 543554 580170 543622 580226
rect 543678 580170 561250 580226
rect 561306 580170 561374 580226
rect 561430 580170 561498 580226
rect 561554 580170 561622 580226
rect 561678 580170 579250 580226
rect 579306 580170 579374 580226
rect 579430 580170 579498 580226
rect 579554 580170 579622 580226
rect 579678 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 3250 580102
rect 3306 580046 3374 580102
rect 3430 580046 3498 580102
rect 3554 580046 3622 580102
rect 3678 580046 21250 580102
rect 21306 580046 21374 580102
rect 21430 580046 21498 580102
rect 21554 580046 21622 580102
rect 21678 580046 39250 580102
rect 39306 580046 39374 580102
rect 39430 580046 39498 580102
rect 39554 580046 39622 580102
rect 39678 580046 57250 580102
rect 57306 580046 57374 580102
rect 57430 580046 57498 580102
rect 57554 580046 57622 580102
rect 57678 580046 75250 580102
rect 75306 580046 75374 580102
rect 75430 580046 75498 580102
rect 75554 580046 75622 580102
rect 75678 580046 93250 580102
rect 93306 580046 93374 580102
rect 93430 580046 93498 580102
rect 93554 580046 93622 580102
rect 93678 580046 111250 580102
rect 111306 580046 111374 580102
rect 111430 580046 111498 580102
rect 111554 580046 111622 580102
rect 111678 580046 129250 580102
rect 129306 580046 129374 580102
rect 129430 580046 129498 580102
rect 129554 580046 129622 580102
rect 129678 580046 147250 580102
rect 147306 580046 147374 580102
rect 147430 580046 147498 580102
rect 147554 580046 147622 580102
rect 147678 580046 165250 580102
rect 165306 580046 165374 580102
rect 165430 580046 165498 580102
rect 165554 580046 165622 580102
rect 165678 580046 183250 580102
rect 183306 580046 183374 580102
rect 183430 580046 183498 580102
rect 183554 580046 183622 580102
rect 183678 580046 201250 580102
rect 201306 580046 201374 580102
rect 201430 580046 201498 580102
rect 201554 580046 201622 580102
rect 201678 580046 219250 580102
rect 219306 580046 219374 580102
rect 219430 580046 219498 580102
rect 219554 580046 219622 580102
rect 219678 580046 237250 580102
rect 237306 580046 237374 580102
rect 237430 580046 237498 580102
rect 237554 580046 237622 580102
rect 237678 580046 255250 580102
rect 255306 580046 255374 580102
rect 255430 580046 255498 580102
rect 255554 580046 255622 580102
rect 255678 580046 273250 580102
rect 273306 580046 273374 580102
rect 273430 580046 273498 580102
rect 273554 580046 273622 580102
rect 273678 580046 291250 580102
rect 291306 580046 291374 580102
rect 291430 580046 291498 580102
rect 291554 580046 291622 580102
rect 291678 580046 309250 580102
rect 309306 580046 309374 580102
rect 309430 580046 309498 580102
rect 309554 580046 309622 580102
rect 309678 580046 327250 580102
rect 327306 580046 327374 580102
rect 327430 580046 327498 580102
rect 327554 580046 327622 580102
rect 327678 580046 345250 580102
rect 345306 580046 345374 580102
rect 345430 580046 345498 580102
rect 345554 580046 345622 580102
rect 345678 580046 363250 580102
rect 363306 580046 363374 580102
rect 363430 580046 363498 580102
rect 363554 580046 363622 580102
rect 363678 580046 381250 580102
rect 381306 580046 381374 580102
rect 381430 580046 381498 580102
rect 381554 580046 381622 580102
rect 381678 580046 399250 580102
rect 399306 580046 399374 580102
rect 399430 580046 399498 580102
rect 399554 580046 399622 580102
rect 399678 580046 417250 580102
rect 417306 580046 417374 580102
rect 417430 580046 417498 580102
rect 417554 580046 417622 580102
rect 417678 580046 435250 580102
rect 435306 580046 435374 580102
rect 435430 580046 435498 580102
rect 435554 580046 435622 580102
rect 435678 580046 453250 580102
rect 453306 580046 453374 580102
rect 453430 580046 453498 580102
rect 453554 580046 453622 580102
rect 453678 580046 471250 580102
rect 471306 580046 471374 580102
rect 471430 580046 471498 580102
rect 471554 580046 471622 580102
rect 471678 580046 489250 580102
rect 489306 580046 489374 580102
rect 489430 580046 489498 580102
rect 489554 580046 489622 580102
rect 489678 580046 507250 580102
rect 507306 580046 507374 580102
rect 507430 580046 507498 580102
rect 507554 580046 507622 580102
rect 507678 580046 525250 580102
rect 525306 580046 525374 580102
rect 525430 580046 525498 580102
rect 525554 580046 525622 580102
rect 525678 580046 543250 580102
rect 543306 580046 543374 580102
rect 543430 580046 543498 580102
rect 543554 580046 543622 580102
rect 543678 580046 561250 580102
rect 561306 580046 561374 580102
rect 561430 580046 561498 580102
rect 561554 580046 561622 580102
rect 561678 580046 579250 580102
rect 579306 580046 579374 580102
rect 579430 580046 579498 580102
rect 579554 580046 579622 580102
rect 579678 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 3250 579978
rect 3306 579922 3374 579978
rect 3430 579922 3498 579978
rect 3554 579922 3622 579978
rect 3678 579922 21250 579978
rect 21306 579922 21374 579978
rect 21430 579922 21498 579978
rect 21554 579922 21622 579978
rect 21678 579922 39250 579978
rect 39306 579922 39374 579978
rect 39430 579922 39498 579978
rect 39554 579922 39622 579978
rect 39678 579922 57250 579978
rect 57306 579922 57374 579978
rect 57430 579922 57498 579978
rect 57554 579922 57622 579978
rect 57678 579922 75250 579978
rect 75306 579922 75374 579978
rect 75430 579922 75498 579978
rect 75554 579922 75622 579978
rect 75678 579922 93250 579978
rect 93306 579922 93374 579978
rect 93430 579922 93498 579978
rect 93554 579922 93622 579978
rect 93678 579922 111250 579978
rect 111306 579922 111374 579978
rect 111430 579922 111498 579978
rect 111554 579922 111622 579978
rect 111678 579922 129250 579978
rect 129306 579922 129374 579978
rect 129430 579922 129498 579978
rect 129554 579922 129622 579978
rect 129678 579922 147250 579978
rect 147306 579922 147374 579978
rect 147430 579922 147498 579978
rect 147554 579922 147622 579978
rect 147678 579922 165250 579978
rect 165306 579922 165374 579978
rect 165430 579922 165498 579978
rect 165554 579922 165622 579978
rect 165678 579922 183250 579978
rect 183306 579922 183374 579978
rect 183430 579922 183498 579978
rect 183554 579922 183622 579978
rect 183678 579922 201250 579978
rect 201306 579922 201374 579978
rect 201430 579922 201498 579978
rect 201554 579922 201622 579978
rect 201678 579922 219250 579978
rect 219306 579922 219374 579978
rect 219430 579922 219498 579978
rect 219554 579922 219622 579978
rect 219678 579922 237250 579978
rect 237306 579922 237374 579978
rect 237430 579922 237498 579978
rect 237554 579922 237622 579978
rect 237678 579922 255250 579978
rect 255306 579922 255374 579978
rect 255430 579922 255498 579978
rect 255554 579922 255622 579978
rect 255678 579922 273250 579978
rect 273306 579922 273374 579978
rect 273430 579922 273498 579978
rect 273554 579922 273622 579978
rect 273678 579922 291250 579978
rect 291306 579922 291374 579978
rect 291430 579922 291498 579978
rect 291554 579922 291622 579978
rect 291678 579922 309250 579978
rect 309306 579922 309374 579978
rect 309430 579922 309498 579978
rect 309554 579922 309622 579978
rect 309678 579922 327250 579978
rect 327306 579922 327374 579978
rect 327430 579922 327498 579978
rect 327554 579922 327622 579978
rect 327678 579922 345250 579978
rect 345306 579922 345374 579978
rect 345430 579922 345498 579978
rect 345554 579922 345622 579978
rect 345678 579922 363250 579978
rect 363306 579922 363374 579978
rect 363430 579922 363498 579978
rect 363554 579922 363622 579978
rect 363678 579922 381250 579978
rect 381306 579922 381374 579978
rect 381430 579922 381498 579978
rect 381554 579922 381622 579978
rect 381678 579922 399250 579978
rect 399306 579922 399374 579978
rect 399430 579922 399498 579978
rect 399554 579922 399622 579978
rect 399678 579922 417250 579978
rect 417306 579922 417374 579978
rect 417430 579922 417498 579978
rect 417554 579922 417622 579978
rect 417678 579922 435250 579978
rect 435306 579922 435374 579978
rect 435430 579922 435498 579978
rect 435554 579922 435622 579978
rect 435678 579922 453250 579978
rect 453306 579922 453374 579978
rect 453430 579922 453498 579978
rect 453554 579922 453622 579978
rect 453678 579922 471250 579978
rect 471306 579922 471374 579978
rect 471430 579922 471498 579978
rect 471554 579922 471622 579978
rect 471678 579922 489250 579978
rect 489306 579922 489374 579978
rect 489430 579922 489498 579978
rect 489554 579922 489622 579978
rect 489678 579922 507250 579978
rect 507306 579922 507374 579978
rect 507430 579922 507498 579978
rect 507554 579922 507622 579978
rect 507678 579922 525250 579978
rect 525306 579922 525374 579978
rect 525430 579922 525498 579978
rect 525554 579922 525622 579978
rect 525678 579922 543250 579978
rect 543306 579922 543374 579978
rect 543430 579922 543498 579978
rect 543554 579922 543622 579978
rect 543678 579922 561250 579978
rect 561306 579922 561374 579978
rect 561430 579922 561498 579978
rect 561554 579922 561622 579978
rect 561678 579922 579250 579978
rect 579306 579922 579374 579978
rect 579430 579922 579498 579978
rect 579554 579922 579622 579978
rect 579678 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 6970 568350
rect 7026 568294 7094 568350
rect 7150 568294 7218 568350
rect 7274 568294 7342 568350
rect 7398 568294 24970 568350
rect 25026 568294 25094 568350
rect 25150 568294 25218 568350
rect 25274 568294 25342 568350
rect 25398 568294 42970 568350
rect 43026 568294 43094 568350
rect 43150 568294 43218 568350
rect 43274 568294 43342 568350
rect 43398 568294 60970 568350
rect 61026 568294 61094 568350
rect 61150 568294 61218 568350
rect 61274 568294 61342 568350
rect 61398 568294 78970 568350
rect 79026 568294 79094 568350
rect 79150 568294 79218 568350
rect 79274 568294 79342 568350
rect 79398 568294 96970 568350
rect 97026 568294 97094 568350
rect 97150 568294 97218 568350
rect 97274 568294 97342 568350
rect 97398 568294 114970 568350
rect 115026 568294 115094 568350
rect 115150 568294 115218 568350
rect 115274 568294 115342 568350
rect 115398 568294 132970 568350
rect 133026 568294 133094 568350
rect 133150 568294 133218 568350
rect 133274 568294 133342 568350
rect 133398 568294 150970 568350
rect 151026 568294 151094 568350
rect 151150 568294 151218 568350
rect 151274 568294 151342 568350
rect 151398 568294 168970 568350
rect 169026 568294 169094 568350
rect 169150 568294 169218 568350
rect 169274 568294 169342 568350
rect 169398 568294 186970 568350
rect 187026 568294 187094 568350
rect 187150 568294 187218 568350
rect 187274 568294 187342 568350
rect 187398 568294 204970 568350
rect 205026 568294 205094 568350
rect 205150 568294 205218 568350
rect 205274 568294 205342 568350
rect 205398 568294 222970 568350
rect 223026 568294 223094 568350
rect 223150 568294 223218 568350
rect 223274 568294 223342 568350
rect 223398 568294 240970 568350
rect 241026 568294 241094 568350
rect 241150 568294 241218 568350
rect 241274 568294 241342 568350
rect 241398 568294 258970 568350
rect 259026 568294 259094 568350
rect 259150 568294 259218 568350
rect 259274 568294 259342 568350
rect 259398 568294 276970 568350
rect 277026 568294 277094 568350
rect 277150 568294 277218 568350
rect 277274 568294 277342 568350
rect 277398 568294 294970 568350
rect 295026 568294 295094 568350
rect 295150 568294 295218 568350
rect 295274 568294 295342 568350
rect 295398 568294 312970 568350
rect 313026 568294 313094 568350
rect 313150 568294 313218 568350
rect 313274 568294 313342 568350
rect 313398 568294 330970 568350
rect 331026 568294 331094 568350
rect 331150 568294 331218 568350
rect 331274 568294 331342 568350
rect 331398 568294 348970 568350
rect 349026 568294 349094 568350
rect 349150 568294 349218 568350
rect 349274 568294 349342 568350
rect 349398 568294 366970 568350
rect 367026 568294 367094 568350
rect 367150 568294 367218 568350
rect 367274 568294 367342 568350
rect 367398 568294 384970 568350
rect 385026 568294 385094 568350
rect 385150 568294 385218 568350
rect 385274 568294 385342 568350
rect 385398 568294 402970 568350
rect 403026 568294 403094 568350
rect 403150 568294 403218 568350
rect 403274 568294 403342 568350
rect 403398 568294 420970 568350
rect 421026 568294 421094 568350
rect 421150 568294 421218 568350
rect 421274 568294 421342 568350
rect 421398 568294 438970 568350
rect 439026 568294 439094 568350
rect 439150 568294 439218 568350
rect 439274 568294 439342 568350
rect 439398 568294 456970 568350
rect 457026 568294 457094 568350
rect 457150 568294 457218 568350
rect 457274 568294 457342 568350
rect 457398 568294 474970 568350
rect 475026 568294 475094 568350
rect 475150 568294 475218 568350
rect 475274 568294 475342 568350
rect 475398 568294 492970 568350
rect 493026 568294 493094 568350
rect 493150 568294 493218 568350
rect 493274 568294 493342 568350
rect 493398 568294 510970 568350
rect 511026 568294 511094 568350
rect 511150 568294 511218 568350
rect 511274 568294 511342 568350
rect 511398 568294 528970 568350
rect 529026 568294 529094 568350
rect 529150 568294 529218 568350
rect 529274 568294 529342 568350
rect 529398 568294 546970 568350
rect 547026 568294 547094 568350
rect 547150 568294 547218 568350
rect 547274 568294 547342 568350
rect 547398 568294 564970 568350
rect 565026 568294 565094 568350
rect 565150 568294 565218 568350
rect 565274 568294 565342 568350
rect 565398 568294 582970 568350
rect 583026 568294 583094 568350
rect 583150 568294 583218 568350
rect 583274 568294 583342 568350
rect 583398 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 6970 568226
rect 7026 568170 7094 568226
rect 7150 568170 7218 568226
rect 7274 568170 7342 568226
rect 7398 568170 24970 568226
rect 25026 568170 25094 568226
rect 25150 568170 25218 568226
rect 25274 568170 25342 568226
rect 25398 568170 42970 568226
rect 43026 568170 43094 568226
rect 43150 568170 43218 568226
rect 43274 568170 43342 568226
rect 43398 568170 60970 568226
rect 61026 568170 61094 568226
rect 61150 568170 61218 568226
rect 61274 568170 61342 568226
rect 61398 568170 78970 568226
rect 79026 568170 79094 568226
rect 79150 568170 79218 568226
rect 79274 568170 79342 568226
rect 79398 568170 96970 568226
rect 97026 568170 97094 568226
rect 97150 568170 97218 568226
rect 97274 568170 97342 568226
rect 97398 568170 114970 568226
rect 115026 568170 115094 568226
rect 115150 568170 115218 568226
rect 115274 568170 115342 568226
rect 115398 568170 132970 568226
rect 133026 568170 133094 568226
rect 133150 568170 133218 568226
rect 133274 568170 133342 568226
rect 133398 568170 150970 568226
rect 151026 568170 151094 568226
rect 151150 568170 151218 568226
rect 151274 568170 151342 568226
rect 151398 568170 168970 568226
rect 169026 568170 169094 568226
rect 169150 568170 169218 568226
rect 169274 568170 169342 568226
rect 169398 568170 186970 568226
rect 187026 568170 187094 568226
rect 187150 568170 187218 568226
rect 187274 568170 187342 568226
rect 187398 568170 204970 568226
rect 205026 568170 205094 568226
rect 205150 568170 205218 568226
rect 205274 568170 205342 568226
rect 205398 568170 222970 568226
rect 223026 568170 223094 568226
rect 223150 568170 223218 568226
rect 223274 568170 223342 568226
rect 223398 568170 240970 568226
rect 241026 568170 241094 568226
rect 241150 568170 241218 568226
rect 241274 568170 241342 568226
rect 241398 568170 258970 568226
rect 259026 568170 259094 568226
rect 259150 568170 259218 568226
rect 259274 568170 259342 568226
rect 259398 568170 276970 568226
rect 277026 568170 277094 568226
rect 277150 568170 277218 568226
rect 277274 568170 277342 568226
rect 277398 568170 294970 568226
rect 295026 568170 295094 568226
rect 295150 568170 295218 568226
rect 295274 568170 295342 568226
rect 295398 568170 312970 568226
rect 313026 568170 313094 568226
rect 313150 568170 313218 568226
rect 313274 568170 313342 568226
rect 313398 568170 330970 568226
rect 331026 568170 331094 568226
rect 331150 568170 331218 568226
rect 331274 568170 331342 568226
rect 331398 568170 348970 568226
rect 349026 568170 349094 568226
rect 349150 568170 349218 568226
rect 349274 568170 349342 568226
rect 349398 568170 366970 568226
rect 367026 568170 367094 568226
rect 367150 568170 367218 568226
rect 367274 568170 367342 568226
rect 367398 568170 384970 568226
rect 385026 568170 385094 568226
rect 385150 568170 385218 568226
rect 385274 568170 385342 568226
rect 385398 568170 402970 568226
rect 403026 568170 403094 568226
rect 403150 568170 403218 568226
rect 403274 568170 403342 568226
rect 403398 568170 420970 568226
rect 421026 568170 421094 568226
rect 421150 568170 421218 568226
rect 421274 568170 421342 568226
rect 421398 568170 438970 568226
rect 439026 568170 439094 568226
rect 439150 568170 439218 568226
rect 439274 568170 439342 568226
rect 439398 568170 456970 568226
rect 457026 568170 457094 568226
rect 457150 568170 457218 568226
rect 457274 568170 457342 568226
rect 457398 568170 474970 568226
rect 475026 568170 475094 568226
rect 475150 568170 475218 568226
rect 475274 568170 475342 568226
rect 475398 568170 492970 568226
rect 493026 568170 493094 568226
rect 493150 568170 493218 568226
rect 493274 568170 493342 568226
rect 493398 568170 510970 568226
rect 511026 568170 511094 568226
rect 511150 568170 511218 568226
rect 511274 568170 511342 568226
rect 511398 568170 528970 568226
rect 529026 568170 529094 568226
rect 529150 568170 529218 568226
rect 529274 568170 529342 568226
rect 529398 568170 546970 568226
rect 547026 568170 547094 568226
rect 547150 568170 547218 568226
rect 547274 568170 547342 568226
rect 547398 568170 564970 568226
rect 565026 568170 565094 568226
rect 565150 568170 565218 568226
rect 565274 568170 565342 568226
rect 565398 568170 582970 568226
rect 583026 568170 583094 568226
rect 583150 568170 583218 568226
rect 583274 568170 583342 568226
rect 583398 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 6970 568102
rect 7026 568046 7094 568102
rect 7150 568046 7218 568102
rect 7274 568046 7342 568102
rect 7398 568046 24970 568102
rect 25026 568046 25094 568102
rect 25150 568046 25218 568102
rect 25274 568046 25342 568102
rect 25398 568046 42970 568102
rect 43026 568046 43094 568102
rect 43150 568046 43218 568102
rect 43274 568046 43342 568102
rect 43398 568046 60970 568102
rect 61026 568046 61094 568102
rect 61150 568046 61218 568102
rect 61274 568046 61342 568102
rect 61398 568046 78970 568102
rect 79026 568046 79094 568102
rect 79150 568046 79218 568102
rect 79274 568046 79342 568102
rect 79398 568046 96970 568102
rect 97026 568046 97094 568102
rect 97150 568046 97218 568102
rect 97274 568046 97342 568102
rect 97398 568046 114970 568102
rect 115026 568046 115094 568102
rect 115150 568046 115218 568102
rect 115274 568046 115342 568102
rect 115398 568046 132970 568102
rect 133026 568046 133094 568102
rect 133150 568046 133218 568102
rect 133274 568046 133342 568102
rect 133398 568046 150970 568102
rect 151026 568046 151094 568102
rect 151150 568046 151218 568102
rect 151274 568046 151342 568102
rect 151398 568046 168970 568102
rect 169026 568046 169094 568102
rect 169150 568046 169218 568102
rect 169274 568046 169342 568102
rect 169398 568046 186970 568102
rect 187026 568046 187094 568102
rect 187150 568046 187218 568102
rect 187274 568046 187342 568102
rect 187398 568046 204970 568102
rect 205026 568046 205094 568102
rect 205150 568046 205218 568102
rect 205274 568046 205342 568102
rect 205398 568046 222970 568102
rect 223026 568046 223094 568102
rect 223150 568046 223218 568102
rect 223274 568046 223342 568102
rect 223398 568046 240970 568102
rect 241026 568046 241094 568102
rect 241150 568046 241218 568102
rect 241274 568046 241342 568102
rect 241398 568046 258970 568102
rect 259026 568046 259094 568102
rect 259150 568046 259218 568102
rect 259274 568046 259342 568102
rect 259398 568046 276970 568102
rect 277026 568046 277094 568102
rect 277150 568046 277218 568102
rect 277274 568046 277342 568102
rect 277398 568046 294970 568102
rect 295026 568046 295094 568102
rect 295150 568046 295218 568102
rect 295274 568046 295342 568102
rect 295398 568046 312970 568102
rect 313026 568046 313094 568102
rect 313150 568046 313218 568102
rect 313274 568046 313342 568102
rect 313398 568046 330970 568102
rect 331026 568046 331094 568102
rect 331150 568046 331218 568102
rect 331274 568046 331342 568102
rect 331398 568046 348970 568102
rect 349026 568046 349094 568102
rect 349150 568046 349218 568102
rect 349274 568046 349342 568102
rect 349398 568046 366970 568102
rect 367026 568046 367094 568102
rect 367150 568046 367218 568102
rect 367274 568046 367342 568102
rect 367398 568046 384970 568102
rect 385026 568046 385094 568102
rect 385150 568046 385218 568102
rect 385274 568046 385342 568102
rect 385398 568046 402970 568102
rect 403026 568046 403094 568102
rect 403150 568046 403218 568102
rect 403274 568046 403342 568102
rect 403398 568046 420970 568102
rect 421026 568046 421094 568102
rect 421150 568046 421218 568102
rect 421274 568046 421342 568102
rect 421398 568046 438970 568102
rect 439026 568046 439094 568102
rect 439150 568046 439218 568102
rect 439274 568046 439342 568102
rect 439398 568046 456970 568102
rect 457026 568046 457094 568102
rect 457150 568046 457218 568102
rect 457274 568046 457342 568102
rect 457398 568046 474970 568102
rect 475026 568046 475094 568102
rect 475150 568046 475218 568102
rect 475274 568046 475342 568102
rect 475398 568046 492970 568102
rect 493026 568046 493094 568102
rect 493150 568046 493218 568102
rect 493274 568046 493342 568102
rect 493398 568046 510970 568102
rect 511026 568046 511094 568102
rect 511150 568046 511218 568102
rect 511274 568046 511342 568102
rect 511398 568046 528970 568102
rect 529026 568046 529094 568102
rect 529150 568046 529218 568102
rect 529274 568046 529342 568102
rect 529398 568046 546970 568102
rect 547026 568046 547094 568102
rect 547150 568046 547218 568102
rect 547274 568046 547342 568102
rect 547398 568046 564970 568102
rect 565026 568046 565094 568102
rect 565150 568046 565218 568102
rect 565274 568046 565342 568102
rect 565398 568046 582970 568102
rect 583026 568046 583094 568102
rect 583150 568046 583218 568102
rect 583274 568046 583342 568102
rect 583398 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 6970 567978
rect 7026 567922 7094 567978
rect 7150 567922 7218 567978
rect 7274 567922 7342 567978
rect 7398 567922 24970 567978
rect 25026 567922 25094 567978
rect 25150 567922 25218 567978
rect 25274 567922 25342 567978
rect 25398 567922 42970 567978
rect 43026 567922 43094 567978
rect 43150 567922 43218 567978
rect 43274 567922 43342 567978
rect 43398 567922 60970 567978
rect 61026 567922 61094 567978
rect 61150 567922 61218 567978
rect 61274 567922 61342 567978
rect 61398 567922 78970 567978
rect 79026 567922 79094 567978
rect 79150 567922 79218 567978
rect 79274 567922 79342 567978
rect 79398 567922 96970 567978
rect 97026 567922 97094 567978
rect 97150 567922 97218 567978
rect 97274 567922 97342 567978
rect 97398 567922 114970 567978
rect 115026 567922 115094 567978
rect 115150 567922 115218 567978
rect 115274 567922 115342 567978
rect 115398 567922 132970 567978
rect 133026 567922 133094 567978
rect 133150 567922 133218 567978
rect 133274 567922 133342 567978
rect 133398 567922 150970 567978
rect 151026 567922 151094 567978
rect 151150 567922 151218 567978
rect 151274 567922 151342 567978
rect 151398 567922 168970 567978
rect 169026 567922 169094 567978
rect 169150 567922 169218 567978
rect 169274 567922 169342 567978
rect 169398 567922 186970 567978
rect 187026 567922 187094 567978
rect 187150 567922 187218 567978
rect 187274 567922 187342 567978
rect 187398 567922 204970 567978
rect 205026 567922 205094 567978
rect 205150 567922 205218 567978
rect 205274 567922 205342 567978
rect 205398 567922 222970 567978
rect 223026 567922 223094 567978
rect 223150 567922 223218 567978
rect 223274 567922 223342 567978
rect 223398 567922 240970 567978
rect 241026 567922 241094 567978
rect 241150 567922 241218 567978
rect 241274 567922 241342 567978
rect 241398 567922 258970 567978
rect 259026 567922 259094 567978
rect 259150 567922 259218 567978
rect 259274 567922 259342 567978
rect 259398 567922 276970 567978
rect 277026 567922 277094 567978
rect 277150 567922 277218 567978
rect 277274 567922 277342 567978
rect 277398 567922 294970 567978
rect 295026 567922 295094 567978
rect 295150 567922 295218 567978
rect 295274 567922 295342 567978
rect 295398 567922 312970 567978
rect 313026 567922 313094 567978
rect 313150 567922 313218 567978
rect 313274 567922 313342 567978
rect 313398 567922 330970 567978
rect 331026 567922 331094 567978
rect 331150 567922 331218 567978
rect 331274 567922 331342 567978
rect 331398 567922 348970 567978
rect 349026 567922 349094 567978
rect 349150 567922 349218 567978
rect 349274 567922 349342 567978
rect 349398 567922 366970 567978
rect 367026 567922 367094 567978
rect 367150 567922 367218 567978
rect 367274 567922 367342 567978
rect 367398 567922 384970 567978
rect 385026 567922 385094 567978
rect 385150 567922 385218 567978
rect 385274 567922 385342 567978
rect 385398 567922 402970 567978
rect 403026 567922 403094 567978
rect 403150 567922 403218 567978
rect 403274 567922 403342 567978
rect 403398 567922 420970 567978
rect 421026 567922 421094 567978
rect 421150 567922 421218 567978
rect 421274 567922 421342 567978
rect 421398 567922 438970 567978
rect 439026 567922 439094 567978
rect 439150 567922 439218 567978
rect 439274 567922 439342 567978
rect 439398 567922 456970 567978
rect 457026 567922 457094 567978
rect 457150 567922 457218 567978
rect 457274 567922 457342 567978
rect 457398 567922 474970 567978
rect 475026 567922 475094 567978
rect 475150 567922 475218 567978
rect 475274 567922 475342 567978
rect 475398 567922 492970 567978
rect 493026 567922 493094 567978
rect 493150 567922 493218 567978
rect 493274 567922 493342 567978
rect 493398 567922 510970 567978
rect 511026 567922 511094 567978
rect 511150 567922 511218 567978
rect 511274 567922 511342 567978
rect 511398 567922 528970 567978
rect 529026 567922 529094 567978
rect 529150 567922 529218 567978
rect 529274 567922 529342 567978
rect 529398 567922 546970 567978
rect 547026 567922 547094 567978
rect 547150 567922 547218 567978
rect 547274 567922 547342 567978
rect 547398 567922 564970 567978
rect 565026 567922 565094 567978
rect 565150 567922 565218 567978
rect 565274 567922 565342 567978
rect 565398 567922 582970 567978
rect 583026 567922 583094 567978
rect 583150 567922 583218 567978
rect 583274 567922 583342 567978
rect 583398 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 3250 562350
rect 3306 562294 3374 562350
rect 3430 562294 3498 562350
rect 3554 562294 3622 562350
rect 3678 562294 21250 562350
rect 21306 562294 21374 562350
rect 21430 562294 21498 562350
rect 21554 562294 21622 562350
rect 21678 562294 39250 562350
rect 39306 562294 39374 562350
rect 39430 562294 39498 562350
rect 39554 562294 39622 562350
rect 39678 562294 57250 562350
rect 57306 562294 57374 562350
rect 57430 562294 57498 562350
rect 57554 562294 57622 562350
rect 57678 562294 75250 562350
rect 75306 562294 75374 562350
rect 75430 562294 75498 562350
rect 75554 562294 75622 562350
rect 75678 562294 93250 562350
rect 93306 562294 93374 562350
rect 93430 562294 93498 562350
rect 93554 562294 93622 562350
rect 93678 562294 111250 562350
rect 111306 562294 111374 562350
rect 111430 562294 111498 562350
rect 111554 562294 111622 562350
rect 111678 562294 129250 562350
rect 129306 562294 129374 562350
rect 129430 562294 129498 562350
rect 129554 562294 129622 562350
rect 129678 562294 147250 562350
rect 147306 562294 147374 562350
rect 147430 562294 147498 562350
rect 147554 562294 147622 562350
rect 147678 562294 165250 562350
rect 165306 562294 165374 562350
rect 165430 562294 165498 562350
rect 165554 562294 165622 562350
rect 165678 562294 183250 562350
rect 183306 562294 183374 562350
rect 183430 562294 183498 562350
rect 183554 562294 183622 562350
rect 183678 562294 201250 562350
rect 201306 562294 201374 562350
rect 201430 562294 201498 562350
rect 201554 562294 201622 562350
rect 201678 562294 219250 562350
rect 219306 562294 219374 562350
rect 219430 562294 219498 562350
rect 219554 562294 219622 562350
rect 219678 562294 237250 562350
rect 237306 562294 237374 562350
rect 237430 562294 237498 562350
rect 237554 562294 237622 562350
rect 237678 562294 255250 562350
rect 255306 562294 255374 562350
rect 255430 562294 255498 562350
rect 255554 562294 255622 562350
rect 255678 562294 273250 562350
rect 273306 562294 273374 562350
rect 273430 562294 273498 562350
rect 273554 562294 273622 562350
rect 273678 562294 291250 562350
rect 291306 562294 291374 562350
rect 291430 562294 291498 562350
rect 291554 562294 291622 562350
rect 291678 562294 309250 562350
rect 309306 562294 309374 562350
rect 309430 562294 309498 562350
rect 309554 562294 309622 562350
rect 309678 562294 327250 562350
rect 327306 562294 327374 562350
rect 327430 562294 327498 562350
rect 327554 562294 327622 562350
rect 327678 562294 345250 562350
rect 345306 562294 345374 562350
rect 345430 562294 345498 562350
rect 345554 562294 345622 562350
rect 345678 562294 363250 562350
rect 363306 562294 363374 562350
rect 363430 562294 363498 562350
rect 363554 562294 363622 562350
rect 363678 562294 381250 562350
rect 381306 562294 381374 562350
rect 381430 562294 381498 562350
rect 381554 562294 381622 562350
rect 381678 562294 399250 562350
rect 399306 562294 399374 562350
rect 399430 562294 399498 562350
rect 399554 562294 399622 562350
rect 399678 562294 417250 562350
rect 417306 562294 417374 562350
rect 417430 562294 417498 562350
rect 417554 562294 417622 562350
rect 417678 562294 435250 562350
rect 435306 562294 435374 562350
rect 435430 562294 435498 562350
rect 435554 562294 435622 562350
rect 435678 562294 453250 562350
rect 453306 562294 453374 562350
rect 453430 562294 453498 562350
rect 453554 562294 453622 562350
rect 453678 562294 471250 562350
rect 471306 562294 471374 562350
rect 471430 562294 471498 562350
rect 471554 562294 471622 562350
rect 471678 562294 489250 562350
rect 489306 562294 489374 562350
rect 489430 562294 489498 562350
rect 489554 562294 489622 562350
rect 489678 562294 507250 562350
rect 507306 562294 507374 562350
rect 507430 562294 507498 562350
rect 507554 562294 507622 562350
rect 507678 562294 525250 562350
rect 525306 562294 525374 562350
rect 525430 562294 525498 562350
rect 525554 562294 525622 562350
rect 525678 562294 543250 562350
rect 543306 562294 543374 562350
rect 543430 562294 543498 562350
rect 543554 562294 543622 562350
rect 543678 562294 561250 562350
rect 561306 562294 561374 562350
rect 561430 562294 561498 562350
rect 561554 562294 561622 562350
rect 561678 562294 579250 562350
rect 579306 562294 579374 562350
rect 579430 562294 579498 562350
rect 579554 562294 579622 562350
rect 579678 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 3250 562226
rect 3306 562170 3374 562226
rect 3430 562170 3498 562226
rect 3554 562170 3622 562226
rect 3678 562170 21250 562226
rect 21306 562170 21374 562226
rect 21430 562170 21498 562226
rect 21554 562170 21622 562226
rect 21678 562170 39250 562226
rect 39306 562170 39374 562226
rect 39430 562170 39498 562226
rect 39554 562170 39622 562226
rect 39678 562170 57250 562226
rect 57306 562170 57374 562226
rect 57430 562170 57498 562226
rect 57554 562170 57622 562226
rect 57678 562170 75250 562226
rect 75306 562170 75374 562226
rect 75430 562170 75498 562226
rect 75554 562170 75622 562226
rect 75678 562170 93250 562226
rect 93306 562170 93374 562226
rect 93430 562170 93498 562226
rect 93554 562170 93622 562226
rect 93678 562170 111250 562226
rect 111306 562170 111374 562226
rect 111430 562170 111498 562226
rect 111554 562170 111622 562226
rect 111678 562170 129250 562226
rect 129306 562170 129374 562226
rect 129430 562170 129498 562226
rect 129554 562170 129622 562226
rect 129678 562170 147250 562226
rect 147306 562170 147374 562226
rect 147430 562170 147498 562226
rect 147554 562170 147622 562226
rect 147678 562170 165250 562226
rect 165306 562170 165374 562226
rect 165430 562170 165498 562226
rect 165554 562170 165622 562226
rect 165678 562170 183250 562226
rect 183306 562170 183374 562226
rect 183430 562170 183498 562226
rect 183554 562170 183622 562226
rect 183678 562170 201250 562226
rect 201306 562170 201374 562226
rect 201430 562170 201498 562226
rect 201554 562170 201622 562226
rect 201678 562170 219250 562226
rect 219306 562170 219374 562226
rect 219430 562170 219498 562226
rect 219554 562170 219622 562226
rect 219678 562170 237250 562226
rect 237306 562170 237374 562226
rect 237430 562170 237498 562226
rect 237554 562170 237622 562226
rect 237678 562170 255250 562226
rect 255306 562170 255374 562226
rect 255430 562170 255498 562226
rect 255554 562170 255622 562226
rect 255678 562170 273250 562226
rect 273306 562170 273374 562226
rect 273430 562170 273498 562226
rect 273554 562170 273622 562226
rect 273678 562170 291250 562226
rect 291306 562170 291374 562226
rect 291430 562170 291498 562226
rect 291554 562170 291622 562226
rect 291678 562170 309250 562226
rect 309306 562170 309374 562226
rect 309430 562170 309498 562226
rect 309554 562170 309622 562226
rect 309678 562170 327250 562226
rect 327306 562170 327374 562226
rect 327430 562170 327498 562226
rect 327554 562170 327622 562226
rect 327678 562170 345250 562226
rect 345306 562170 345374 562226
rect 345430 562170 345498 562226
rect 345554 562170 345622 562226
rect 345678 562170 363250 562226
rect 363306 562170 363374 562226
rect 363430 562170 363498 562226
rect 363554 562170 363622 562226
rect 363678 562170 381250 562226
rect 381306 562170 381374 562226
rect 381430 562170 381498 562226
rect 381554 562170 381622 562226
rect 381678 562170 399250 562226
rect 399306 562170 399374 562226
rect 399430 562170 399498 562226
rect 399554 562170 399622 562226
rect 399678 562170 417250 562226
rect 417306 562170 417374 562226
rect 417430 562170 417498 562226
rect 417554 562170 417622 562226
rect 417678 562170 435250 562226
rect 435306 562170 435374 562226
rect 435430 562170 435498 562226
rect 435554 562170 435622 562226
rect 435678 562170 453250 562226
rect 453306 562170 453374 562226
rect 453430 562170 453498 562226
rect 453554 562170 453622 562226
rect 453678 562170 471250 562226
rect 471306 562170 471374 562226
rect 471430 562170 471498 562226
rect 471554 562170 471622 562226
rect 471678 562170 489250 562226
rect 489306 562170 489374 562226
rect 489430 562170 489498 562226
rect 489554 562170 489622 562226
rect 489678 562170 507250 562226
rect 507306 562170 507374 562226
rect 507430 562170 507498 562226
rect 507554 562170 507622 562226
rect 507678 562170 525250 562226
rect 525306 562170 525374 562226
rect 525430 562170 525498 562226
rect 525554 562170 525622 562226
rect 525678 562170 543250 562226
rect 543306 562170 543374 562226
rect 543430 562170 543498 562226
rect 543554 562170 543622 562226
rect 543678 562170 561250 562226
rect 561306 562170 561374 562226
rect 561430 562170 561498 562226
rect 561554 562170 561622 562226
rect 561678 562170 579250 562226
rect 579306 562170 579374 562226
rect 579430 562170 579498 562226
rect 579554 562170 579622 562226
rect 579678 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 3250 562102
rect 3306 562046 3374 562102
rect 3430 562046 3498 562102
rect 3554 562046 3622 562102
rect 3678 562046 21250 562102
rect 21306 562046 21374 562102
rect 21430 562046 21498 562102
rect 21554 562046 21622 562102
rect 21678 562046 39250 562102
rect 39306 562046 39374 562102
rect 39430 562046 39498 562102
rect 39554 562046 39622 562102
rect 39678 562046 57250 562102
rect 57306 562046 57374 562102
rect 57430 562046 57498 562102
rect 57554 562046 57622 562102
rect 57678 562046 75250 562102
rect 75306 562046 75374 562102
rect 75430 562046 75498 562102
rect 75554 562046 75622 562102
rect 75678 562046 93250 562102
rect 93306 562046 93374 562102
rect 93430 562046 93498 562102
rect 93554 562046 93622 562102
rect 93678 562046 111250 562102
rect 111306 562046 111374 562102
rect 111430 562046 111498 562102
rect 111554 562046 111622 562102
rect 111678 562046 129250 562102
rect 129306 562046 129374 562102
rect 129430 562046 129498 562102
rect 129554 562046 129622 562102
rect 129678 562046 147250 562102
rect 147306 562046 147374 562102
rect 147430 562046 147498 562102
rect 147554 562046 147622 562102
rect 147678 562046 165250 562102
rect 165306 562046 165374 562102
rect 165430 562046 165498 562102
rect 165554 562046 165622 562102
rect 165678 562046 183250 562102
rect 183306 562046 183374 562102
rect 183430 562046 183498 562102
rect 183554 562046 183622 562102
rect 183678 562046 201250 562102
rect 201306 562046 201374 562102
rect 201430 562046 201498 562102
rect 201554 562046 201622 562102
rect 201678 562046 219250 562102
rect 219306 562046 219374 562102
rect 219430 562046 219498 562102
rect 219554 562046 219622 562102
rect 219678 562046 237250 562102
rect 237306 562046 237374 562102
rect 237430 562046 237498 562102
rect 237554 562046 237622 562102
rect 237678 562046 255250 562102
rect 255306 562046 255374 562102
rect 255430 562046 255498 562102
rect 255554 562046 255622 562102
rect 255678 562046 273250 562102
rect 273306 562046 273374 562102
rect 273430 562046 273498 562102
rect 273554 562046 273622 562102
rect 273678 562046 291250 562102
rect 291306 562046 291374 562102
rect 291430 562046 291498 562102
rect 291554 562046 291622 562102
rect 291678 562046 309250 562102
rect 309306 562046 309374 562102
rect 309430 562046 309498 562102
rect 309554 562046 309622 562102
rect 309678 562046 327250 562102
rect 327306 562046 327374 562102
rect 327430 562046 327498 562102
rect 327554 562046 327622 562102
rect 327678 562046 345250 562102
rect 345306 562046 345374 562102
rect 345430 562046 345498 562102
rect 345554 562046 345622 562102
rect 345678 562046 363250 562102
rect 363306 562046 363374 562102
rect 363430 562046 363498 562102
rect 363554 562046 363622 562102
rect 363678 562046 381250 562102
rect 381306 562046 381374 562102
rect 381430 562046 381498 562102
rect 381554 562046 381622 562102
rect 381678 562046 399250 562102
rect 399306 562046 399374 562102
rect 399430 562046 399498 562102
rect 399554 562046 399622 562102
rect 399678 562046 417250 562102
rect 417306 562046 417374 562102
rect 417430 562046 417498 562102
rect 417554 562046 417622 562102
rect 417678 562046 435250 562102
rect 435306 562046 435374 562102
rect 435430 562046 435498 562102
rect 435554 562046 435622 562102
rect 435678 562046 453250 562102
rect 453306 562046 453374 562102
rect 453430 562046 453498 562102
rect 453554 562046 453622 562102
rect 453678 562046 471250 562102
rect 471306 562046 471374 562102
rect 471430 562046 471498 562102
rect 471554 562046 471622 562102
rect 471678 562046 489250 562102
rect 489306 562046 489374 562102
rect 489430 562046 489498 562102
rect 489554 562046 489622 562102
rect 489678 562046 507250 562102
rect 507306 562046 507374 562102
rect 507430 562046 507498 562102
rect 507554 562046 507622 562102
rect 507678 562046 525250 562102
rect 525306 562046 525374 562102
rect 525430 562046 525498 562102
rect 525554 562046 525622 562102
rect 525678 562046 543250 562102
rect 543306 562046 543374 562102
rect 543430 562046 543498 562102
rect 543554 562046 543622 562102
rect 543678 562046 561250 562102
rect 561306 562046 561374 562102
rect 561430 562046 561498 562102
rect 561554 562046 561622 562102
rect 561678 562046 579250 562102
rect 579306 562046 579374 562102
rect 579430 562046 579498 562102
rect 579554 562046 579622 562102
rect 579678 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 3250 561978
rect 3306 561922 3374 561978
rect 3430 561922 3498 561978
rect 3554 561922 3622 561978
rect 3678 561922 21250 561978
rect 21306 561922 21374 561978
rect 21430 561922 21498 561978
rect 21554 561922 21622 561978
rect 21678 561922 39250 561978
rect 39306 561922 39374 561978
rect 39430 561922 39498 561978
rect 39554 561922 39622 561978
rect 39678 561922 57250 561978
rect 57306 561922 57374 561978
rect 57430 561922 57498 561978
rect 57554 561922 57622 561978
rect 57678 561922 75250 561978
rect 75306 561922 75374 561978
rect 75430 561922 75498 561978
rect 75554 561922 75622 561978
rect 75678 561922 93250 561978
rect 93306 561922 93374 561978
rect 93430 561922 93498 561978
rect 93554 561922 93622 561978
rect 93678 561922 111250 561978
rect 111306 561922 111374 561978
rect 111430 561922 111498 561978
rect 111554 561922 111622 561978
rect 111678 561922 129250 561978
rect 129306 561922 129374 561978
rect 129430 561922 129498 561978
rect 129554 561922 129622 561978
rect 129678 561922 147250 561978
rect 147306 561922 147374 561978
rect 147430 561922 147498 561978
rect 147554 561922 147622 561978
rect 147678 561922 165250 561978
rect 165306 561922 165374 561978
rect 165430 561922 165498 561978
rect 165554 561922 165622 561978
rect 165678 561922 183250 561978
rect 183306 561922 183374 561978
rect 183430 561922 183498 561978
rect 183554 561922 183622 561978
rect 183678 561922 201250 561978
rect 201306 561922 201374 561978
rect 201430 561922 201498 561978
rect 201554 561922 201622 561978
rect 201678 561922 219250 561978
rect 219306 561922 219374 561978
rect 219430 561922 219498 561978
rect 219554 561922 219622 561978
rect 219678 561922 237250 561978
rect 237306 561922 237374 561978
rect 237430 561922 237498 561978
rect 237554 561922 237622 561978
rect 237678 561922 255250 561978
rect 255306 561922 255374 561978
rect 255430 561922 255498 561978
rect 255554 561922 255622 561978
rect 255678 561922 273250 561978
rect 273306 561922 273374 561978
rect 273430 561922 273498 561978
rect 273554 561922 273622 561978
rect 273678 561922 291250 561978
rect 291306 561922 291374 561978
rect 291430 561922 291498 561978
rect 291554 561922 291622 561978
rect 291678 561922 309250 561978
rect 309306 561922 309374 561978
rect 309430 561922 309498 561978
rect 309554 561922 309622 561978
rect 309678 561922 327250 561978
rect 327306 561922 327374 561978
rect 327430 561922 327498 561978
rect 327554 561922 327622 561978
rect 327678 561922 345250 561978
rect 345306 561922 345374 561978
rect 345430 561922 345498 561978
rect 345554 561922 345622 561978
rect 345678 561922 363250 561978
rect 363306 561922 363374 561978
rect 363430 561922 363498 561978
rect 363554 561922 363622 561978
rect 363678 561922 381250 561978
rect 381306 561922 381374 561978
rect 381430 561922 381498 561978
rect 381554 561922 381622 561978
rect 381678 561922 399250 561978
rect 399306 561922 399374 561978
rect 399430 561922 399498 561978
rect 399554 561922 399622 561978
rect 399678 561922 417250 561978
rect 417306 561922 417374 561978
rect 417430 561922 417498 561978
rect 417554 561922 417622 561978
rect 417678 561922 435250 561978
rect 435306 561922 435374 561978
rect 435430 561922 435498 561978
rect 435554 561922 435622 561978
rect 435678 561922 453250 561978
rect 453306 561922 453374 561978
rect 453430 561922 453498 561978
rect 453554 561922 453622 561978
rect 453678 561922 471250 561978
rect 471306 561922 471374 561978
rect 471430 561922 471498 561978
rect 471554 561922 471622 561978
rect 471678 561922 489250 561978
rect 489306 561922 489374 561978
rect 489430 561922 489498 561978
rect 489554 561922 489622 561978
rect 489678 561922 507250 561978
rect 507306 561922 507374 561978
rect 507430 561922 507498 561978
rect 507554 561922 507622 561978
rect 507678 561922 525250 561978
rect 525306 561922 525374 561978
rect 525430 561922 525498 561978
rect 525554 561922 525622 561978
rect 525678 561922 543250 561978
rect 543306 561922 543374 561978
rect 543430 561922 543498 561978
rect 543554 561922 543622 561978
rect 543678 561922 561250 561978
rect 561306 561922 561374 561978
rect 561430 561922 561498 561978
rect 561554 561922 561622 561978
rect 561678 561922 579250 561978
rect 579306 561922 579374 561978
rect 579430 561922 579498 561978
rect 579554 561922 579622 561978
rect 579678 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 6970 550350
rect 7026 550294 7094 550350
rect 7150 550294 7218 550350
rect 7274 550294 7342 550350
rect 7398 550294 24970 550350
rect 25026 550294 25094 550350
rect 25150 550294 25218 550350
rect 25274 550294 25342 550350
rect 25398 550294 42970 550350
rect 43026 550294 43094 550350
rect 43150 550294 43218 550350
rect 43274 550294 43342 550350
rect 43398 550294 60970 550350
rect 61026 550294 61094 550350
rect 61150 550294 61218 550350
rect 61274 550294 61342 550350
rect 61398 550294 78970 550350
rect 79026 550294 79094 550350
rect 79150 550294 79218 550350
rect 79274 550294 79342 550350
rect 79398 550294 96970 550350
rect 97026 550294 97094 550350
rect 97150 550294 97218 550350
rect 97274 550294 97342 550350
rect 97398 550294 114970 550350
rect 115026 550294 115094 550350
rect 115150 550294 115218 550350
rect 115274 550294 115342 550350
rect 115398 550294 132970 550350
rect 133026 550294 133094 550350
rect 133150 550294 133218 550350
rect 133274 550294 133342 550350
rect 133398 550294 150970 550350
rect 151026 550294 151094 550350
rect 151150 550294 151218 550350
rect 151274 550294 151342 550350
rect 151398 550294 168970 550350
rect 169026 550294 169094 550350
rect 169150 550294 169218 550350
rect 169274 550294 169342 550350
rect 169398 550294 186970 550350
rect 187026 550294 187094 550350
rect 187150 550294 187218 550350
rect 187274 550294 187342 550350
rect 187398 550294 204970 550350
rect 205026 550294 205094 550350
rect 205150 550294 205218 550350
rect 205274 550294 205342 550350
rect 205398 550294 222970 550350
rect 223026 550294 223094 550350
rect 223150 550294 223218 550350
rect 223274 550294 223342 550350
rect 223398 550294 240970 550350
rect 241026 550294 241094 550350
rect 241150 550294 241218 550350
rect 241274 550294 241342 550350
rect 241398 550294 258970 550350
rect 259026 550294 259094 550350
rect 259150 550294 259218 550350
rect 259274 550294 259342 550350
rect 259398 550294 276970 550350
rect 277026 550294 277094 550350
rect 277150 550294 277218 550350
rect 277274 550294 277342 550350
rect 277398 550294 294970 550350
rect 295026 550294 295094 550350
rect 295150 550294 295218 550350
rect 295274 550294 295342 550350
rect 295398 550294 312970 550350
rect 313026 550294 313094 550350
rect 313150 550294 313218 550350
rect 313274 550294 313342 550350
rect 313398 550294 330970 550350
rect 331026 550294 331094 550350
rect 331150 550294 331218 550350
rect 331274 550294 331342 550350
rect 331398 550294 348970 550350
rect 349026 550294 349094 550350
rect 349150 550294 349218 550350
rect 349274 550294 349342 550350
rect 349398 550294 366970 550350
rect 367026 550294 367094 550350
rect 367150 550294 367218 550350
rect 367274 550294 367342 550350
rect 367398 550294 384970 550350
rect 385026 550294 385094 550350
rect 385150 550294 385218 550350
rect 385274 550294 385342 550350
rect 385398 550294 402970 550350
rect 403026 550294 403094 550350
rect 403150 550294 403218 550350
rect 403274 550294 403342 550350
rect 403398 550294 420970 550350
rect 421026 550294 421094 550350
rect 421150 550294 421218 550350
rect 421274 550294 421342 550350
rect 421398 550294 438970 550350
rect 439026 550294 439094 550350
rect 439150 550294 439218 550350
rect 439274 550294 439342 550350
rect 439398 550294 456970 550350
rect 457026 550294 457094 550350
rect 457150 550294 457218 550350
rect 457274 550294 457342 550350
rect 457398 550294 474970 550350
rect 475026 550294 475094 550350
rect 475150 550294 475218 550350
rect 475274 550294 475342 550350
rect 475398 550294 492970 550350
rect 493026 550294 493094 550350
rect 493150 550294 493218 550350
rect 493274 550294 493342 550350
rect 493398 550294 510970 550350
rect 511026 550294 511094 550350
rect 511150 550294 511218 550350
rect 511274 550294 511342 550350
rect 511398 550294 528970 550350
rect 529026 550294 529094 550350
rect 529150 550294 529218 550350
rect 529274 550294 529342 550350
rect 529398 550294 546970 550350
rect 547026 550294 547094 550350
rect 547150 550294 547218 550350
rect 547274 550294 547342 550350
rect 547398 550294 564970 550350
rect 565026 550294 565094 550350
rect 565150 550294 565218 550350
rect 565274 550294 565342 550350
rect 565398 550294 582970 550350
rect 583026 550294 583094 550350
rect 583150 550294 583218 550350
rect 583274 550294 583342 550350
rect 583398 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 6970 550226
rect 7026 550170 7094 550226
rect 7150 550170 7218 550226
rect 7274 550170 7342 550226
rect 7398 550170 24970 550226
rect 25026 550170 25094 550226
rect 25150 550170 25218 550226
rect 25274 550170 25342 550226
rect 25398 550170 42970 550226
rect 43026 550170 43094 550226
rect 43150 550170 43218 550226
rect 43274 550170 43342 550226
rect 43398 550170 60970 550226
rect 61026 550170 61094 550226
rect 61150 550170 61218 550226
rect 61274 550170 61342 550226
rect 61398 550170 78970 550226
rect 79026 550170 79094 550226
rect 79150 550170 79218 550226
rect 79274 550170 79342 550226
rect 79398 550170 96970 550226
rect 97026 550170 97094 550226
rect 97150 550170 97218 550226
rect 97274 550170 97342 550226
rect 97398 550170 114970 550226
rect 115026 550170 115094 550226
rect 115150 550170 115218 550226
rect 115274 550170 115342 550226
rect 115398 550170 132970 550226
rect 133026 550170 133094 550226
rect 133150 550170 133218 550226
rect 133274 550170 133342 550226
rect 133398 550170 150970 550226
rect 151026 550170 151094 550226
rect 151150 550170 151218 550226
rect 151274 550170 151342 550226
rect 151398 550170 168970 550226
rect 169026 550170 169094 550226
rect 169150 550170 169218 550226
rect 169274 550170 169342 550226
rect 169398 550170 186970 550226
rect 187026 550170 187094 550226
rect 187150 550170 187218 550226
rect 187274 550170 187342 550226
rect 187398 550170 204970 550226
rect 205026 550170 205094 550226
rect 205150 550170 205218 550226
rect 205274 550170 205342 550226
rect 205398 550170 222970 550226
rect 223026 550170 223094 550226
rect 223150 550170 223218 550226
rect 223274 550170 223342 550226
rect 223398 550170 240970 550226
rect 241026 550170 241094 550226
rect 241150 550170 241218 550226
rect 241274 550170 241342 550226
rect 241398 550170 258970 550226
rect 259026 550170 259094 550226
rect 259150 550170 259218 550226
rect 259274 550170 259342 550226
rect 259398 550170 276970 550226
rect 277026 550170 277094 550226
rect 277150 550170 277218 550226
rect 277274 550170 277342 550226
rect 277398 550170 294970 550226
rect 295026 550170 295094 550226
rect 295150 550170 295218 550226
rect 295274 550170 295342 550226
rect 295398 550170 312970 550226
rect 313026 550170 313094 550226
rect 313150 550170 313218 550226
rect 313274 550170 313342 550226
rect 313398 550170 330970 550226
rect 331026 550170 331094 550226
rect 331150 550170 331218 550226
rect 331274 550170 331342 550226
rect 331398 550170 348970 550226
rect 349026 550170 349094 550226
rect 349150 550170 349218 550226
rect 349274 550170 349342 550226
rect 349398 550170 366970 550226
rect 367026 550170 367094 550226
rect 367150 550170 367218 550226
rect 367274 550170 367342 550226
rect 367398 550170 384970 550226
rect 385026 550170 385094 550226
rect 385150 550170 385218 550226
rect 385274 550170 385342 550226
rect 385398 550170 402970 550226
rect 403026 550170 403094 550226
rect 403150 550170 403218 550226
rect 403274 550170 403342 550226
rect 403398 550170 420970 550226
rect 421026 550170 421094 550226
rect 421150 550170 421218 550226
rect 421274 550170 421342 550226
rect 421398 550170 438970 550226
rect 439026 550170 439094 550226
rect 439150 550170 439218 550226
rect 439274 550170 439342 550226
rect 439398 550170 456970 550226
rect 457026 550170 457094 550226
rect 457150 550170 457218 550226
rect 457274 550170 457342 550226
rect 457398 550170 474970 550226
rect 475026 550170 475094 550226
rect 475150 550170 475218 550226
rect 475274 550170 475342 550226
rect 475398 550170 492970 550226
rect 493026 550170 493094 550226
rect 493150 550170 493218 550226
rect 493274 550170 493342 550226
rect 493398 550170 510970 550226
rect 511026 550170 511094 550226
rect 511150 550170 511218 550226
rect 511274 550170 511342 550226
rect 511398 550170 528970 550226
rect 529026 550170 529094 550226
rect 529150 550170 529218 550226
rect 529274 550170 529342 550226
rect 529398 550170 546970 550226
rect 547026 550170 547094 550226
rect 547150 550170 547218 550226
rect 547274 550170 547342 550226
rect 547398 550170 564970 550226
rect 565026 550170 565094 550226
rect 565150 550170 565218 550226
rect 565274 550170 565342 550226
rect 565398 550170 582970 550226
rect 583026 550170 583094 550226
rect 583150 550170 583218 550226
rect 583274 550170 583342 550226
rect 583398 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 6970 550102
rect 7026 550046 7094 550102
rect 7150 550046 7218 550102
rect 7274 550046 7342 550102
rect 7398 550046 24970 550102
rect 25026 550046 25094 550102
rect 25150 550046 25218 550102
rect 25274 550046 25342 550102
rect 25398 550046 42970 550102
rect 43026 550046 43094 550102
rect 43150 550046 43218 550102
rect 43274 550046 43342 550102
rect 43398 550046 60970 550102
rect 61026 550046 61094 550102
rect 61150 550046 61218 550102
rect 61274 550046 61342 550102
rect 61398 550046 78970 550102
rect 79026 550046 79094 550102
rect 79150 550046 79218 550102
rect 79274 550046 79342 550102
rect 79398 550046 96970 550102
rect 97026 550046 97094 550102
rect 97150 550046 97218 550102
rect 97274 550046 97342 550102
rect 97398 550046 114970 550102
rect 115026 550046 115094 550102
rect 115150 550046 115218 550102
rect 115274 550046 115342 550102
rect 115398 550046 132970 550102
rect 133026 550046 133094 550102
rect 133150 550046 133218 550102
rect 133274 550046 133342 550102
rect 133398 550046 150970 550102
rect 151026 550046 151094 550102
rect 151150 550046 151218 550102
rect 151274 550046 151342 550102
rect 151398 550046 168970 550102
rect 169026 550046 169094 550102
rect 169150 550046 169218 550102
rect 169274 550046 169342 550102
rect 169398 550046 186970 550102
rect 187026 550046 187094 550102
rect 187150 550046 187218 550102
rect 187274 550046 187342 550102
rect 187398 550046 204970 550102
rect 205026 550046 205094 550102
rect 205150 550046 205218 550102
rect 205274 550046 205342 550102
rect 205398 550046 222970 550102
rect 223026 550046 223094 550102
rect 223150 550046 223218 550102
rect 223274 550046 223342 550102
rect 223398 550046 240970 550102
rect 241026 550046 241094 550102
rect 241150 550046 241218 550102
rect 241274 550046 241342 550102
rect 241398 550046 258970 550102
rect 259026 550046 259094 550102
rect 259150 550046 259218 550102
rect 259274 550046 259342 550102
rect 259398 550046 276970 550102
rect 277026 550046 277094 550102
rect 277150 550046 277218 550102
rect 277274 550046 277342 550102
rect 277398 550046 294970 550102
rect 295026 550046 295094 550102
rect 295150 550046 295218 550102
rect 295274 550046 295342 550102
rect 295398 550046 312970 550102
rect 313026 550046 313094 550102
rect 313150 550046 313218 550102
rect 313274 550046 313342 550102
rect 313398 550046 330970 550102
rect 331026 550046 331094 550102
rect 331150 550046 331218 550102
rect 331274 550046 331342 550102
rect 331398 550046 348970 550102
rect 349026 550046 349094 550102
rect 349150 550046 349218 550102
rect 349274 550046 349342 550102
rect 349398 550046 366970 550102
rect 367026 550046 367094 550102
rect 367150 550046 367218 550102
rect 367274 550046 367342 550102
rect 367398 550046 384970 550102
rect 385026 550046 385094 550102
rect 385150 550046 385218 550102
rect 385274 550046 385342 550102
rect 385398 550046 402970 550102
rect 403026 550046 403094 550102
rect 403150 550046 403218 550102
rect 403274 550046 403342 550102
rect 403398 550046 420970 550102
rect 421026 550046 421094 550102
rect 421150 550046 421218 550102
rect 421274 550046 421342 550102
rect 421398 550046 438970 550102
rect 439026 550046 439094 550102
rect 439150 550046 439218 550102
rect 439274 550046 439342 550102
rect 439398 550046 456970 550102
rect 457026 550046 457094 550102
rect 457150 550046 457218 550102
rect 457274 550046 457342 550102
rect 457398 550046 474970 550102
rect 475026 550046 475094 550102
rect 475150 550046 475218 550102
rect 475274 550046 475342 550102
rect 475398 550046 492970 550102
rect 493026 550046 493094 550102
rect 493150 550046 493218 550102
rect 493274 550046 493342 550102
rect 493398 550046 510970 550102
rect 511026 550046 511094 550102
rect 511150 550046 511218 550102
rect 511274 550046 511342 550102
rect 511398 550046 528970 550102
rect 529026 550046 529094 550102
rect 529150 550046 529218 550102
rect 529274 550046 529342 550102
rect 529398 550046 546970 550102
rect 547026 550046 547094 550102
rect 547150 550046 547218 550102
rect 547274 550046 547342 550102
rect 547398 550046 564970 550102
rect 565026 550046 565094 550102
rect 565150 550046 565218 550102
rect 565274 550046 565342 550102
rect 565398 550046 582970 550102
rect 583026 550046 583094 550102
rect 583150 550046 583218 550102
rect 583274 550046 583342 550102
rect 583398 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 6970 549978
rect 7026 549922 7094 549978
rect 7150 549922 7218 549978
rect 7274 549922 7342 549978
rect 7398 549922 24970 549978
rect 25026 549922 25094 549978
rect 25150 549922 25218 549978
rect 25274 549922 25342 549978
rect 25398 549922 42970 549978
rect 43026 549922 43094 549978
rect 43150 549922 43218 549978
rect 43274 549922 43342 549978
rect 43398 549922 60970 549978
rect 61026 549922 61094 549978
rect 61150 549922 61218 549978
rect 61274 549922 61342 549978
rect 61398 549922 78970 549978
rect 79026 549922 79094 549978
rect 79150 549922 79218 549978
rect 79274 549922 79342 549978
rect 79398 549922 96970 549978
rect 97026 549922 97094 549978
rect 97150 549922 97218 549978
rect 97274 549922 97342 549978
rect 97398 549922 114970 549978
rect 115026 549922 115094 549978
rect 115150 549922 115218 549978
rect 115274 549922 115342 549978
rect 115398 549922 132970 549978
rect 133026 549922 133094 549978
rect 133150 549922 133218 549978
rect 133274 549922 133342 549978
rect 133398 549922 150970 549978
rect 151026 549922 151094 549978
rect 151150 549922 151218 549978
rect 151274 549922 151342 549978
rect 151398 549922 168970 549978
rect 169026 549922 169094 549978
rect 169150 549922 169218 549978
rect 169274 549922 169342 549978
rect 169398 549922 186970 549978
rect 187026 549922 187094 549978
rect 187150 549922 187218 549978
rect 187274 549922 187342 549978
rect 187398 549922 204970 549978
rect 205026 549922 205094 549978
rect 205150 549922 205218 549978
rect 205274 549922 205342 549978
rect 205398 549922 222970 549978
rect 223026 549922 223094 549978
rect 223150 549922 223218 549978
rect 223274 549922 223342 549978
rect 223398 549922 240970 549978
rect 241026 549922 241094 549978
rect 241150 549922 241218 549978
rect 241274 549922 241342 549978
rect 241398 549922 258970 549978
rect 259026 549922 259094 549978
rect 259150 549922 259218 549978
rect 259274 549922 259342 549978
rect 259398 549922 276970 549978
rect 277026 549922 277094 549978
rect 277150 549922 277218 549978
rect 277274 549922 277342 549978
rect 277398 549922 294970 549978
rect 295026 549922 295094 549978
rect 295150 549922 295218 549978
rect 295274 549922 295342 549978
rect 295398 549922 312970 549978
rect 313026 549922 313094 549978
rect 313150 549922 313218 549978
rect 313274 549922 313342 549978
rect 313398 549922 330970 549978
rect 331026 549922 331094 549978
rect 331150 549922 331218 549978
rect 331274 549922 331342 549978
rect 331398 549922 348970 549978
rect 349026 549922 349094 549978
rect 349150 549922 349218 549978
rect 349274 549922 349342 549978
rect 349398 549922 366970 549978
rect 367026 549922 367094 549978
rect 367150 549922 367218 549978
rect 367274 549922 367342 549978
rect 367398 549922 384970 549978
rect 385026 549922 385094 549978
rect 385150 549922 385218 549978
rect 385274 549922 385342 549978
rect 385398 549922 402970 549978
rect 403026 549922 403094 549978
rect 403150 549922 403218 549978
rect 403274 549922 403342 549978
rect 403398 549922 420970 549978
rect 421026 549922 421094 549978
rect 421150 549922 421218 549978
rect 421274 549922 421342 549978
rect 421398 549922 438970 549978
rect 439026 549922 439094 549978
rect 439150 549922 439218 549978
rect 439274 549922 439342 549978
rect 439398 549922 456970 549978
rect 457026 549922 457094 549978
rect 457150 549922 457218 549978
rect 457274 549922 457342 549978
rect 457398 549922 474970 549978
rect 475026 549922 475094 549978
rect 475150 549922 475218 549978
rect 475274 549922 475342 549978
rect 475398 549922 492970 549978
rect 493026 549922 493094 549978
rect 493150 549922 493218 549978
rect 493274 549922 493342 549978
rect 493398 549922 510970 549978
rect 511026 549922 511094 549978
rect 511150 549922 511218 549978
rect 511274 549922 511342 549978
rect 511398 549922 528970 549978
rect 529026 549922 529094 549978
rect 529150 549922 529218 549978
rect 529274 549922 529342 549978
rect 529398 549922 546970 549978
rect 547026 549922 547094 549978
rect 547150 549922 547218 549978
rect 547274 549922 547342 549978
rect 547398 549922 564970 549978
rect 565026 549922 565094 549978
rect 565150 549922 565218 549978
rect 565274 549922 565342 549978
rect 565398 549922 582970 549978
rect 583026 549922 583094 549978
rect 583150 549922 583218 549978
rect 583274 549922 583342 549978
rect 583398 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 3250 544350
rect 3306 544294 3374 544350
rect 3430 544294 3498 544350
rect 3554 544294 3622 544350
rect 3678 544294 21250 544350
rect 21306 544294 21374 544350
rect 21430 544294 21498 544350
rect 21554 544294 21622 544350
rect 21678 544294 39250 544350
rect 39306 544294 39374 544350
rect 39430 544294 39498 544350
rect 39554 544294 39622 544350
rect 39678 544294 57250 544350
rect 57306 544294 57374 544350
rect 57430 544294 57498 544350
rect 57554 544294 57622 544350
rect 57678 544294 75250 544350
rect 75306 544294 75374 544350
rect 75430 544294 75498 544350
rect 75554 544294 75622 544350
rect 75678 544294 93250 544350
rect 93306 544294 93374 544350
rect 93430 544294 93498 544350
rect 93554 544294 93622 544350
rect 93678 544294 111250 544350
rect 111306 544294 111374 544350
rect 111430 544294 111498 544350
rect 111554 544294 111622 544350
rect 111678 544294 129250 544350
rect 129306 544294 129374 544350
rect 129430 544294 129498 544350
rect 129554 544294 129622 544350
rect 129678 544294 147250 544350
rect 147306 544294 147374 544350
rect 147430 544294 147498 544350
rect 147554 544294 147622 544350
rect 147678 544294 165250 544350
rect 165306 544294 165374 544350
rect 165430 544294 165498 544350
rect 165554 544294 165622 544350
rect 165678 544294 183250 544350
rect 183306 544294 183374 544350
rect 183430 544294 183498 544350
rect 183554 544294 183622 544350
rect 183678 544294 201250 544350
rect 201306 544294 201374 544350
rect 201430 544294 201498 544350
rect 201554 544294 201622 544350
rect 201678 544294 219250 544350
rect 219306 544294 219374 544350
rect 219430 544294 219498 544350
rect 219554 544294 219622 544350
rect 219678 544294 237250 544350
rect 237306 544294 237374 544350
rect 237430 544294 237498 544350
rect 237554 544294 237622 544350
rect 237678 544294 255250 544350
rect 255306 544294 255374 544350
rect 255430 544294 255498 544350
rect 255554 544294 255622 544350
rect 255678 544294 273250 544350
rect 273306 544294 273374 544350
rect 273430 544294 273498 544350
rect 273554 544294 273622 544350
rect 273678 544294 291250 544350
rect 291306 544294 291374 544350
rect 291430 544294 291498 544350
rect 291554 544294 291622 544350
rect 291678 544294 309250 544350
rect 309306 544294 309374 544350
rect 309430 544294 309498 544350
rect 309554 544294 309622 544350
rect 309678 544294 327250 544350
rect 327306 544294 327374 544350
rect 327430 544294 327498 544350
rect 327554 544294 327622 544350
rect 327678 544294 345250 544350
rect 345306 544294 345374 544350
rect 345430 544294 345498 544350
rect 345554 544294 345622 544350
rect 345678 544294 363250 544350
rect 363306 544294 363374 544350
rect 363430 544294 363498 544350
rect 363554 544294 363622 544350
rect 363678 544294 381250 544350
rect 381306 544294 381374 544350
rect 381430 544294 381498 544350
rect 381554 544294 381622 544350
rect 381678 544294 399250 544350
rect 399306 544294 399374 544350
rect 399430 544294 399498 544350
rect 399554 544294 399622 544350
rect 399678 544294 417250 544350
rect 417306 544294 417374 544350
rect 417430 544294 417498 544350
rect 417554 544294 417622 544350
rect 417678 544294 435250 544350
rect 435306 544294 435374 544350
rect 435430 544294 435498 544350
rect 435554 544294 435622 544350
rect 435678 544294 453250 544350
rect 453306 544294 453374 544350
rect 453430 544294 453498 544350
rect 453554 544294 453622 544350
rect 453678 544294 471250 544350
rect 471306 544294 471374 544350
rect 471430 544294 471498 544350
rect 471554 544294 471622 544350
rect 471678 544294 489250 544350
rect 489306 544294 489374 544350
rect 489430 544294 489498 544350
rect 489554 544294 489622 544350
rect 489678 544294 507250 544350
rect 507306 544294 507374 544350
rect 507430 544294 507498 544350
rect 507554 544294 507622 544350
rect 507678 544294 525250 544350
rect 525306 544294 525374 544350
rect 525430 544294 525498 544350
rect 525554 544294 525622 544350
rect 525678 544294 543250 544350
rect 543306 544294 543374 544350
rect 543430 544294 543498 544350
rect 543554 544294 543622 544350
rect 543678 544294 561250 544350
rect 561306 544294 561374 544350
rect 561430 544294 561498 544350
rect 561554 544294 561622 544350
rect 561678 544294 579250 544350
rect 579306 544294 579374 544350
rect 579430 544294 579498 544350
rect 579554 544294 579622 544350
rect 579678 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 3250 544226
rect 3306 544170 3374 544226
rect 3430 544170 3498 544226
rect 3554 544170 3622 544226
rect 3678 544170 21250 544226
rect 21306 544170 21374 544226
rect 21430 544170 21498 544226
rect 21554 544170 21622 544226
rect 21678 544170 39250 544226
rect 39306 544170 39374 544226
rect 39430 544170 39498 544226
rect 39554 544170 39622 544226
rect 39678 544170 57250 544226
rect 57306 544170 57374 544226
rect 57430 544170 57498 544226
rect 57554 544170 57622 544226
rect 57678 544170 75250 544226
rect 75306 544170 75374 544226
rect 75430 544170 75498 544226
rect 75554 544170 75622 544226
rect 75678 544170 93250 544226
rect 93306 544170 93374 544226
rect 93430 544170 93498 544226
rect 93554 544170 93622 544226
rect 93678 544170 111250 544226
rect 111306 544170 111374 544226
rect 111430 544170 111498 544226
rect 111554 544170 111622 544226
rect 111678 544170 129250 544226
rect 129306 544170 129374 544226
rect 129430 544170 129498 544226
rect 129554 544170 129622 544226
rect 129678 544170 147250 544226
rect 147306 544170 147374 544226
rect 147430 544170 147498 544226
rect 147554 544170 147622 544226
rect 147678 544170 165250 544226
rect 165306 544170 165374 544226
rect 165430 544170 165498 544226
rect 165554 544170 165622 544226
rect 165678 544170 183250 544226
rect 183306 544170 183374 544226
rect 183430 544170 183498 544226
rect 183554 544170 183622 544226
rect 183678 544170 201250 544226
rect 201306 544170 201374 544226
rect 201430 544170 201498 544226
rect 201554 544170 201622 544226
rect 201678 544170 219250 544226
rect 219306 544170 219374 544226
rect 219430 544170 219498 544226
rect 219554 544170 219622 544226
rect 219678 544170 237250 544226
rect 237306 544170 237374 544226
rect 237430 544170 237498 544226
rect 237554 544170 237622 544226
rect 237678 544170 255250 544226
rect 255306 544170 255374 544226
rect 255430 544170 255498 544226
rect 255554 544170 255622 544226
rect 255678 544170 273250 544226
rect 273306 544170 273374 544226
rect 273430 544170 273498 544226
rect 273554 544170 273622 544226
rect 273678 544170 291250 544226
rect 291306 544170 291374 544226
rect 291430 544170 291498 544226
rect 291554 544170 291622 544226
rect 291678 544170 309250 544226
rect 309306 544170 309374 544226
rect 309430 544170 309498 544226
rect 309554 544170 309622 544226
rect 309678 544170 327250 544226
rect 327306 544170 327374 544226
rect 327430 544170 327498 544226
rect 327554 544170 327622 544226
rect 327678 544170 345250 544226
rect 345306 544170 345374 544226
rect 345430 544170 345498 544226
rect 345554 544170 345622 544226
rect 345678 544170 363250 544226
rect 363306 544170 363374 544226
rect 363430 544170 363498 544226
rect 363554 544170 363622 544226
rect 363678 544170 381250 544226
rect 381306 544170 381374 544226
rect 381430 544170 381498 544226
rect 381554 544170 381622 544226
rect 381678 544170 399250 544226
rect 399306 544170 399374 544226
rect 399430 544170 399498 544226
rect 399554 544170 399622 544226
rect 399678 544170 417250 544226
rect 417306 544170 417374 544226
rect 417430 544170 417498 544226
rect 417554 544170 417622 544226
rect 417678 544170 435250 544226
rect 435306 544170 435374 544226
rect 435430 544170 435498 544226
rect 435554 544170 435622 544226
rect 435678 544170 453250 544226
rect 453306 544170 453374 544226
rect 453430 544170 453498 544226
rect 453554 544170 453622 544226
rect 453678 544170 471250 544226
rect 471306 544170 471374 544226
rect 471430 544170 471498 544226
rect 471554 544170 471622 544226
rect 471678 544170 489250 544226
rect 489306 544170 489374 544226
rect 489430 544170 489498 544226
rect 489554 544170 489622 544226
rect 489678 544170 507250 544226
rect 507306 544170 507374 544226
rect 507430 544170 507498 544226
rect 507554 544170 507622 544226
rect 507678 544170 525250 544226
rect 525306 544170 525374 544226
rect 525430 544170 525498 544226
rect 525554 544170 525622 544226
rect 525678 544170 543250 544226
rect 543306 544170 543374 544226
rect 543430 544170 543498 544226
rect 543554 544170 543622 544226
rect 543678 544170 561250 544226
rect 561306 544170 561374 544226
rect 561430 544170 561498 544226
rect 561554 544170 561622 544226
rect 561678 544170 579250 544226
rect 579306 544170 579374 544226
rect 579430 544170 579498 544226
rect 579554 544170 579622 544226
rect 579678 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 3250 544102
rect 3306 544046 3374 544102
rect 3430 544046 3498 544102
rect 3554 544046 3622 544102
rect 3678 544046 21250 544102
rect 21306 544046 21374 544102
rect 21430 544046 21498 544102
rect 21554 544046 21622 544102
rect 21678 544046 39250 544102
rect 39306 544046 39374 544102
rect 39430 544046 39498 544102
rect 39554 544046 39622 544102
rect 39678 544046 57250 544102
rect 57306 544046 57374 544102
rect 57430 544046 57498 544102
rect 57554 544046 57622 544102
rect 57678 544046 75250 544102
rect 75306 544046 75374 544102
rect 75430 544046 75498 544102
rect 75554 544046 75622 544102
rect 75678 544046 93250 544102
rect 93306 544046 93374 544102
rect 93430 544046 93498 544102
rect 93554 544046 93622 544102
rect 93678 544046 111250 544102
rect 111306 544046 111374 544102
rect 111430 544046 111498 544102
rect 111554 544046 111622 544102
rect 111678 544046 129250 544102
rect 129306 544046 129374 544102
rect 129430 544046 129498 544102
rect 129554 544046 129622 544102
rect 129678 544046 147250 544102
rect 147306 544046 147374 544102
rect 147430 544046 147498 544102
rect 147554 544046 147622 544102
rect 147678 544046 165250 544102
rect 165306 544046 165374 544102
rect 165430 544046 165498 544102
rect 165554 544046 165622 544102
rect 165678 544046 183250 544102
rect 183306 544046 183374 544102
rect 183430 544046 183498 544102
rect 183554 544046 183622 544102
rect 183678 544046 201250 544102
rect 201306 544046 201374 544102
rect 201430 544046 201498 544102
rect 201554 544046 201622 544102
rect 201678 544046 219250 544102
rect 219306 544046 219374 544102
rect 219430 544046 219498 544102
rect 219554 544046 219622 544102
rect 219678 544046 237250 544102
rect 237306 544046 237374 544102
rect 237430 544046 237498 544102
rect 237554 544046 237622 544102
rect 237678 544046 255250 544102
rect 255306 544046 255374 544102
rect 255430 544046 255498 544102
rect 255554 544046 255622 544102
rect 255678 544046 273250 544102
rect 273306 544046 273374 544102
rect 273430 544046 273498 544102
rect 273554 544046 273622 544102
rect 273678 544046 291250 544102
rect 291306 544046 291374 544102
rect 291430 544046 291498 544102
rect 291554 544046 291622 544102
rect 291678 544046 309250 544102
rect 309306 544046 309374 544102
rect 309430 544046 309498 544102
rect 309554 544046 309622 544102
rect 309678 544046 327250 544102
rect 327306 544046 327374 544102
rect 327430 544046 327498 544102
rect 327554 544046 327622 544102
rect 327678 544046 345250 544102
rect 345306 544046 345374 544102
rect 345430 544046 345498 544102
rect 345554 544046 345622 544102
rect 345678 544046 363250 544102
rect 363306 544046 363374 544102
rect 363430 544046 363498 544102
rect 363554 544046 363622 544102
rect 363678 544046 381250 544102
rect 381306 544046 381374 544102
rect 381430 544046 381498 544102
rect 381554 544046 381622 544102
rect 381678 544046 399250 544102
rect 399306 544046 399374 544102
rect 399430 544046 399498 544102
rect 399554 544046 399622 544102
rect 399678 544046 417250 544102
rect 417306 544046 417374 544102
rect 417430 544046 417498 544102
rect 417554 544046 417622 544102
rect 417678 544046 435250 544102
rect 435306 544046 435374 544102
rect 435430 544046 435498 544102
rect 435554 544046 435622 544102
rect 435678 544046 453250 544102
rect 453306 544046 453374 544102
rect 453430 544046 453498 544102
rect 453554 544046 453622 544102
rect 453678 544046 471250 544102
rect 471306 544046 471374 544102
rect 471430 544046 471498 544102
rect 471554 544046 471622 544102
rect 471678 544046 489250 544102
rect 489306 544046 489374 544102
rect 489430 544046 489498 544102
rect 489554 544046 489622 544102
rect 489678 544046 507250 544102
rect 507306 544046 507374 544102
rect 507430 544046 507498 544102
rect 507554 544046 507622 544102
rect 507678 544046 525250 544102
rect 525306 544046 525374 544102
rect 525430 544046 525498 544102
rect 525554 544046 525622 544102
rect 525678 544046 543250 544102
rect 543306 544046 543374 544102
rect 543430 544046 543498 544102
rect 543554 544046 543622 544102
rect 543678 544046 561250 544102
rect 561306 544046 561374 544102
rect 561430 544046 561498 544102
rect 561554 544046 561622 544102
rect 561678 544046 579250 544102
rect 579306 544046 579374 544102
rect 579430 544046 579498 544102
rect 579554 544046 579622 544102
rect 579678 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 3250 543978
rect 3306 543922 3374 543978
rect 3430 543922 3498 543978
rect 3554 543922 3622 543978
rect 3678 543922 21250 543978
rect 21306 543922 21374 543978
rect 21430 543922 21498 543978
rect 21554 543922 21622 543978
rect 21678 543922 39250 543978
rect 39306 543922 39374 543978
rect 39430 543922 39498 543978
rect 39554 543922 39622 543978
rect 39678 543922 57250 543978
rect 57306 543922 57374 543978
rect 57430 543922 57498 543978
rect 57554 543922 57622 543978
rect 57678 543922 75250 543978
rect 75306 543922 75374 543978
rect 75430 543922 75498 543978
rect 75554 543922 75622 543978
rect 75678 543922 93250 543978
rect 93306 543922 93374 543978
rect 93430 543922 93498 543978
rect 93554 543922 93622 543978
rect 93678 543922 111250 543978
rect 111306 543922 111374 543978
rect 111430 543922 111498 543978
rect 111554 543922 111622 543978
rect 111678 543922 129250 543978
rect 129306 543922 129374 543978
rect 129430 543922 129498 543978
rect 129554 543922 129622 543978
rect 129678 543922 147250 543978
rect 147306 543922 147374 543978
rect 147430 543922 147498 543978
rect 147554 543922 147622 543978
rect 147678 543922 165250 543978
rect 165306 543922 165374 543978
rect 165430 543922 165498 543978
rect 165554 543922 165622 543978
rect 165678 543922 183250 543978
rect 183306 543922 183374 543978
rect 183430 543922 183498 543978
rect 183554 543922 183622 543978
rect 183678 543922 201250 543978
rect 201306 543922 201374 543978
rect 201430 543922 201498 543978
rect 201554 543922 201622 543978
rect 201678 543922 219250 543978
rect 219306 543922 219374 543978
rect 219430 543922 219498 543978
rect 219554 543922 219622 543978
rect 219678 543922 237250 543978
rect 237306 543922 237374 543978
rect 237430 543922 237498 543978
rect 237554 543922 237622 543978
rect 237678 543922 255250 543978
rect 255306 543922 255374 543978
rect 255430 543922 255498 543978
rect 255554 543922 255622 543978
rect 255678 543922 273250 543978
rect 273306 543922 273374 543978
rect 273430 543922 273498 543978
rect 273554 543922 273622 543978
rect 273678 543922 291250 543978
rect 291306 543922 291374 543978
rect 291430 543922 291498 543978
rect 291554 543922 291622 543978
rect 291678 543922 309250 543978
rect 309306 543922 309374 543978
rect 309430 543922 309498 543978
rect 309554 543922 309622 543978
rect 309678 543922 327250 543978
rect 327306 543922 327374 543978
rect 327430 543922 327498 543978
rect 327554 543922 327622 543978
rect 327678 543922 345250 543978
rect 345306 543922 345374 543978
rect 345430 543922 345498 543978
rect 345554 543922 345622 543978
rect 345678 543922 363250 543978
rect 363306 543922 363374 543978
rect 363430 543922 363498 543978
rect 363554 543922 363622 543978
rect 363678 543922 381250 543978
rect 381306 543922 381374 543978
rect 381430 543922 381498 543978
rect 381554 543922 381622 543978
rect 381678 543922 399250 543978
rect 399306 543922 399374 543978
rect 399430 543922 399498 543978
rect 399554 543922 399622 543978
rect 399678 543922 417250 543978
rect 417306 543922 417374 543978
rect 417430 543922 417498 543978
rect 417554 543922 417622 543978
rect 417678 543922 435250 543978
rect 435306 543922 435374 543978
rect 435430 543922 435498 543978
rect 435554 543922 435622 543978
rect 435678 543922 453250 543978
rect 453306 543922 453374 543978
rect 453430 543922 453498 543978
rect 453554 543922 453622 543978
rect 453678 543922 471250 543978
rect 471306 543922 471374 543978
rect 471430 543922 471498 543978
rect 471554 543922 471622 543978
rect 471678 543922 489250 543978
rect 489306 543922 489374 543978
rect 489430 543922 489498 543978
rect 489554 543922 489622 543978
rect 489678 543922 507250 543978
rect 507306 543922 507374 543978
rect 507430 543922 507498 543978
rect 507554 543922 507622 543978
rect 507678 543922 525250 543978
rect 525306 543922 525374 543978
rect 525430 543922 525498 543978
rect 525554 543922 525622 543978
rect 525678 543922 543250 543978
rect 543306 543922 543374 543978
rect 543430 543922 543498 543978
rect 543554 543922 543622 543978
rect 543678 543922 561250 543978
rect 561306 543922 561374 543978
rect 561430 543922 561498 543978
rect 561554 543922 561622 543978
rect 561678 543922 579250 543978
rect 579306 543922 579374 543978
rect 579430 543922 579498 543978
rect 579554 543922 579622 543978
rect 579678 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 6970 532350
rect 7026 532294 7094 532350
rect 7150 532294 7218 532350
rect 7274 532294 7342 532350
rect 7398 532294 24970 532350
rect 25026 532294 25094 532350
rect 25150 532294 25218 532350
rect 25274 532294 25342 532350
rect 25398 532294 42970 532350
rect 43026 532294 43094 532350
rect 43150 532294 43218 532350
rect 43274 532294 43342 532350
rect 43398 532294 60970 532350
rect 61026 532294 61094 532350
rect 61150 532294 61218 532350
rect 61274 532294 61342 532350
rect 61398 532294 78970 532350
rect 79026 532294 79094 532350
rect 79150 532294 79218 532350
rect 79274 532294 79342 532350
rect 79398 532294 96970 532350
rect 97026 532294 97094 532350
rect 97150 532294 97218 532350
rect 97274 532294 97342 532350
rect 97398 532294 114970 532350
rect 115026 532294 115094 532350
rect 115150 532294 115218 532350
rect 115274 532294 115342 532350
rect 115398 532294 132970 532350
rect 133026 532294 133094 532350
rect 133150 532294 133218 532350
rect 133274 532294 133342 532350
rect 133398 532294 150970 532350
rect 151026 532294 151094 532350
rect 151150 532294 151218 532350
rect 151274 532294 151342 532350
rect 151398 532294 168970 532350
rect 169026 532294 169094 532350
rect 169150 532294 169218 532350
rect 169274 532294 169342 532350
rect 169398 532294 186970 532350
rect 187026 532294 187094 532350
rect 187150 532294 187218 532350
rect 187274 532294 187342 532350
rect 187398 532294 204970 532350
rect 205026 532294 205094 532350
rect 205150 532294 205218 532350
rect 205274 532294 205342 532350
rect 205398 532294 222970 532350
rect 223026 532294 223094 532350
rect 223150 532294 223218 532350
rect 223274 532294 223342 532350
rect 223398 532294 240970 532350
rect 241026 532294 241094 532350
rect 241150 532294 241218 532350
rect 241274 532294 241342 532350
rect 241398 532294 258970 532350
rect 259026 532294 259094 532350
rect 259150 532294 259218 532350
rect 259274 532294 259342 532350
rect 259398 532294 276970 532350
rect 277026 532294 277094 532350
rect 277150 532294 277218 532350
rect 277274 532294 277342 532350
rect 277398 532294 294970 532350
rect 295026 532294 295094 532350
rect 295150 532294 295218 532350
rect 295274 532294 295342 532350
rect 295398 532294 312970 532350
rect 313026 532294 313094 532350
rect 313150 532294 313218 532350
rect 313274 532294 313342 532350
rect 313398 532294 330970 532350
rect 331026 532294 331094 532350
rect 331150 532294 331218 532350
rect 331274 532294 331342 532350
rect 331398 532294 348970 532350
rect 349026 532294 349094 532350
rect 349150 532294 349218 532350
rect 349274 532294 349342 532350
rect 349398 532294 366970 532350
rect 367026 532294 367094 532350
rect 367150 532294 367218 532350
rect 367274 532294 367342 532350
rect 367398 532294 384970 532350
rect 385026 532294 385094 532350
rect 385150 532294 385218 532350
rect 385274 532294 385342 532350
rect 385398 532294 402970 532350
rect 403026 532294 403094 532350
rect 403150 532294 403218 532350
rect 403274 532294 403342 532350
rect 403398 532294 420970 532350
rect 421026 532294 421094 532350
rect 421150 532294 421218 532350
rect 421274 532294 421342 532350
rect 421398 532294 438970 532350
rect 439026 532294 439094 532350
rect 439150 532294 439218 532350
rect 439274 532294 439342 532350
rect 439398 532294 456970 532350
rect 457026 532294 457094 532350
rect 457150 532294 457218 532350
rect 457274 532294 457342 532350
rect 457398 532294 474970 532350
rect 475026 532294 475094 532350
rect 475150 532294 475218 532350
rect 475274 532294 475342 532350
rect 475398 532294 492970 532350
rect 493026 532294 493094 532350
rect 493150 532294 493218 532350
rect 493274 532294 493342 532350
rect 493398 532294 510970 532350
rect 511026 532294 511094 532350
rect 511150 532294 511218 532350
rect 511274 532294 511342 532350
rect 511398 532294 528970 532350
rect 529026 532294 529094 532350
rect 529150 532294 529218 532350
rect 529274 532294 529342 532350
rect 529398 532294 546970 532350
rect 547026 532294 547094 532350
rect 547150 532294 547218 532350
rect 547274 532294 547342 532350
rect 547398 532294 564970 532350
rect 565026 532294 565094 532350
rect 565150 532294 565218 532350
rect 565274 532294 565342 532350
rect 565398 532294 582970 532350
rect 583026 532294 583094 532350
rect 583150 532294 583218 532350
rect 583274 532294 583342 532350
rect 583398 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 6970 532226
rect 7026 532170 7094 532226
rect 7150 532170 7218 532226
rect 7274 532170 7342 532226
rect 7398 532170 24970 532226
rect 25026 532170 25094 532226
rect 25150 532170 25218 532226
rect 25274 532170 25342 532226
rect 25398 532170 42970 532226
rect 43026 532170 43094 532226
rect 43150 532170 43218 532226
rect 43274 532170 43342 532226
rect 43398 532170 60970 532226
rect 61026 532170 61094 532226
rect 61150 532170 61218 532226
rect 61274 532170 61342 532226
rect 61398 532170 78970 532226
rect 79026 532170 79094 532226
rect 79150 532170 79218 532226
rect 79274 532170 79342 532226
rect 79398 532170 96970 532226
rect 97026 532170 97094 532226
rect 97150 532170 97218 532226
rect 97274 532170 97342 532226
rect 97398 532170 114970 532226
rect 115026 532170 115094 532226
rect 115150 532170 115218 532226
rect 115274 532170 115342 532226
rect 115398 532170 132970 532226
rect 133026 532170 133094 532226
rect 133150 532170 133218 532226
rect 133274 532170 133342 532226
rect 133398 532170 150970 532226
rect 151026 532170 151094 532226
rect 151150 532170 151218 532226
rect 151274 532170 151342 532226
rect 151398 532170 168970 532226
rect 169026 532170 169094 532226
rect 169150 532170 169218 532226
rect 169274 532170 169342 532226
rect 169398 532170 186970 532226
rect 187026 532170 187094 532226
rect 187150 532170 187218 532226
rect 187274 532170 187342 532226
rect 187398 532170 204970 532226
rect 205026 532170 205094 532226
rect 205150 532170 205218 532226
rect 205274 532170 205342 532226
rect 205398 532170 222970 532226
rect 223026 532170 223094 532226
rect 223150 532170 223218 532226
rect 223274 532170 223342 532226
rect 223398 532170 240970 532226
rect 241026 532170 241094 532226
rect 241150 532170 241218 532226
rect 241274 532170 241342 532226
rect 241398 532170 258970 532226
rect 259026 532170 259094 532226
rect 259150 532170 259218 532226
rect 259274 532170 259342 532226
rect 259398 532170 276970 532226
rect 277026 532170 277094 532226
rect 277150 532170 277218 532226
rect 277274 532170 277342 532226
rect 277398 532170 294970 532226
rect 295026 532170 295094 532226
rect 295150 532170 295218 532226
rect 295274 532170 295342 532226
rect 295398 532170 312970 532226
rect 313026 532170 313094 532226
rect 313150 532170 313218 532226
rect 313274 532170 313342 532226
rect 313398 532170 330970 532226
rect 331026 532170 331094 532226
rect 331150 532170 331218 532226
rect 331274 532170 331342 532226
rect 331398 532170 348970 532226
rect 349026 532170 349094 532226
rect 349150 532170 349218 532226
rect 349274 532170 349342 532226
rect 349398 532170 366970 532226
rect 367026 532170 367094 532226
rect 367150 532170 367218 532226
rect 367274 532170 367342 532226
rect 367398 532170 384970 532226
rect 385026 532170 385094 532226
rect 385150 532170 385218 532226
rect 385274 532170 385342 532226
rect 385398 532170 402970 532226
rect 403026 532170 403094 532226
rect 403150 532170 403218 532226
rect 403274 532170 403342 532226
rect 403398 532170 420970 532226
rect 421026 532170 421094 532226
rect 421150 532170 421218 532226
rect 421274 532170 421342 532226
rect 421398 532170 438970 532226
rect 439026 532170 439094 532226
rect 439150 532170 439218 532226
rect 439274 532170 439342 532226
rect 439398 532170 456970 532226
rect 457026 532170 457094 532226
rect 457150 532170 457218 532226
rect 457274 532170 457342 532226
rect 457398 532170 474970 532226
rect 475026 532170 475094 532226
rect 475150 532170 475218 532226
rect 475274 532170 475342 532226
rect 475398 532170 492970 532226
rect 493026 532170 493094 532226
rect 493150 532170 493218 532226
rect 493274 532170 493342 532226
rect 493398 532170 510970 532226
rect 511026 532170 511094 532226
rect 511150 532170 511218 532226
rect 511274 532170 511342 532226
rect 511398 532170 528970 532226
rect 529026 532170 529094 532226
rect 529150 532170 529218 532226
rect 529274 532170 529342 532226
rect 529398 532170 546970 532226
rect 547026 532170 547094 532226
rect 547150 532170 547218 532226
rect 547274 532170 547342 532226
rect 547398 532170 564970 532226
rect 565026 532170 565094 532226
rect 565150 532170 565218 532226
rect 565274 532170 565342 532226
rect 565398 532170 582970 532226
rect 583026 532170 583094 532226
rect 583150 532170 583218 532226
rect 583274 532170 583342 532226
rect 583398 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 6970 532102
rect 7026 532046 7094 532102
rect 7150 532046 7218 532102
rect 7274 532046 7342 532102
rect 7398 532046 24970 532102
rect 25026 532046 25094 532102
rect 25150 532046 25218 532102
rect 25274 532046 25342 532102
rect 25398 532046 42970 532102
rect 43026 532046 43094 532102
rect 43150 532046 43218 532102
rect 43274 532046 43342 532102
rect 43398 532046 60970 532102
rect 61026 532046 61094 532102
rect 61150 532046 61218 532102
rect 61274 532046 61342 532102
rect 61398 532046 78970 532102
rect 79026 532046 79094 532102
rect 79150 532046 79218 532102
rect 79274 532046 79342 532102
rect 79398 532046 96970 532102
rect 97026 532046 97094 532102
rect 97150 532046 97218 532102
rect 97274 532046 97342 532102
rect 97398 532046 114970 532102
rect 115026 532046 115094 532102
rect 115150 532046 115218 532102
rect 115274 532046 115342 532102
rect 115398 532046 132970 532102
rect 133026 532046 133094 532102
rect 133150 532046 133218 532102
rect 133274 532046 133342 532102
rect 133398 532046 150970 532102
rect 151026 532046 151094 532102
rect 151150 532046 151218 532102
rect 151274 532046 151342 532102
rect 151398 532046 168970 532102
rect 169026 532046 169094 532102
rect 169150 532046 169218 532102
rect 169274 532046 169342 532102
rect 169398 532046 186970 532102
rect 187026 532046 187094 532102
rect 187150 532046 187218 532102
rect 187274 532046 187342 532102
rect 187398 532046 204970 532102
rect 205026 532046 205094 532102
rect 205150 532046 205218 532102
rect 205274 532046 205342 532102
rect 205398 532046 222970 532102
rect 223026 532046 223094 532102
rect 223150 532046 223218 532102
rect 223274 532046 223342 532102
rect 223398 532046 240970 532102
rect 241026 532046 241094 532102
rect 241150 532046 241218 532102
rect 241274 532046 241342 532102
rect 241398 532046 258970 532102
rect 259026 532046 259094 532102
rect 259150 532046 259218 532102
rect 259274 532046 259342 532102
rect 259398 532046 276970 532102
rect 277026 532046 277094 532102
rect 277150 532046 277218 532102
rect 277274 532046 277342 532102
rect 277398 532046 294970 532102
rect 295026 532046 295094 532102
rect 295150 532046 295218 532102
rect 295274 532046 295342 532102
rect 295398 532046 312970 532102
rect 313026 532046 313094 532102
rect 313150 532046 313218 532102
rect 313274 532046 313342 532102
rect 313398 532046 330970 532102
rect 331026 532046 331094 532102
rect 331150 532046 331218 532102
rect 331274 532046 331342 532102
rect 331398 532046 348970 532102
rect 349026 532046 349094 532102
rect 349150 532046 349218 532102
rect 349274 532046 349342 532102
rect 349398 532046 366970 532102
rect 367026 532046 367094 532102
rect 367150 532046 367218 532102
rect 367274 532046 367342 532102
rect 367398 532046 384970 532102
rect 385026 532046 385094 532102
rect 385150 532046 385218 532102
rect 385274 532046 385342 532102
rect 385398 532046 402970 532102
rect 403026 532046 403094 532102
rect 403150 532046 403218 532102
rect 403274 532046 403342 532102
rect 403398 532046 420970 532102
rect 421026 532046 421094 532102
rect 421150 532046 421218 532102
rect 421274 532046 421342 532102
rect 421398 532046 438970 532102
rect 439026 532046 439094 532102
rect 439150 532046 439218 532102
rect 439274 532046 439342 532102
rect 439398 532046 456970 532102
rect 457026 532046 457094 532102
rect 457150 532046 457218 532102
rect 457274 532046 457342 532102
rect 457398 532046 474970 532102
rect 475026 532046 475094 532102
rect 475150 532046 475218 532102
rect 475274 532046 475342 532102
rect 475398 532046 492970 532102
rect 493026 532046 493094 532102
rect 493150 532046 493218 532102
rect 493274 532046 493342 532102
rect 493398 532046 510970 532102
rect 511026 532046 511094 532102
rect 511150 532046 511218 532102
rect 511274 532046 511342 532102
rect 511398 532046 528970 532102
rect 529026 532046 529094 532102
rect 529150 532046 529218 532102
rect 529274 532046 529342 532102
rect 529398 532046 546970 532102
rect 547026 532046 547094 532102
rect 547150 532046 547218 532102
rect 547274 532046 547342 532102
rect 547398 532046 564970 532102
rect 565026 532046 565094 532102
rect 565150 532046 565218 532102
rect 565274 532046 565342 532102
rect 565398 532046 582970 532102
rect 583026 532046 583094 532102
rect 583150 532046 583218 532102
rect 583274 532046 583342 532102
rect 583398 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 6970 531978
rect 7026 531922 7094 531978
rect 7150 531922 7218 531978
rect 7274 531922 7342 531978
rect 7398 531922 24970 531978
rect 25026 531922 25094 531978
rect 25150 531922 25218 531978
rect 25274 531922 25342 531978
rect 25398 531922 42970 531978
rect 43026 531922 43094 531978
rect 43150 531922 43218 531978
rect 43274 531922 43342 531978
rect 43398 531922 60970 531978
rect 61026 531922 61094 531978
rect 61150 531922 61218 531978
rect 61274 531922 61342 531978
rect 61398 531922 78970 531978
rect 79026 531922 79094 531978
rect 79150 531922 79218 531978
rect 79274 531922 79342 531978
rect 79398 531922 96970 531978
rect 97026 531922 97094 531978
rect 97150 531922 97218 531978
rect 97274 531922 97342 531978
rect 97398 531922 114970 531978
rect 115026 531922 115094 531978
rect 115150 531922 115218 531978
rect 115274 531922 115342 531978
rect 115398 531922 132970 531978
rect 133026 531922 133094 531978
rect 133150 531922 133218 531978
rect 133274 531922 133342 531978
rect 133398 531922 150970 531978
rect 151026 531922 151094 531978
rect 151150 531922 151218 531978
rect 151274 531922 151342 531978
rect 151398 531922 168970 531978
rect 169026 531922 169094 531978
rect 169150 531922 169218 531978
rect 169274 531922 169342 531978
rect 169398 531922 186970 531978
rect 187026 531922 187094 531978
rect 187150 531922 187218 531978
rect 187274 531922 187342 531978
rect 187398 531922 204970 531978
rect 205026 531922 205094 531978
rect 205150 531922 205218 531978
rect 205274 531922 205342 531978
rect 205398 531922 222970 531978
rect 223026 531922 223094 531978
rect 223150 531922 223218 531978
rect 223274 531922 223342 531978
rect 223398 531922 240970 531978
rect 241026 531922 241094 531978
rect 241150 531922 241218 531978
rect 241274 531922 241342 531978
rect 241398 531922 258970 531978
rect 259026 531922 259094 531978
rect 259150 531922 259218 531978
rect 259274 531922 259342 531978
rect 259398 531922 276970 531978
rect 277026 531922 277094 531978
rect 277150 531922 277218 531978
rect 277274 531922 277342 531978
rect 277398 531922 294970 531978
rect 295026 531922 295094 531978
rect 295150 531922 295218 531978
rect 295274 531922 295342 531978
rect 295398 531922 312970 531978
rect 313026 531922 313094 531978
rect 313150 531922 313218 531978
rect 313274 531922 313342 531978
rect 313398 531922 330970 531978
rect 331026 531922 331094 531978
rect 331150 531922 331218 531978
rect 331274 531922 331342 531978
rect 331398 531922 348970 531978
rect 349026 531922 349094 531978
rect 349150 531922 349218 531978
rect 349274 531922 349342 531978
rect 349398 531922 366970 531978
rect 367026 531922 367094 531978
rect 367150 531922 367218 531978
rect 367274 531922 367342 531978
rect 367398 531922 384970 531978
rect 385026 531922 385094 531978
rect 385150 531922 385218 531978
rect 385274 531922 385342 531978
rect 385398 531922 402970 531978
rect 403026 531922 403094 531978
rect 403150 531922 403218 531978
rect 403274 531922 403342 531978
rect 403398 531922 420970 531978
rect 421026 531922 421094 531978
rect 421150 531922 421218 531978
rect 421274 531922 421342 531978
rect 421398 531922 438970 531978
rect 439026 531922 439094 531978
rect 439150 531922 439218 531978
rect 439274 531922 439342 531978
rect 439398 531922 456970 531978
rect 457026 531922 457094 531978
rect 457150 531922 457218 531978
rect 457274 531922 457342 531978
rect 457398 531922 474970 531978
rect 475026 531922 475094 531978
rect 475150 531922 475218 531978
rect 475274 531922 475342 531978
rect 475398 531922 492970 531978
rect 493026 531922 493094 531978
rect 493150 531922 493218 531978
rect 493274 531922 493342 531978
rect 493398 531922 510970 531978
rect 511026 531922 511094 531978
rect 511150 531922 511218 531978
rect 511274 531922 511342 531978
rect 511398 531922 528970 531978
rect 529026 531922 529094 531978
rect 529150 531922 529218 531978
rect 529274 531922 529342 531978
rect 529398 531922 546970 531978
rect 547026 531922 547094 531978
rect 547150 531922 547218 531978
rect 547274 531922 547342 531978
rect 547398 531922 564970 531978
rect 565026 531922 565094 531978
rect 565150 531922 565218 531978
rect 565274 531922 565342 531978
rect 565398 531922 582970 531978
rect 583026 531922 583094 531978
rect 583150 531922 583218 531978
rect 583274 531922 583342 531978
rect 583398 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 3250 526350
rect 3306 526294 3374 526350
rect 3430 526294 3498 526350
rect 3554 526294 3622 526350
rect 3678 526294 21250 526350
rect 21306 526294 21374 526350
rect 21430 526294 21498 526350
rect 21554 526294 21622 526350
rect 21678 526294 39250 526350
rect 39306 526294 39374 526350
rect 39430 526294 39498 526350
rect 39554 526294 39622 526350
rect 39678 526294 57250 526350
rect 57306 526294 57374 526350
rect 57430 526294 57498 526350
rect 57554 526294 57622 526350
rect 57678 526294 75250 526350
rect 75306 526294 75374 526350
rect 75430 526294 75498 526350
rect 75554 526294 75622 526350
rect 75678 526294 93250 526350
rect 93306 526294 93374 526350
rect 93430 526294 93498 526350
rect 93554 526294 93622 526350
rect 93678 526294 111250 526350
rect 111306 526294 111374 526350
rect 111430 526294 111498 526350
rect 111554 526294 111622 526350
rect 111678 526294 129250 526350
rect 129306 526294 129374 526350
rect 129430 526294 129498 526350
rect 129554 526294 129622 526350
rect 129678 526294 147250 526350
rect 147306 526294 147374 526350
rect 147430 526294 147498 526350
rect 147554 526294 147622 526350
rect 147678 526294 165250 526350
rect 165306 526294 165374 526350
rect 165430 526294 165498 526350
rect 165554 526294 165622 526350
rect 165678 526294 183250 526350
rect 183306 526294 183374 526350
rect 183430 526294 183498 526350
rect 183554 526294 183622 526350
rect 183678 526294 201250 526350
rect 201306 526294 201374 526350
rect 201430 526294 201498 526350
rect 201554 526294 201622 526350
rect 201678 526294 219250 526350
rect 219306 526294 219374 526350
rect 219430 526294 219498 526350
rect 219554 526294 219622 526350
rect 219678 526294 237250 526350
rect 237306 526294 237374 526350
rect 237430 526294 237498 526350
rect 237554 526294 237622 526350
rect 237678 526294 255250 526350
rect 255306 526294 255374 526350
rect 255430 526294 255498 526350
rect 255554 526294 255622 526350
rect 255678 526294 273250 526350
rect 273306 526294 273374 526350
rect 273430 526294 273498 526350
rect 273554 526294 273622 526350
rect 273678 526294 291250 526350
rect 291306 526294 291374 526350
rect 291430 526294 291498 526350
rect 291554 526294 291622 526350
rect 291678 526294 309250 526350
rect 309306 526294 309374 526350
rect 309430 526294 309498 526350
rect 309554 526294 309622 526350
rect 309678 526294 327250 526350
rect 327306 526294 327374 526350
rect 327430 526294 327498 526350
rect 327554 526294 327622 526350
rect 327678 526294 345250 526350
rect 345306 526294 345374 526350
rect 345430 526294 345498 526350
rect 345554 526294 345622 526350
rect 345678 526294 363250 526350
rect 363306 526294 363374 526350
rect 363430 526294 363498 526350
rect 363554 526294 363622 526350
rect 363678 526294 381250 526350
rect 381306 526294 381374 526350
rect 381430 526294 381498 526350
rect 381554 526294 381622 526350
rect 381678 526294 399250 526350
rect 399306 526294 399374 526350
rect 399430 526294 399498 526350
rect 399554 526294 399622 526350
rect 399678 526294 417250 526350
rect 417306 526294 417374 526350
rect 417430 526294 417498 526350
rect 417554 526294 417622 526350
rect 417678 526294 435250 526350
rect 435306 526294 435374 526350
rect 435430 526294 435498 526350
rect 435554 526294 435622 526350
rect 435678 526294 453250 526350
rect 453306 526294 453374 526350
rect 453430 526294 453498 526350
rect 453554 526294 453622 526350
rect 453678 526294 471250 526350
rect 471306 526294 471374 526350
rect 471430 526294 471498 526350
rect 471554 526294 471622 526350
rect 471678 526294 489250 526350
rect 489306 526294 489374 526350
rect 489430 526294 489498 526350
rect 489554 526294 489622 526350
rect 489678 526294 507250 526350
rect 507306 526294 507374 526350
rect 507430 526294 507498 526350
rect 507554 526294 507622 526350
rect 507678 526294 525250 526350
rect 525306 526294 525374 526350
rect 525430 526294 525498 526350
rect 525554 526294 525622 526350
rect 525678 526294 543250 526350
rect 543306 526294 543374 526350
rect 543430 526294 543498 526350
rect 543554 526294 543622 526350
rect 543678 526294 561250 526350
rect 561306 526294 561374 526350
rect 561430 526294 561498 526350
rect 561554 526294 561622 526350
rect 561678 526294 579250 526350
rect 579306 526294 579374 526350
rect 579430 526294 579498 526350
rect 579554 526294 579622 526350
rect 579678 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 3250 526226
rect 3306 526170 3374 526226
rect 3430 526170 3498 526226
rect 3554 526170 3622 526226
rect 3678 526170 21250 526226
rect 21306 526170 21374 526226
rect 21430 526170 21498 526226
rect 21554 526170 21622 526226
rect 21678 526170 39250 526226
rect 39306 526170 39374 526226
rect 39430 526170 39498 526226
rect 39554 526170 39622 526226
rect 39678 526170 57250 526226
rect 57306 526170 57374 526226
rect 57430 526170 57498 526226
rect 57554 526170 57622 526226
rect 57678 526170 75250 526226
rect 75306 526170 75374 526226
rect 75430 526170 75498 526226
rect 75554 526170 75622 526226
rect 75678 526170 93250 526226
rect 93306 526170 93374 526226
rect 93430 526170 93498 526226
rect 93554 526170 93622 526226
rect 93678 526170 111250 526226
rect 111306 526170 111374 526226
rect 111430 526170 111498 526226
rect 111554 526170 111622 526226
rect 111678 526170 129250 526226
rect 129306 526170 129374 526226
rect 129430 526170 129498 526226
rect 129554 526170 129622 526226
rect 129678 526170 147250 526226
rect 147306 526170 147374 526226
rect 147430 526170 147498 526226
rect 147554 526170 147622 526226
rect 147678 526170 165250 526226
rect 165306 526170 165374 526226
rect 165430 526170 165498 526226
rect 165554 526170 165622 526226
rect 165678 526170 183250 526226
rect 183306 526170 183374 526226
rect 183430 526170 183498 526226
rect 183554 526170 183622 526226
rect 183678 526170 201250 526226
rect 201306 526170 201374 526226
rect 201430 526170 201498 526226
rect 201554 526170 201622 526226
rect 201678 526170 219250 526226
rect 219306 526170 219374 526226
rect 219430 526170 219498 526226
rect 219554 526170 219622 526226
rect 219678 526170 237250 526226
rect 237306 526170 237374 526226
rect 237430 526170 237498 526226
rect 237554 526170 237622 526226
rect 237678 526170 255250 526226
rect 255306 526170 255374 526226
rect 255430 526170 255498 526226
rect 255554 526170 255622 526226
rect 255678 526170 273250 526226
rect 273306 526170 273374 526226
rect 273430 526170 273498 526226
rect 273554 526170 273622 526226
rect 273678 526170 291250 526226
rect 291306 526170 291374 526226
rect 291430 526170 291498 526226
rect 291554 526170 291622 526226
rect 291678 526170 309250 526226
rect 309306 526170 309374 526226
rect 309430 526170 309498 526226
rect 309554 526170 309622 526226
rect 309678 526170 327250 526226
rect 327306 526170 327374 526226
rect 327430 526170 327498 526226
rect 327554 526170 327622 526226
rect 327678 526170 345250 526226
rect 345306 526170 345374 526226
rect 345430 526170 345498 526226
rect 345554 526170 345622 526226
rect 345678 526170 363250 526226
rect 363306 526170 363374 526226
rect 363430 526170 363498 526226
rect 363554 526170 363622 526226
rect 363678 526170 381250 526226
rect 381306 526170 381374 526226
rect 381430 526170 381498 526226
rect 381554 526170 381622 526226
rect 381678 526170 399250 526226
rect 399306 526170 399374 526226
rect 399430 526170 399498 526226
rect 399554 526170 399622 526226
rect 399678 526170 417250 526226
rect 417306 526170 417374 526226
rect 417430 526170 417498 526226
rect 417554 526170 417622 526226
rect 417678 526170 435250 526226
rect 435306 526170 435374 526226
rect 435430 526170 435498 526226
rect 435554 526170 435622 526226
rect 435678 526170 453250 526226
rect 453306 526170 453374 526226
rect 453430 526170 453498 526226
rect 453554 526170 453622 526226
rect 453678 526170 471250 526226
rect 471306 526170 471374 526226
rect 471430 526170 471498 526226
rect 471554 526170 471622 526226
rect 471678 526170 489250 526226
rect 489306 526170 489374 526226
rect 489430 526170 489498 526226
rect 489554 526170 489622 526226
rect 489678 526170 507250 526226
rect 507306 526170 507374 526226
rect 507430 526170 507498 526226
rect 507554 526170 507622 526226
rect 507678 526170 525250 526226
rect 525306 526170 525374 526226
rect 525430 526170 525498 526226
rect 525554 526170 525622 526226
rect 525678 526170 543250 526226
rect 543306 526170 543374 526226
rect 543430 526170 543498 526226
rect 543554 526170 543622 526226
rect 543678 526170 561250 526226
rect 561306 526170 561374 526226
rect 561430 526170 561498 526226
rect 561554 526170 561622 526226
rect 561678 526170 579250 526226
rect 579306 526170 579374 526226
rect 579430 526170 579498 526226
rect 579554 526170 579622 526226
rect 579678 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 3250 526102
rect 3306 526046 3374 526102
rect 3430 526046 3498 526102
rect 3554 526046 3622 526102
rect 3678 526046 21250 526102
rect 21306 526046 21374 526102
rect 21430 526046 21498 526102
rect 21554 526046 21622 526102
rect 21678 526046 39250 526102
rect 39306 526046 39374 526102
rect 39430 526046 39498 526102
rect 39554 526046 39622 526102
rect 39678 526046 57250 526102
rect 57306 526046 57374 526102
rect 57430 526046 57498 526102
rect 57554 526046 57622 526102
rect 57678 526046 75250 526102
rect 75306 526046 75374 526102
rect 75430 526046 75498 526102
rect 75554 526046 75622 526102
rect 75678 526046 93250 526102
rect 93306 526046 93374 526102
rect 93430 526046 93498 526102
rect 93554 526046 93622 526102
rect 93678 526046 111250 526102
rect 111306 526046 111374 526102
rect 111430 526046 111498 526102
rect 111554 526046 111622 526102
rect 111678 526046 129250 526102
rect 129306 526046 129374 526102
rect 129430 526046 129498 526102
rect 129554 526046 129622 526102
rect 129678 526046 147250 526102
rect 147306 526046 147374 526102
rect 147430 526046 147498 526102
rect 147554 526046 147622 526102
rect 147678 526046 165250 526102
rect 165306 526046 165374 526102
rect 165430 526046 165498 526102
rect 165554 526046 165622 526102
rect 165678 526046 183250 526102
rect 183306 526046 183374 526102
rect 183430 526046 183498 526102
rect 183554 526046 183622 526102
rect 183678 526046 201250 526102
rect 201306 526046 201374 526102
rect 201430 526046 201498 526102
rect 201554 526046 201622 526102
rect 201678 526046 219250 526102
rect 219306 526046 219374 526102
rect 219430 526046 219498 526102
rect 219554 526046 219622 526102
rect 219678 526046 237250 526102
rect 237306 526046 237374 526102
rect 237430 526046 237498 526102
rect 237554 526046 237622 526102
rect 237678 526046 255250 526102
rect 255306 526046 255374 526102
rect 255430 526046 255498 526102
rect 255554 526046 255622 526102
rect 255678 526046 273250 526102
rect 273306 526046 273374 526102
rect 273430 526046 273498 526102
rect 273554 526046 273622 526102
rect 273678 526046 291250 526102
rect 291306 526046 291374 526102
rect 291430 526046 291498 526102
rect 291554 526046 291622 526102
rect 291678 526046 309250 526102
rect 309306 526046 309374 526102
rect 309430 526046 309498 526102
rect 309554 526046 309622 526102
rect 309678 526046 327250 526102
rect 327306 526046 327374 526102
rect 327430 526046 327498 526102
rect 327554 526046 327622 526102
rect 327678 526046 345250 526102
rect 345306 526046 345374 526102
rect 345430 526046 345498 526102
rect 345554 526046 345622 526102
rect 345678 526046 363250 526102
rect 363306 526046 363374 526102
rect 363430 526046 363498 526102
rect 363554 526046 363622 526102
rect 363678 526046 381250 526102
rect 381306 526046 381374 526102
rect 381430 526046 381498 526102
rect 381554 526046 381622 526102
rect 381678 526046 399250 526102
rect 399306 526046 399374 526102
rect 399430 526046 399498 526102
rect 399554 526046 399622 526102
rect 399678 526046 417250 526102
rect 417306 526046 417374 526102
rect 417430 526046 417498 526102
rect 417554 526046 417622 526102
rect 417678 526046 435250 526102
rect 435306 526046 435374 526102
rect 435430 526046 435498 526102
rect 435554 526046 435622 526102
rect 435678 526046 453250 526102
rect 453306 526046 453374 526102
rect 453430 526046 453498 526102
rect 453554 526046 453622 526102
rect 453678 526046 471250 526102
rect 471306 526046 471374 526102
rect 471430 526046 471498 526102
rect 471554 526046 471622 526102
rect 471678 526046 489250 526102
rect 489306 526046 489374 526102
rect 489430 526046 489498 526102
rect 489554 526046 489622 526102
rect 489678 526046 507250 526102
rect 507306 526046 507374 526102
rect 507430 526046 507498 526102
rect 507554 526046 507622 526102
rect 507678 526046 525250 526102
rect 525306 526046 525374 526102
rect 525430 526046 525498 526102
rect 525554 526046 525622 526102
rect 525678 526046 543250 526102
rect 543306 526046 543374 526102
rect 543430 526046 543498 526102
rect 543554 526046 543622 526102
rect 543678 526046 561250 526102
rect 561306 526046 561374 526102
rect 561430 526046 561498 526102
rect 561554 526046 561622 526102
rect 561678 526046 579250 526102
rect 579306 526046 579374 526102
rect 579430 526046 579498 526102
rect 579554 526046 579622 526102
rect 579678 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 3250 525978
rect 3306 525922 3374 525978
rect 3430 525922 3498 525978
rect 3554 525922 3622 525978
rect 3678 525922 21250 525978
rect 21306 525922 21374 525978
rect 21430 525922 21498 525978
rect 21554 525922 21622 525978
rect 21678 525922 39250 525978
rect 39306 525922 39374 525978
rect 39430 525922 39498 525978
rect 39554 525922 39622 525978
rect 39678 525922 57250 525978
rect 57306 525922 57374 525978
rect 57430 525922 57498 525978
rect 57554 525922 57622 525978
rect 57678 525922 75250 525978
rect 75306 525922 75374 525978
rect 75430 525922 75498 525978
rect 75554 525922 75622 525978
rect 75678 525922 93250 525978
rect 93306 525922 93374 525978
rect 93430 525922 93498 525978
rect 93554 525922 93622 525978
rect 93678 525922 111250 525978
rect 111306 525922 111374 525978
rect 111430 525922 111498 525978
rect 111554 525922 111622 525978
rect 111678 525922 129250 525978
rect 129306 525922 129374 525978
rect 129430 525922 129498 525978
rect 129554 525922 129622 525978
rect 129678 525922 147250 525978
rect 147306 525922 147374 525978
rect 147430 525922 147498 525978
rect 147554 525922 147622 525978
rect 147678 525922 165250 525978
rect 165306 525922 165374 525978
rect 165430 525922 165498 525978
rect 165554 525922 165622 525978
rect 165678 525922 183250 525978
rect 183306 525922 183374 525978
rect 183430 525922 183498 525978
rect 183554 525922 183622 525978
rect 183678 525922 201250 525978
rect 201306 525922 201374 525978
rect 201430 525922 201498 525978
rect 201554 525922 201622 525978
rect 201678 525922 219250 525978
rect 219306 525922 219374 525978
rect 219430 525922 219498 525978
rect 219554 525922 219622 525978
rect 219678 525922 237250 525978
rect 237306 525922 237374 525978
rect 237430 525922 237498 525978
rect 237554 525922 237622 525978
rect 237678 525922 255250 525978
rect 255306 525922 255374 525978
rect 255430 525922 255498 525978
rect 255554 525922 255622 525978
rect 255678 525922 273250 525978
rect 273306 525922 273374 525978
rect 273430 525922 273498 525978
rect 273554 525922 273622 525978
rect 273678 525922 291250 525978
rect 291306 525922 291374 525978
rect 291430 525922 291498 525978
rect 291554 525922 291622 525978
rect 291678 525922 309250 525978
rect 309306 525922 309374 525978
rect 309430 525922 309498 525978
rect 309554 525922 309622 525978
rect 309678 525922 327250 525978
rect 327306 525922 327374 525978
rect 327430 525922 327498 525978
rect 327554 525922 327622 525978
rect 327678 525922 345250 525978
rect 345306 525922 345374 525978
rect 345430 525922 345498 525978
rect 345554 525922 345622 525978
rect 345678 525922 363250 525978
rect 363306 525922 363374 525978
rect 363430 525922 363498 525978
rect 363554 525922 363622 525978
rect 363678 525922 381250 525978
rect 381306 525922 381374 525978
rect 381430 525922 381498 525978
rect 381554 525922 381622 525978
rect 381678 525922 399250 525978
rect 399306 525922 399374 525978
rect 399430 525922 399498 525978
rect 399554 525922 399622 525978
rect 399678 525922 417250 525978
rect 417306 525922 417374 525978
rect 417430 525922 417498 525978
rect 417554 525922 417622 525978
rect 417678 525922 435250 525978
rect 435306 525922 435374 525978
rect 435430 525922 435498 525978
rect 435554 525922 435622 525978
rect 435678 525922 453250 525978
rect 453306 525922 453374 525978
rect 453430 525922 453498 525978
rect 453554 525922 453622 525978
rect 453678 525922 471250 525978
rect 471306 525922 471374 525978
rect 471430 525922 471498 525978
rect 471554 525922 471622 525978
rect 471678 525922 489250 525978
rect 489306 525922 489374 525978
rect 489430 525922 489498 525978
rect 489554 525922 489622 525978
rect 489678 525922 507250 525978
rect 507306 525922 507374 525978
rect 507430 525922 507498 525978
rect 507554 525922 507622 525978
rect 507678 525922 525250 525978
rect 525306 525922 525374 525978
rect 525430 525922 525498 525978
rect 525554 525922 525622 525978
rect 525678 525922 543250 525978
rect 543306 525922 543374 525978
rect 543430 525922 543498 525978
rect 543554 525922 543622 525978
rect 543678 525922 561250 525978
rect 561306 525922 561374 525978
rect 561430 525922 561498 525978
rect 561554 525922 561622 525978
rect 561678 525922 579250 525978
rect 579306 525922 579374 525978
rect 579430 525922 579498 525978
rect 579554 525922 579622 525978
rect 579678 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 6970 514350
rect 7026 514294 7094 514350
rect 7150 514294 7218 514350
rect 7274 514294 7342 514350
rect 7398 514294 24970 514350
rect 25026 514294 25094 514350
rect 25150 514294 25218 514350
rect 25274 514294 25342 514350
rect 25398 514294 42970 514350
rect 43026 514294 43094 514350
rect 43150 514294 43218 514350
rect 43274 514294 43342 514350
rect 43398 514294 60970 514350
rect 61026 514294 61094 514350
rect 61150 514294 61218 514350
rect 61274 514294 61342 514350
rect 61398 514294 78970 514350
rect 79026 514294 79094 514350
rect 79150 514294 79218 514350
rect 79274 514294 79342 514350
rect 79398 514294 96970 514350
rect 97026 514294 97094 514350
rect 97150 514294 97218 514350
rect 97274 514294 97342 514350
rect 97398 514294 114970 514350
rect 115026 514294 115094 514350
rect 115150 514294 115218 514350
rect 115274 514294 115342 514350
rect 115398 514294 132970 514350
rect 133026 514294 133094 514350
rect 133150 514294 133218 514350
rect 133274 514294 133342 514350
rect 133398 514294 150970 514350
rect 151026 514294 151094 514350
rect 151150 514294 151218 514350
rect 151274 514294 151342 514350
rect 151398 514294 168970 514350
rect 169026 514294 169094 514350
rect 169150 514294 169218 514350
rect 169274 514294 169342 514350
rect 169398 514294 186970 514350
rect 187026 514294 187094 514350
rect 187150 514294 187218 514350
rect 187274 514294 187342 514350
rect 187398 514294 204970 514350
rect 205026 514294 205094 514350
rect 205150 514294 205218 514350
rect 205274 514294 205342 514350
rect 205398 514294 222970 514350
rect 223026 514294 223094 514350
rect 223150 514294 223218 514350
rect 223274 514294 223342 514350
rect 223398 514294 240970 514350
rect 241026 514294 241094 514350
rect 241150 514294 241218 514350
rect 241274 514294 241342 514350
rect 241398 514294 258970 514350
rect 259026 514294 259094 514350
rect 259150 514294 259218 514350
rect 259274 514294 259342 514350
rect 259398 514294 276970 514350
rect 277026 514294 277094 514350
rect 277150 514294 277218 514350
rect 277274 514294 277342 514350
rect 277398 514294 294970 514350
rect 295026 514294 295094 514350
rect 295150 514294 295218 514350
rect 295274 514294 295342 514350
rect 295398 514294 312970 514350
rect 313026 514294 313094 514350
rect 313150 514294 313218 514350
rect 313274 514294 313342 514350
rect 313398 514294 330970 514350
rect 331026 514294 331094 514350
rect 331150 514294 331218 514350
rect 331274 514294 331342 514350
rect 331398 514294 348970 514350
rect 349026 514294 349094 514350
rect 349150 514294 349218 514350
rect 349274 514294 349342 514350
rect 349398 514294 366970 514350
rect 367026 514294 367094 514350
rect 367150 514294 367218 514350
rect 367274 514294 367342 514350
rect 367398 514294 384970 514350
rect 385026 514294 385094 514350
rect 385150 514294 385218 514350
rect 385274 514294 385342 514350
rect 385398 514294 402970 514350
rect 403026 514294 403094 514350
rect 403150 514294 403218 514350
rect 403274 514294 403342 514350
rect 403398 514294 420970 514350
rect 421026 514294 421094 514350
rect 421150 514294 421218 514350
rect 421274 514294 421342 514350
rect 421398 514294 438970 514350
rect 439026 514294 439094 514350
rect 439150 514294 439218 514350
rect 439274 514294 439342 514350
rect 439398 514294 456970 514350
rect 457026 514294 457094 514350
rect 457150 514294 457218 514350
rect 457274 514294 457342 514350
rect 457398 514294 474970 514350
rect 475026 514294 475094 514350
rect 475150 514294 475218 514350
rect 475274 514294 475342 514350
rect 475398 514294 492970 514350
rect 493026 514294 493094 514350
rect 493150 514294 493218 514350
rect 493274 514294 493342 514350
rect 493398 514294 510970 514350
rect 511026 514294 511094 514350
rect 511150 514294 511218 514350
rect 511274 514294 511342 514350
rect 511398 514294 528970 514350
rect 529026 514294 529094 514350
rect 529150 514294 529218 514350
rect 529274 514294 529342 514350
rect 529398 514294 546970 514350
rect 547026 514294 547094 514350
rect 547150 514294 547218 514350
rect 547274 514294 547342 514350
rect 547398 514294 564970 514350
rect 565026 514294 565094 514350
rect 565150 514294 565218 514350
rect 565274 514294 565342 514350
rect 565398 514294 582970 514350
rect 583026 514294 583094 514350
rect 583150 514294 583218 514350
rect 583274 514294 583342 514350
rect 583398 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 6970 514226
rect 7026 514170 7094 514226
rect 7150 514170 7218 514226
rect 7274 514170 7342 514226
rect 7398 514170 24970 514226
rect 25026 514170 25094 514226
rect 25150 514170 25218 514226
rect 25274 514170 25342 514226
rect 25398 514170 42970 514226
rect 43026 514170 43094 514226
rect 43150 514170 43218 514226
rect 43274 514170 43342 514226
rect 43398 514170 60970 514226
rect 61026 514170 61094 514226
rect 61150 514170 61218 514226
rect 61274 514170 61342 514226
rect 61398 514170 78970 514226
rect 79026 514170 79094 514226
rect 79150 514170 79218 514226
rect 79274 514170 79342 514226
rect 79398 514170 96970 514226
rect 97026 514170 97094 514226
rect 97150 514170 97218 514226
rect 97274 514170 97342 514226
rect 97398 514170 114970 514226
rect 115026 514170 115094 514226
rect 115150 514170 115218 514226
rect 115274 514170 115342 514226
rect 115398 514170 132970 514226
rect 133026 514170 133094 514226
rect 133150 514170 133218 514226
rect 133274 514170 133342 514226
rect 133398 514170 150970 514226
rect 151026 514170 151094 514226
rect 151150 514170 151218 514226
rect 151274 514170 151342 514226
rect 151398 514170 168970 514226
rect 169026 514170 169094 514226
rect 169150 514170 169218 514226
rect 169274 514170 169342 514226
rect 169398 514170 186970 514226
rect 187026 514170 187094 514226
rect 187150 514170 187218 514226
rect 187274 514170 187342 514226
rect 187398 514170 204970 514226
rect 205026 514170 205094 514226
rect 205150 514170 205218 514226
rect 205274 514170 205342 514226
rect 205398 514170 222970 514226
rect 223026 514170 223094 514226
rect 223150 514170 223218 514226
rect 223274 514170 223342 514226
rect 223398 514170 240970 514226
rect 241026 514170 241094 514226
rect 241150 514170 241218 514226
rect 241274 514170 241342 514226
rect 241398 514170 258970 514226
rect 259026 514170 259094 514226
rect 259150 514170 259218 514226
rect 259274 514170 259342 514226
rect 259398 514170 276970 514226
rect 277026 514170 277094 514226
rect 277150 514170 277218 514226
rect 277274 514170 277342 514226
rect 277398 514170 294970 514226
rect 295026 514170 295094 514226
rect 295150 514170 295218 514226
rect 295274 514170 295342 514226
rect 295398 514170 312970 514226
rect 313026 514170 313094 514226
rect 313150 514170 313218 514226
rect 313274 514170 313342 514226
rect 313398 514170 330970 514226
rect 331026 514170 331094 514226
rect 331150 514170 331218 514226
rect 331274 514170 331342 514226
rect 331398 514170 348970 514226
rect 349026 514170 349094 514226
rect 349150 514170 349218 514226
rect 349274 514170 349342 514226
rect 349398 514170 366970 514226
rect 367026 514170 367094 514226
rect 367150 514170 367218 514226
rect 367274 514170 367342 514226
rect 367398 514170 384970 514226
rect 385026 514170 385094 514226
rect 385150 514170 385218 514226
rect 385274 514170 385342 514226
rect 385398 514170 402970 514226
rect 403026 514170 403094 514226
rect 403150 514170 403218 514226
rect 403274 514170 403342 514226
rect 403398 514170 420970 514226
rect 421026 514170 421094 514226
rect 421150 514170 421218 514226
rect 421274 514170 421342 514226
rect 421398 514170 438970 514226
rect 439026 514170 439094 514226
rect 439150 514170 439218 514226
rect 439274 514170 439342 514226
rect 439398 514170 456970 514226
rect 457026 514170 457094 514226
rect 457150 514170 457218 514226
rect 457274 514170 457342 514226
rect 457398 514170 474970 514226
rect 475026 514170 475094 514226
rect 475150 514170 475218 514226
rect 475274 514170 475342 514226
rect 475398 514170 492970 514226
rect 493026 514170 493094 514226
rect 493150 514170 493218 514226
rect 493274 514170 493342 514226
rect 493398 514170 510970 514226
rect 511026 514170 511094 514226
rect 511150 514170 511218 514226
rect 511274 514170 511342 514226
rect 511398 514170 528970 514226
rect 529026 514170 529094 514226
rect 529150 514170 529218 514226
rect 529274 514170 529342 514226
rect 529398 514170 546970 514226
rect 547026 514170 547094 514226
rect 547150 514170 547218 514226
rect 547274 514170 547342 514226
rect 547398 514170 564970 514226
rect 565026 514170 565094 514226
rect 565150 514170 565218 514226
rect 565274 514170 565342 514226
rect 565398 514170 582970 514226
rect 583026 514170 583094 514226
rect 583150 514170 583218 514226
rect 583274 514170 583342 514226
rect 583398 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 6970 514102
rect 7026 514046 7094 514102
rect 7150 514046 7218 514102
rect 7274 514046 7342 514102
rect 7398 514046 24970 514102
rect 25026 514046 25094 514102
rect 25150 514046 25218 514102
rect 25274 514046 25342 514102
rect 25398 514046 42970 514102
rect 43026 514046 43094 514102
rect 43150 514046 43218 514102
rect 43274 514046 43342 514102
rect 43398 514046 60970 514102
rect 61026 514046 61094 514102
rect 61150 514046 61218 514102
rect 61274 514046 61342 514102
rect 61398 514046 78970 514102
rect 79026 514046 79094 514102
rect 79150 514046 79218 514102
rect 79274 514046 79342 514102
rect 79398 514046 96970 514102
rect 97026 514046 97094 514102
rect 97150 514046 97218 514102
rect 97274 514046 97342 514102
rect 97398 514046 114970 514102
rect 115026 514046 115094 514102
rect 115150 514046 115218 514102
rect 115274 514046 115342 514102
rect 115398 514046 132970 514102
rect 133026 514046 133094 514102
rect 133150 514046 133218 514102
rect 133274 514046 133342 514102
rect 133398 514046 150970 514102
rect 151026 514046 151094 514102
rect 151150 514046 151218 514102
rect 151274 514046 151342 514102
rect 151398 514046 168970 514102
rect 169026 514046 169094 514102
rect 169150 514046 169218 514102
rect 169274 514046 169342 514102
rect 169398 514046 186970 514102
rect 187026 514046 187094 514102
rect 187150 514046 187218 514102
rect 187274 514046 187342 514102
rect 187398 514046 204970 514102
rect 205026 514046 205094 514102
rect 205150 514046 205218 514102
rect 205274 514046 205342 514102
rect 205398 514046 222970 514102
rect 223026 514046 223094 514102
rect 223150 514046 223218 514102
rect 223274 514046 223342 514102
rect 223398 514046 240970 514102
rect 241026 514046 241094 514102
rect 241150 514046 241218 514102
rect 241274 514046 241342 514102
rect 241398 514046 258970 514102
rect 259026 514046 259094 514102
rect 259150 514046 259218 514102
rect 259274 514046 259342 514102
rect 259398 514046 276970 514102
rect 277026 514046 277094 514102
rect 277150 514046 277218 514102
rect 277274 514046 277342 514102
rect 277398 514046 294970 514102
rect 295026 514046 295094 514102
rect 295150 514046 295218 514102
rect 295274 514046 295342 514102
rect 295398 514046 312970 514102
rect 313026 514046 313094 514102
rect 313150 514046 313218 514102
rect 313274 514046 313342 514102
rect 313398 514046 330970 514102
rect 331026 514046 331094 514102
rect 331150 514046 331218 514102
rect 331274 514046 331342 514102
rect 331398 514046 348970 514102
rect 349026 514046 349094 514102
rect 349150 514046 349218 514102
rect 349274 514046 349342 514102
rect 349398 514046 366970 514102
rect 367026 514046 367094 514102
rect 367150 514046 367218 514102
rect 367274 514046 367342 514102
rect 367398 514046 384970 514102
rect 385026 514046 385094 514102
rect 385150 514046 385218 514102
rect 385274 514046 385342 514102
rect 385398 514046 402970 514102
rect 403026 514046 403094 514102
rect 403150 514046 403218 514102
rect 403274 514046 403342 514102
rect 403398 514046 420970 514102
rect 421026 514046 421094 514102
rect 421150 514046 421218 514102
rect 421274 514046 421342 514102
rect 421398 514046 438970 514102
rect 439026 514046 439094 514102
rect 439150 514046 439218 514102
rect 439274 514046 439342 514102
rect 439398 514046 456970 514102
rect 457026 514046 457094 514102
rect 457150 514046 457218 514102
rect 457274 514046 457342 514102
rect 457398 514046 474970 514102
rect 475026 514046 475094 514102
rect 475150 514046 475218 514102
rect 475274 514046 475342 514102
rect 475398 514046 492970 514102
rect 493026 514046 493094 514102
rect 493150 514046 493218 514102
rect 493274 514046 493342 514102
rect 493398 514046 510970 514102
rect 511026 514046 511094 514102
rect 511150 514046 511218 514102
rect 511274 514046 511342 514102
rect 511398 514046 528970 514102
rect 529026 514046 529094 514102
rect 529150 514046 529218 514102
rect 529274 514046 529342 514102
rect 529398 514046 546970 514102
rect 547026 514046 547094 514102
rect 547150 514046 547218 514102
rect 547274 514046 547342 514102
rect 547398 514046 564970 514102
rect 565026 514046 565094 514102
rect 565150 514046 565218 514102
rect 565274 514046 565342 514102
rect 565398 514046 582970 514102
rect 583026 514046 583094 514102
rect 583150 514046 583218 514102
rect 583274 514046 583342 514102
rect 583398 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 6970 513978
rect 7026 513922 7094 513978
rect 7150 513922 7218 513978
rect 7274 513922 7342 513978
rect 7398 513922 24970 513978
rect 25026 513922 25094 513978
rect 25150 513922 25218 513978
rect 25274 513922 25342 513978
rect 25398 513922 42970 513978
rect 43026 513922 43094 513978
rect 43150 513922 43218 513978
rect 43274 513922 43342 513978
rect 43398 513922 60970 513978
rect 61026 513922 61094 513978
rect 61150 513922 61218 513978
rect 61274 513922 61342 513978
rect 61398 513922 78970 513978
rect 79026 513922 79094 513978
rect 79150 513922 79218 513978
rect 79274 513922 79342 513978
rect 79398 513922 96970 513978
rect 97026 513922 97094 513978
rect 97150 513922 97218 513978
rect 97274 513922 97342 513978
rect 97398 513922 114970 513978
rect 115026 513922 115094 513978
rect 115150 513922 115218 513978
rect 115274 513922 115342 513978
rect 115398 513922 132970 513978
rect 133026 513922 133094 513978
rect 133150 513922 133218 513978
rect 133274 513922 133342 513978
rect 133398 513922 150970 513978
rect 151026 513922 151094 513978
rect 151150 513922 151218 513978
rect 151274 513922 151342 513978
rect 151398 513922 168970 513978
rect 169026 513922 169094 513978
rect 169150 513922 169218 513978
rect 169274 513922 169342 513978
rect 169398 513922 186970 513978
rect 187026 513922 187094 513978
rect 187150 513922 187218 513978
rect 187274 513922 187342 513978
rect 187398 513922 204970 513978
rect 205026 513922 205094 513978
rect 205150 513922 205218 513978
rect 205274 513922 205342 513978
rect 205398 513922 222970 513978
rect 223026 513922 223094 513978
rect 223150 513922 223218 513978
rect 223274 513922 223342 513978
rect 223398 513922 240970 513978
rect 241026 513922 241094 513978
rect 241150 513922 241218 513978
rect 241274 513922 241342 513978
rect 241398 513922 258970 513978
rect 259026 513922 259094 513978
rect 259150 513922 259218 513978
rect 259274 513922 259342 513978
rect 259398 513922 276970 513978
rect 277026 513922 277094 513978
rect 277150 513922 277218 513978
rect 277274 513922 277342 513978
rect 277398 513922 294970 513978
rect 295026 513922 295094 513978
rect 295150 513922 295218 513978
rect 295274 513922 295342 513978
rect 295398 513922 312970 513978
rect 313026 513922 313094 513978
rect 313150 513922 313218 513978
rect 313274 513922 313342 513978
rect 313398 513922 330970 513978
rect 331026 513922 331094 513978
rect 331150 513922 331218 513978
rect 331274 513922 331342 513978
rect 331398 513922 348970 513978
rect 349026 513922 349094 513978
rect 349150 513922 349218 513978
rect 349274 513922 349342 513978
rect 349398 513922 366970 513978
rect 367026 513922 367094 513978
rect 367150 513922 367218 513978
rect 367274 513922 367342 513978
rect 367398 513922 384970 513978
rect 385026 513922 385094 513978
rect 385150 513922 385218 513978
rect 385274 513922 385342 513978
rect 385398 513922 402970 513978
rect 403026 513922 403094 513978
rect 403150 513922 403218 513978
rect 403274 513922 403342 513978
rect 403398 513922 420970 513978
rect 421026 513922 421094 513978
rect 421150 513922 421218 513978
rect 421274 513922 421342 513978
rect 421398 513922 438970 513978
rect 439026 513922 439094 513978
rect 439150 513922 439218 513978
rect 439274 513922 439342 513978
rect 439398 513922 456970 513978
rect 457026 513922 457094 513978
rect 457150 513922 457218 513978
rect 457274 513922 457342 513978
rect 457398 513922 474970 513978
rect 475026 513922 475094 513978
rect 475150 513922 475218 513978
rect 475274 513922 475342 513978
rect 475398 513922 492970 513978
rect 493026 513922 493094 513978
rect 493150 513922 493218 513978
rect 493274 513922 493342 513978
rect 493398 513922 510970 513978
rect 511026 513922 511094 513978
rect 511150 513922 511218 513978
rect 511274 513922 511342 513978
rect 511398 513922 528970 513978
rect 529026 513922 529094 513978
rect 529150 513922 529218 513978
rect 529274 513922 529342 513978
rect 529398 513922 546970 513978
rect 547026 513922 547094 513978
rect 547150 513922 547218 513978
rect 547274 513922 547342 513978
rect 547398 513922 564970 513978
rect 565026 513922 565094 513978
rect 565150 513922 565218 513978
rect 565274 513922 565342 513978
rect 565398 513922 582970 513978
rect 583026 513922 583094 513978
rect 583150 513922 583218 513978
rect 583274 513922 583342 513978
rect 583398 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 3250 508350
rect 3306 508294 3374 508350
rect 3430 508294 3498 508350
rect 3554 508294 3622 508350
rect 3678 508294 21250 508350
rect 21306 508294 21374 508350
rect 21430 508294 21498 508350
rect 21554 508294 21622 508350
rect 21678 508294 39250 508350
rect 39306 508294 39374 508350
rect 39430 508294 39498 508350
rect 39554 508294 39622 508350
rect 39678 508294 57250 508350
rect 57306 508294 57374 508350
rect 57430 508294 57498 508350
rect 57554 508294 57622 508350
rect 57678 508294 75250 508350
rect 75306 508294 75374 508350
rect 75430 508294 75498 508350
rect 75554 508294 75622 508350
rect 75678 508294 93250 508350
rect 93306 508294 93374 508350
rect 93430 508294 93498 508350
rect 93554 508294 93622 508350
rect 93678 508294 111250 508350
rect 111306 508294 111374 508350
rect 111430 508294 111498 508350
rect 111554 508294 111622 508350
rect 111678 508294 129250 508350
rect 129306 508294 129374 508350
rect 129430 508294 129498 508350
rect 129554 508294 129622 508350
rect 129678 508294 147250 508350
rect 147306 508294 147374 508350
rect 147430 508294 147498 508350
rect 147554 508294 147622 508350
rect 147678 508294 165250 508350
rect 165306 508294 165374 508350
rect 165430 508294 165498 508350
rect 165554 508294 165622 508350
rect 165678 508294 183250 508350
rect 183306 508294 183374 508350
rect 183430 508294 183498 508350
rect 183554 508294 183622 508350
rect 183678 508294 201250 508350
rect 201306 508294 201374 508350
rect 201430 508294 201498 508350
rect 201554 508294 201622 508350
rect 201678 508294 219250 508350
rect 219306 508294 219374 508350
rect 219430 508294 219498 508350
rect 219554 508294 219622 508350
rect 219678 508294 237250 508350
rect 237306 508294 237374 508350
rect 237430 508294 237498 508350
rect 237554 508294 237622 508350
rect 237678 508294 255250 508350
rect 255306 508294 255374 508350
rect 255430 508294 255498 508350
rect 255554 508294 255622 508350
rect 255678 508294 273250 508350
rect 273306 508294 273374 508350
rect 273430 508294 273498 508350
rect 273554 508294 273622 508350
rect 273678 508294 291250 508350
rect 291306 508294 291374 508350
rect 291430 508294 291498 508350
rect 291554 508294 291622 508350
rect 291678 508294 309250 508350
rect 309306 508294 309374 508350
rect 309430 508294 309498 508350
rect 309554 508294 309622 508350
rect 309678 508294 327250 508350
rect 327306 508294 327374 508350
rect 327430 508294 327498 508350
rect 327554 508294 327622 508350
rect 327678 508294 345250 508350
rect 345306 508294 345374 508350
rect 345430 508294 345498 508350
rect 345554 508294 345622 508350
rect 345678 508294 363250 508350
rect 363306 508294 363374 508350
rect 363430 508294 363498 508350
rect 363554 508294 363622 508350
rect 363678 508294 381250 508350
rect 381306 508294 381374 508350
rect 381430 508294 381498 508350
rect 381554 508294 381622 508350
rect 381678 508294 399250 508350
rect 399306 508294 399374 508350
rect 399430 508294 399498 508350
rect 399554 508294 399622 508350
rect 399678 508294 417250 508350
rect 417306 508294 417374 508350
rect 417430 508294 417498 508350
rect 417554 508294 417622 508350
rect 417678 508294 435250 508350
rect 435306 508294 435374 508350
rect 435430 508294 435498 508350
rect 435554 508294 435622 508350
rect 435678 508294 453250 508350
rect 453306 508294 453374 508350
rect 453430 508294 453498 508350
rect 453554 508294 453622 508350
rect 453678 508294 471250 508350
rect 471306 508294 471374 508350
rect 471430 508294 471498 508350
rect 471554 508294 471622 508350
rect 471678 508294 489250 508350
rect 489306 508294 489374 508350
rect 489430 508294 489498 508350
rect 489554 508294 489622 508350
rect 489678 508294 507250 508350
rect 507306 508294 507374 508350
rect 507430 508294 507498 508350
rect 507554 508294 507622 508350
rect 507678 508294 525250 508350
rect 525306 508294 525374 508350
rect 525430 508294 525498 508350
rect 525554 508294 525622 508350
rect 525678 508294 543250 508350
rect 543306 508294 543374 508350
rect 543430 508294 543498 508350
rect 543554 508294 543622 508350
rect 543678 508294 561250 508350
rect 561306 508294 561374 508350
rect 561430 508294 561498 508350
rect 561554 508294 561622 508350
rect 561678 508294 579250 508350
rect 579306 508294 579374 508350
rect 579430 508294 579498 508350
rect 579554 508294 579622 508350
rect 579678 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 3250 508226
rect 3306 508170 3374 508226
rect 3430 508170 3498 508226
rect 3554 508170 3622 508226
rect 3678 508170 21250 508226
rect 21306 508170 21374 508226
rect 21430 508170 21498 508226
rect 21554 508170 21622 508226
rect 21678 508170 39250 508226
rect 39306 508170 39374 508226
rect 39430 508170 39498 508226
rect 39554 508170 39622 508226
rect 39678 508170 57250 508226
rect 57306 508170 57374 508226
rect 57430 508170 57498 508226
rect 57554 508170 57622 508226
rect 57678 508170 75250 508226
rect 75306 508170 75374 508226
rect 75430 508170 75498 508226
rect 75554 508170 75622 508226
rect 75678 508170 93250 508226
rect 93306 508170 93374 508226
rect 93430 508170 93498 508226
rect 93554 508170 93622 508226
rect 93678 508170 111250 508226
rect 111306 508170 111374 508226
rect 111430 508170 111498 508226
rect 111554 508170 111622 508226
rect 111678 508170 129250 508226
rect 129306 508170 129374 508226
rect 129430 508170 129498 508226
rect 129554 508170 129622 508226
rect 129678 508170 147250 508226
rect 147306 508170 147374 508226
rect 147430 508170 147498 508226
rect 147554 508170 147622 508226
rect 147678 508170 165250 508226
rect 165306 508170 165374 508226
rect 165430 508170 165498 508226
rect 165554 508170 165622 508226
rect 165678 508170 183250 508226
rect 183306 508170 183374 508226
rect 183430 508170 183498 508226
rect 183554 508170 183622 508226
rect 183678 508170 201250 508226
rect 201306 508170 201374 508226
rect 201430 508170 201498 508226
rect 201554 508170 201622 508226
rect 201678 508170 219250 508226
rect 219306 508170 219374 508226
rect 219430 508170 219498 508226
rect 219554 508170 219622 508226
rect 219678 508170 237250 508226
rect 237306 508170 237374 508226
rect 237430 508170 237498 508226
rect 237554 508170 237622 508226
rect 237678 508170 255250 508226
rect 255306 508170 255374 508226
rect 255430 508170 255498 508226
rect 255554 508170 255622 508226
rect 255678 508170 273250 508226
rect 273306 508170 273374 508226
rect 273430 508170 273498 508226
rect 273554 508170 273622 508226
rect 273678 508170 291250 508226
rect 291306 508170 291374 508226
rect 291430 508170 291498 508226
rect 291554 508170 291622 508226
rect 291678 508170 309250 508226
rect 309306 508170 309374 508226
rect 309430 508170 309498 508226
rect 309554 508170 309622 508226
rect 309678 508170 327250 508226
rect 327306 508170 327374 508226
rect 327430 508170 327498 508226
rect 327554 508170 327622 508226
rect 327678 508170 345250 508226
rect 345306 508170 345374 508226
rect 345430 508170 345498 508226
rect 345554 508170 345622 508226
rect 345678 508170 363250 508226
rect 363306 508170 363374 508226
rect 363430 508170 363498 508226
rect 363554 508170 363622 508226
rect 363678 508170 381250 508226
rect 381306 508170 381374 508226
rect 381430 508170 381498 508226
rect 381554 508170 381622 508226
rect 381678 508170 399250 508226
rect 399306 508170 399374 508226
rect 399430 508170 399498 508226
rect 399554 508170 399622 508226
rect 399678 508170 417250 508226
rect 417306 508170 417374 508226
rect 417430 508170 417498 508226
rect 417554 508170 417622 508226
rect 417678 508170 435250 508226
rect 435306 508170 435374 508226
rect 435430 508170 435498 508226
rect 435554 508170 435622 508226
rect 435678 508170 453250 508226
rect 453306 508170 453374 508226
rect 453430 508170 453498 508226
rect 453554 508170 453622 508226
rect 453678 508170 471250 508226
rect 471306 508170 471374 508226
rect 471430 508170 471498 508226
rect 471554 508170 471622 508226
rect 471678 508170 489250 508226
rect 489306 508170 489374 508226
rect 489430 508170 489498 508226
rect 489554 508170 489622 508226
rect 489678 508170 507250 508226
rect 507306 508170 507374 508226
rect 507430 508170 507498 508226
rect 507554 508170 507622 508226
rect 507678 508170 525250 508226
rect 525306 508170 525374 508226
rect 525430 508170 525498 508226
rect 525554 508170 525622 508226
rect 525678 508170 543250 508226
rect 543306 508170 543374 508226
rect 543430 508170 543498 508226
rect 543554 508170 543622 508226
rect 543678 508170 561250 508226
rect 561306 508170 561374 508226
rect 561430 508170 561498 508226
rect 561554 508170 561622 508226
rect 561678 508170 579250 508226
rect 579306 508170 579374 508226
rect 579430 508170 579498 508226
rect 579554 508170 579622 508226
rect 579678 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 3250 508102
rect 3306 508046 3374 508102
rect 3430 508046 3498 508102
rect 3554 508046 3622 508102
rect 3678 508046 21250 508102
rect 21306 508046 21374 508102
rect 21430 508046 21498 508102
rect 21554 508046 21622 508102
rect 21678 508046 39250 508102
rect 39306 508046 39374 508102
rect 39430 508046 39498 508102
rect 39554 508046 39622 508102
rect 39678 508046 57250 508102
rect 57306 508046 57374 508102
rect 57430 508046 57498 508102
rect 57554 508046 57622 508102
rect 57678 508046 75250 508102
rect 75306 508046 75374 508102
rect 75430 508046 75498 508102
rect 75554 508046 75622 508102
rect 75678 508046 93250 508102
rect 93306 508046 93374 508102
rect 93430 508046 93498 508102
rect 93554 508046 93622 508102
rect 93678 508046 111250 508102
rect 111306 508046 111374 508102
rect 111430 508046 111498 508102
rect 111554 508046 111622 508102
rect 111678 508046 129250 508102
rect 129306 508046 129374 508102
rect 129430 508046 129498 508102
rect 129554 508046 129622 508102
rect 129678 508046 147250 508102
rect 147306 508046 147374 508102
rect 147430 508046 147498 508102
rect 147554 508046 147622 508102
rect 147678 508046 165250 508102
rect 165306 508046 165374 508102
rect 165430 508046 165498 508102
rect 165554 508046 165622 508102
rect 165678 508046 183250 508102
rect 183306 508046 183374 508102
rect 183430 508046 183498 508102
rect 183554 508046 183622 508102
rect 183678 508046 201250 508102
rect 201306 508046 201374 508102
rect 201430 508046 201498 508102
rect 201554 508046 201622 508102
rect 201678 508046 219250 508102
rect 219306 508046 219374 508102
rect 219430 508046 219498 508102
rect 219554 508046 219622 508102
rect 219678 508046 237250 508102
rect 237306 508046 237374 508102
rect 237430 508046 237498 508102
rect 237554 508046 237622 508102
rect 237678 508046 255250 508102
rect 255306 508046 255374 508102
rect 255430 508046 255498 508102
rect 255554 508046 255622 508102
rect 255678 508046 273250 508102
rect 273306 508046 273374 508102
rect 273430 508046 273498 508102
rect 273554 508046 273622 508102
rect 273678 508046 291250 508102
rect 291306 508046 291374 508102
rect 291430 508046 291498 508102
rect 291554 508046 291622 508102
rect 291678 508046 309250 508102
rect 309306 508046 309374 508102
rect 309430 508046 309498 508102
rect 309554 508046 309622 508102
rect 309678 508046 327250 508102
rect 327306 508046 327374 508102
rect 327430 508046 327498 508102
rect 327554 508046 327622 508102
rect 327678 508046 345250 508102
rect 345306 508046 345374 508102
rect 345430 508046 345498 508102
rect 345554 508046 345622 508102
rect 345678 508046 363250 508102
rect 363306 508046 363374 508102
rect 363430 508046 363498 508102
rect 363554 508046 363622 508102
rect 363678 508046 381250 508102
rect 381306 508046 381374 508102
rect 381430 508046 381498 508102
rect 381554 508046 381622 508102
rect 381678 508046 399250 508102
rect 399306 508046 399374 508102
rect 399430 508046 399498 508102
rect 399554 508046 399622 508102
rect 399678 508046 417250 508102
rect 417306 508046 417374 508102
rect 417430 508046 417498 508102
rect 417554 508046 417622 508102
rect 417678 508046 435250 508102
rect 435306 508046 435374 508102
rect 435430 508046 435498 508102
rect 435554 508046 435622 508102
rect 435678 508046 453250 508102
rect 453306 508046 453374 508102
rect 453430 508046 453498 508102
rect 453554 508046 453622 508102
rect 453678 508046 471250 508102
rect 471306 508046 471374 508102
rect 471430 508046 471498 508102
rect 471554 508046 471622 508102
rect 471678 508046 489250 508102
rect 489306 508046 489374 508102
rect 489430 508046 489498 508102
rect 489554 508046 489622 508102
rect 489678 508046 507250 508102
rect 507306 508046 507374 508102
rect 507430 508046 507498 508102
rect 507554 508046 507622 508102
rect 507678 508046 525250 508102
rect 525306 508046 525374 508102
rect 525430 508046 525498 508102
rect 525554 508046 525622 508102
rect 525678 508046 543250 508102
rect 543306 508046 543374 508102
rect 543430 508046 543498 508102
rect 543554 508046 543622 508102
rect 543678 508046 561250 508102
rect 561306 508046 561374 508102
rect 561430 508046 561498 508102
rect 561554 508046 561622 508102
rect 561678 508046 579250 508102
rect 579306 508046 579374 508102
rect 579430 508046 579498 508102
rect 579554 508046 579622 508102
rect 579678 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 3250 507978
rect 3306 507922 3374 507978
rect 3430 507922 3498 507978
rect 3554 507922 3622 507978
rect 3678 507922 21250 507978
rect 21306 507922 21374 507978
rect 21430 507922 21498 507978
rect 21554 507922 21622 507978
rect 21678 507922 39250 507978
rect 39306 507922 39374 507978
rect 39430 507922 39498 507978
rect 39554 507922 39622 507978
rect 39678 507922 57250 507978
rect 57306 507922 57374 507978
rect 57430 507922 57498 507978
rect 57554 507922 57622 507978
rect 57678 507922 75250 507978
rect 75306 507922 75374 507978
rect 75430 507922 75498 507978
rect 75554 507922 75622 507978
rect 75678 507922 93250 507978
rect 93306 507922 93374 507978
rect 93430 507922 93498 507978
rect 93554 507922 93622 507978
rect 93678 507922 111250 507978
rect 111306 507922 111374 507978
rect 111430 507922 111498 507978
rect 111554 507922 111622 507978
rect 111678 507922 129250 507978
rect 129306 507922 129374 507978
rect 129430 507922 129498 507978
rect 129554 507922 129622 507978
rect 129678 507922 147250 507978
rect 147306 507922 147374 507978
rect 147430 507922 147498 507978
rect 147554 507922 147622 507978
rect 147678 507922 165250 507978
rect 165306 507922 165374 507978
rect 165430 507922 165498 507978
rect 165554 507922 165622 507978
rect 165678 507922 183250 507978
rect 183306 507922 183374 507978
rect 183430 507922 183498 507978
rect 183554 507922 183622 507978
rect 183678 507922 201250 507978
rect 201306 507922 201374 507978
rect 201430 507922 201498 507978
rect 201554 507922 201622 507978
rect 201678 507922 219250 507978
rect 219306 507922 219374 507978
rect 219430 507922 219498 507978
rect 219554 507922 219622 507978
rect 219678 507922 237250 507978
rect 237306 507922 237374 507978
rect 237430 507922 237498 507978
rect 237554 507922 237622 507978
rect 237678 507922 255250 507978
rect 255306 507922 255374 507978
rect 255430 507922 255498 507978
rect 255554 507922 255622 507978
rect 255678 507922 273250 507978
rect 273306 507922 273374 507978
rect 273430 507922 273498 507978
rect 273554 507922 273622 507978
rect 273678 507922 291250 507978
rect 291306 507922 291374 507978
rect 291430 507922 291498 507978
rect 291554 507922 291622 507978
rect 291678 507922 309250 507978
rect 309306 507922 309374 507978
rect 309430 507922 309498 507978
rect 309554 507922 309622 507978
rect 309678 507922 327250 507978
rect 327306 507922 327374 507978
rect 327430 507922 327498 507978
rect 327554 507922 327622 507978
rect 327678 507922 345250 507978
rect 345306 507922 345374 507978
rect 345430 507922 345498 507978
rect 345554 507922 345622 507978
rect 345678 507922 363250 507978
rect 363306 507922 363374 507978
rect 363430 507922 363498 507978
rect 363554 507922 363622 507978
rect 363678 507922 381250 507978
rect 381306 507922 381374 507978
rect 381430 507922 381498 507978
rect 381554 507922 381622 507978
rect 381678 507922 399250 507978
rect 399306 507922 399374 507978
rect 399430 507922 399498 507978
rect 399554 507922 399622 507978
rect 399678 507922 417250 507978
rect 417306 507922 417374 507978
rect 417430 507922 417498 507978
rect 417554 507922 417622 507978
rect 417678 507922 435250 507978
rect 435306 507922 435374 507978
rect 435430 507922 435498 507978
rect 435554 507922 435622 507978
rect 435678 507922 453250 507978
rect 453306 507922 453374 507978
rect 453430 507922 453498 507978
rect 453554 507922 453622 507978
rect 453678 507922 471250 507978
rect 471306 507922 471374 507978
rect 471430 507922 471498 507978
rect 471554 507922 471622 507978
rect 471678 507922 489250 507978
rect 489306 507922 489374 507978
rect 489430 507922 489498 507978
rect 489554 507922 489622 507978
rect 489678 507922 507250 507978
rect 507306 507922 507374 507978
rect 507430 507922 507498 507978
rect 507554 507922 507622 507978
rect 507678 507922 525250 507978
rect 525306 507922 525374 507978
rect 525430 507922 525498 507978
rect 525554 507922 525622 507978
rect 525678 507922 543250 507978
rect 543306 507922 543374 507978
rect 543430 507922 543498 507978
rect 543554 507922 543622 507978
rect 543678 507922 561250 507978
rect 561306 507922 561374 507978
rect 561430 507922 561498 507978
rect 561554 507922 561622 507978
rect 561678 507922 579250 507978
rect 579306 507922 579374 507978
rect 579430 507922 579498 507978
rect 579554 507922 579622 507978
rect 579678 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 6970 496350
rect 7026 496294 7094 496350
rect 7150 496294 7218 496350
rect 7274 496294 7342 496350
rect 7398 496294 24970 496350
rect 25026 496294 25094 496350
rect 25150 496294 25218 496350
rect 25274 496294 25342 496350
rect 25398 496294 42970 496350
rect 43026 496294 43094 496350
rect 43150 496294 43218 496350
rect 43274 496294 43342 496350
rect 43398 496294 60970 496350
rect 61026 496294 61094 496350
rect 61150 496294 61218 496350
rect 61274 496294 61342 496350
rect 61398 496294 78970 496350
rect 79026 496294 79094 496350
rect 79150 496294 79218 496350
rect 79274 496294 79342 496350
rect 79398 496294 96970 496350
rect 97026 496294 97094 496350
rect 97150 496294 97218 496350
rect 97274 496294 97342 496350
rect 97398 496294 114970 496350
rect 115026 496294 115094 496350
rect 115150 496294 115218 496350
rect 115274 496294 115342 496350
rect 115398 496294 132970 496350
rect 133026 496294 133094 496350
rect 133150 496294 133218 496350
rect 133274 496294 133342 496350
rect 133398 496294 150970 496350
rect 151026 496294 151094 496350
rect 151150 496294 151218 496350
rect 151274 496294 151342 496350
rect 151398 496294 168970 496350
rect 169026 496294 169094 496350
rect 169150 496294 169218 496350
rect 169274 496294 169342 496350
rect 169398 496294 186970 496350
rect 187026 496294 187094 496350
rect 187150 496294 187218 496350
rect 187274 496294 187342 496350
rect 187398 496333 510970 496350
rect 187398 496294 219878 496333
rect -1916 496277 219878 496294
rect 219934 496277 220002 496333
rect 220058 496277 250598 496333
rect 250654 496277 250722 496333
rect 250778 496277 281318 496333
rect 281374 496277 281442 496333
rect 281498 496277 312038 496333
rect 312094 496277 312162 496333
rect 312218 496277 342758 496333
rect 342814 496277 342882 496333
rect 342938 496277 373478 496333
rect 373534 496277 373602 496333
rect 373658 496277 404198 496333
rect 404254 496277 404322 496333
rect 404378 496277 434918 496333
rect 434974 496277 435042 496333
rect 435098 496277 465638 496333
rect 465694 496277 465762 496333
rect 465818 496277 496358 496333
rect 496414 496277 496482 496333
rect 496538 496294 510970 496333
rect 511026 496294 511094 496350
rect 511150 496294 511218 496350
rect 511274 496294 511342 496350
rect 511398 496294 528970 496350
rect 529026 496294 529094 496350
rect 529150 496294 529218 496350
rect 529274 496294 529342 496350
rect 529398 496294 546970 496350
rect 547026 496294 547094 496350
rect 547150 496294 547218 496350
rect 547274 496294 547342 496350
rect 547398 496294 564970 496350
rect 565026 496294 565094 496350
rect 565150 496294 565218 496350
rect 565274 496294 565342 496350
rect 565398 496294 582970 496350
rect 583026 496294 583094 496350
rect 583150 496294 583218 496350
rect 583274 496294 583342 496350
rect 583398 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 496538 496277 597980 496294
rect -1916 496226 597980 496277
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 6970 496226
rect 7026 496170 7094 496226
rect 7150 496170 7218 496226
rect 7274 496170 7342 496226
rect 7398 496170 24970 496226
rect 25026 496170 25094 496226
rect 25150 496170 25218 496226
rect 25274 496170 25342 496226
rect 25398 496170 42970 496226
rect 43026 496170 43094 496226
rect 43150 496170 43218 496226
rect 43274 496170 43342 496226
rect 43398 496170 60970 496226
rect 61026 496170 61094 496226
rect 61150 496170 61218 496226
rect 61274 496170 61342 496226
rect 61398 496170 78970 496226
rect 79026 496170 79094 496226
rect 79150 496170 79218 496226
rect 79274 496170 79342 496226
rect 79398 496170 96970 496226
rect 97026 496170 97094 496226
rect 97150 496170 97218 496226
rect 97274 496170 97342 496226
rect 97398 496170 114970 496226
rect 115026 496170 115094 496226
rect 115150 496170 115218 496226
rect 115274 496170 115342 496226
rect 115398 496170 132970 496226
rect 133026 496170 133094 496226
rect 133150 496170 133218 496226
rect 133274 496170 133342 496226
rect 133398 496170 150970 496226
rect 151026 496170 151094 496226
rect 151150 496170 151218 496226
rect 151274 496170 151342 496226
rect 151398 496170 168970 496226
rect 169026 496170 169094 496226
rect 169150 496170 169218 496226
rect 169274 496170 169342 496226
rect 169398 496170 186970 496226
rect 187026 496170 187094 496226
rect 187150 496170 187218 496226
rect 187274 496170 187342 496226
rect 187398 496209 510970 496226
rect 187398 496170 219878 496209
rect -1916 496153 219878 496170
rect 219934 496153 220002 496209
rect 220058 496153 250598 496209
rect 250654 496153 250722 496209
rect 250778 496153 281318 496209
rect 281374 496153 281442 496209
rect 281498 496153 312038 496209
rect 312094 496153 312162 496209
rect 312218 496153 342758 496209
rect 342814 496153 342882 496209
rect 342938 496153 373478 496209
rect 373534 496153 373602 496209
rect 373658 496153 404198 496209
rect 404254 496153 404322 496209
rect 404378 496153 434918 496209
rect 434974 496153 435042 496209
rect 435098 496153 465638 496209
rect 465694 496153 465762 496209
rect 465818 496153 496358 496209
rect 496414 496153 496482 496209
rect 496538 496170 510970 496209
rect 511026 496170 511094 496226
rect 511150 496170 511218 496226
rect 511274 496170 511342 496226
rect 511398 496170 528970 496226
rect 529026 496170 529094 496226
rect 529150 496170 529218 496226
rect 529274 496170 529342 496226
rect 529398 496170 546970 496226
rect 547026 496170 547094 496226
rect 547150 496170 547218 496226
rect 547274 496170 547342 496226
rect 547398 496170 564970 496226
rect 565026 496170 565094 496226
rect 565150 496170 565218 496226
rect 565274 496170 565342 496226
rect 565398 496170 582970 496226
rect 583026 496170 583094 496226
rect 583150 496170 583218 496226
rect 583274 496170 583342 496226
rect 583398 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 496538 496153 597980 496170
rect -1916 496102 597980 496153
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 6970 496102
rect 7026 496046 7094 496102
rect 7150 496046 7218 496102
rect 7274 496046 7342 496102
rect 7398 496046 24970 496102
rect 25026 496046 25094 496102
rect 25150 496046 25218 496102
rect 25274 496046 25342 496102
rect 25398 496046 42970 496102
rect 43026 496046 43094 496102
rect 43150 496046 43218 496102
rect 43274 496046 43342 496102
rect 43398 496046 60970 496102
rect 61026 496046 61094 496102
rect 61150 496046 61218 496102
rect 61274 496046 61342 496102
rect 61398 496046 78970 496102
rect 79026 496046 79094 496102
rect 79150 496046 79218 496102
rect 79274 496046 79342 496102
rect 79398 496046 96970 496102
rect 97026 496046 97094 496102
rect 97150 496046 97218 496102
rect 97274 496046 97342 496102
rect 97398 496046 114970 496102
rect 115026 496046 115094 496102
rect 115150 496046 115218 496102
rect 115274 496046 115342 496102
rect 115398 496046 132970 496102
rect 133026 496046 133094 496102
rect 133150 496046 133218 496102
rect 133274 496046 133342 496102
rect 133398 496046 150970 496102
rect 151026 496046 151094 496102
rect 151150 496046 151218 496102
rect 151274 496046 151342 496102
rect 151398 496046 168970 496102
rect 169026 496046 169094 496102
rect 169150 496046 169218 496102
rect 169274 496046 169342 496102
rect 169398 496046 186970 496102
rect 187026 496046 187094 496102
rect 187150 496046 187218 496102
rect 187274 496046 187342 496102
rect 187398 496085 510970 496102
rect 187398 496046 219878 496085
rect -1916 496029 219878 496046
rect 219934 496029 220002 496085
rect 220058 496029 250598 496085
rect 250654 496029 250722 496085
rect 250778 496029 281318 496085
rect 281374 496029 281442 496085
rect 281498 496029 312038 496085
rect 312094 496029 312162 496085
rect 312218 496029 342758 496085
rect 342814 496029 342882 496085
rect 342938 496029 373478 496085
rect 373534 496029 373602 496085
rect 373658 496029 404198 496085
rect 404254 496029 404322 496085
rect 404378 496029 434918 496085
rect 434974 496029 435042 496085
rect 435098 496029 465638 496085
rect 465694 496029 465762 496085
rect 465818 496029 496358 496085
rect 496414 496029 496482 496085
rect 496538 496046 510970 496085
rect 511026 496046 511094 496102
rect 511150 496046 511218 496102
rect 511274 496046 511342 496102
rect 511398 496046 528970 496102
rect 529026 496046 529094 496102
rect 529150 496046 529218 496102
rect 529274 496046 529342 496102
rect 529398 496046 546970 496102
rect 547026 496046 547094 496102
rect 547150 496046 547218 496102
rect 547274 496046 547342 496102
rect 547398 496046 564970 496102
rect 565026 496046 565094 496102
rect 565150 496046 565218 496102
rect 565274 496046 565342 496102
rect 565398 496046 582970 496102
rect 583026 496046 583094 496102
rect 583150 496046 583218 496102
rect 583274 496046 583342 496102
rect 583398 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 496538 496029 597980 496046
rect -1916 495978 597980 496029
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 6970 495978
rect 7026 495922 7094 495978
rect 7150 495922 7218 495978
rect 7274 495922 7342 495978
rect 7398 495922 24970 495978
rect 25026 495922 25094 495978
rect 25150 495922 25218 495978
rect 25274 495922 25342 495978
rect 25398 495922 42970 495978
rect 43026 495922 43094 495978
rect 43150 495922 43218 495978
rect 43274 495922 43342 495978
rect 43398 495922 60970 495978
rect 61026 495922 61094 495978
rect 61150 495922 61218 495978
rect 61274 495922 61342 495978
rect 61398 495922 78970 495978
rect 79026 495922 79094 495978
rect 79150 495922 79218 495978
rect 79274 495922 79342 495978
rect 79398 495922 96970 495978
rect 97026 495922 97094 495978
rect 97150 495922 97218 495978
rect 97274 495922 97342 495978
rect 97398 495922 114970 495978
rect 115026 495922 115094 495978
rect 115150 495922 115218 495978
rect 115274 495922 115342 495978
rect 115398 495922 132970 495978
rect 133026 495922 133094 495978
rect 133150 495922 133218 495978
rect 133274 495922 133342 495978
rect 133398 495922 150970 495978
rect 151026 495922 151094 495978
rect 151150 495922 151218 495978
rect 151274 495922 151342 495978
rect 151398 495922 168970 495978
rect 169026 495922 169094 495978
rect 169150 495922 169218 495978
rect 169274 495922 169342 495978
rect 169398 495922 186970 495978
rect 187026 495922 187094 495978
rect 187150 495922 187218 495978
rect 187274 495922 187342 495978
rect 187398 495961 510970 495978
rect 187398 495922 219878 495961
rect -1916 495905 219878 495922
rect 219934 495905 220002 495961
rect 220058 495905 250598 495961
rect 250654 495905 250722 495961
rect 250778 495905 281318 495961
rect 281374 495905 281442 495961
rect 281498 495905 312038 495961
rect 312094 495905 312162 495961
rect 312218 495905 342758 495961
rect 342814 495905 342882 495961
rect 342938 495905 373478 495961
rect 373534 495905 373602 495961
rect 373658 495905 404198 495961
rect 404254 495905 404322 495961
rect 404378 495905 434918 495961
rect 434974 495905 435042 495961
rect 435098 495905 465638 495961
rect 465694 495905 465762 495961
rect 465818 495905 496358 495961
rect 496414 495905 496482 495961
rect 496538 495922 510970 495961
rect 511026 495922 511094 495978
rect 511150 495922 511218 495978
rect 511274 495922 511342 495978
rect 511398 495922 528970 495978
rect 529026 495922 529094 495978
rect 529150 495922 529218 495978
rect 529274 495922 529342 495978
rect 529398 495922 546970 495978
rect 547026 495922 547094 495978
rect 547150 495922 547218 495978
rect 547274 495922 547342 495978
rect 547398 495922 564970 495978
rect 565026 495922 565094 495978
rect 565150 495922 565218 495978
rect 565274 495922 565342 495978
rect 565398 495922 582970 495978
rect 583026 495922 583094 495978
rect 583150 495922 583218 495978
rect 583274 495922 583342 495978
rect 583398 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 496538 495905 597980 495922
rect -1916 495826 597980 495905
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 3250 490350
rect 3306 490294 3374 490350
rect 3430 490294 3498 490350
rect 3554 490294 3622 490350
rect 3678 490294 21250 490350
rect 21306 490294 21374 490350
rect 21430 490294 21498 490350
rect 21554 490294 21622 490350
rect 21678 490294 39250 490350
rect 39306 490294 39374 490350
rect 39430 490294 39498 490350
rect 39554 490294 39622 490350
rect 39678 490294 57250 490350
rect 57306 490294 57374 490350
rect 57430 490294 57498 490350
rect 57554 490294 57622 490350
rect 57678 490294 75250 490350
rect 75306 490294 75374 490350
rect 75430 490294 75498 490350
rect 75554 490294 75622 490350
rect 75678 490294 93250 490350
rect 93306 490294 93374 490350
rect 93430 490294 93498 490350
rect 93554 490294 93622 490350
rect 93678 490294 111250 490350
rect 111306 490294 111374 490350
rect 111430 490294 111498 490350
rect 111554 490294 111622 490350
rect 111678 490294 129250 490350
rect 129306 490294 129374 490350
rect 129430 490294 129498 490350
rect 129554 490294 129622 490350
rect 129678 490294 147250 490350
rect 147306 490294 147374 490350
rect 147430 490294 147498 490350
rect 147554 490294 147622 490350
rect 147678 490294 165250 490350
rect 165306 490294 165374 490350
rect 165430 490294 165498 490350
rect 165554 490294 165622 490350
rect 165678 490294 183250 490350
rect 183306 490294 183374 490350
rect 183430 490294 183498 490350
rect 183554 490294 183622 490350
rect 183678 490294 201250 490350
rect 201306 490294 201374 490350
rect 201430 490294 201498 490350
rect 201554 490294 201622 490350
rect 201678 490294 204518 490350
rect 204574 490294 204642 490350
rect 204698 490294 235238 490350
rect 235294 490294 235362 490350
rect 235418 490294 265958 490350
rect 266014 490294 266082 490350
rect 266138 490294 296678 490350
rect 296734 490294 296802 490350
rect 296858 490294 327398 490350
rect 327454 490294 327522 490350
rect 327578 490294 358118 490350
rect 358174 490294 358242 490350
rect 358298 490294 388838 490350
rect 388894 490294 388962 490350
rect 389018 490294 419558 490350
rect 419614 490294 419682 490350
rect 419738 490294 450278 490350
rect 450334 490294 450402 490350
rect 450458 490294 480998 490350
rect 481054 490294 481122 490350
rect 481178 490294 507250 490350
rect 507306 490294 507374 490350
rect 507430 490294 507498 490350
rect 507554 490294 507622 490350
rect 507678 490294 525250 490350
rect 525306 490294 525374 490350
rect 525430 490294 525498 490350
rect 525554 490294 525622 490350
rect 525678 490294 543250 490350
rect 543306 490294 543374 490350
rect 543430 490294 543498 490350
rect 543554 490294 543622 490350
rect 543678 490294 561250 490350
rect 561306 490294 561374 490350
rect 561430 490294 561498 490350
rect 561554 490294 561622 490350
rect 561678 490294 579250 490350
rect 579306 490294 579374 490350
rect 579430 490294 579498 490350
rect 579554 490294 579622 490350
rect 579678 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 3250 490226
rect 3306 490170 3374 490226
rect 3430 490170 3498 490226
rect 3554 490170 3622 490226
rect 3678 490170 21250 490226
rect 21306 490170 21374 490226
rect 21430 490170 21498 490226
rect 21554 490170 21622 490226
rect 21678 490170 39250 490226
rect 39306 490170 39374 490226
rect 39430 490170 39498 490226
rect 39554 490170 39622 490226
rect 39678 490170 57250 490226
rect 57306 490170 57374 490226
rect 57430 490170 57498 490226
rect 57554 490170 57622 490226
rect 57678 490170 75250 490226
rect 75306 490170 75374 490226
rect 75430 490170 75498 490226
rect 75554 490170 75622 490226
rect 75678 490170 93250 490226
rect 93306 490170 93374 490226
rect 93430 490170 93498 490226
rect 93554 490170 93622 490226
rect 93678 490170 111250 490226
rect 111306 490170 111374 490226
rect 111430 490170 111498 490226
rect 111554 490170 111622 490226
rect 111678 490170 129250 490226
rect 129306 490170 129374 490226
rect 129430 490170 129498 490226
rect 129554 490170 129622 490226
rect 129678 490170 147250 490226
rect 147306 490170 147374 490226
rect 147430 490170 147498 490226
rect 147554 490170 147622 490226
rect 147678 490170 165250 490226
rect 165306 490170 165374 490226
rect 165430 490170 165498 490226
rect 165554 490170 165622 490226
rect 165678 490170 183250 490226
rect 183306 490170 183374 490226
rect 183430 490170 183498 490226
rect 183554 490170 183622 490226
rect 183678 490170 201250 490226
rect 201306 490170 201374 490226
rect 201430 490170 201498 490226
rect 201554 490170 201622 490226
rect 201678 490170 204518 490226
rect 204574 490170 204642 490226
rect 204698 490170 235238 490226
rect 235294 490170 235362 490226
rect 235418 490170 265958 490226
rect 266014 490170 266082 490226
rect 266138 490170 296678 490226
rect 296734 490170 296802 490226
rect 296858 490170 327398 490226
rect 327454 490170 327522 490226
rect 327578 490170 358118 490226
rect 358174 490170 358242 490226
rect 358298 490170 388838 490226
rect 388894 490170 388962 490226
rect 389018 490170 419558 490226
rect 419614 490170 419682 490226
rect 419738 490170 450278 490226
rect 450334 490170 450402 490226
rect 450458 490170 480998 490226
rect 481054 490170 481122 490226
rect 481178 490170 507250 490226
rect 507306 490170 507374 490226
rect 507430 490170 507498 490226
rect 507554 490170 507622 490226
rect 507678 490170 525250 490226
rect 525306 490170 525374 490226
rect 525430 490170 525498 490226
rect 525554 490170 525622 490226
rect 525678 490170 543250 490226
rect 543306 490170 543374 490226
rect 543430 490170 543498 490226
rect 543554 490170 543622 490226
rect 543678 490170 561250 490226
rect 561306 490170 561374 490226
rect 561430 490170 561498 490226
rect 561554 490170 561622 490226
rect 561678 490170 579250 490226
rect 579306 490170 579374 490226
rect 579430 490170 579498 490226
rect 579554 490170 579622 490226
rect 579678 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 3250 490102
rect 3306 490046 3374 490102
rect 3430 490046 3498 490102
rect 3554 490046 3622 490102
rect 3678 490046 21250 490102
rect 21306 490046 21374 490102
rect 21430 490046 21498 490102
rect 21554 490046 21622 490102
rect 21678 490046 39250 490102
rect 39306 490046 39374 490102
rect 39430 490046 39498 490102
rect 39554 490046 39622 490102
rect 39678 490046 57250 490102
rect 57306 490046 57374 490102
rect 57430 490046 57498 490102
rect 57554 490046 57622 490102
rect 57678 490046 75250 490102
rect 75306 490046 75374 490102
rect 75430 490046 75498 490102
rect 75554 490046 75622 490102
rect 75678 490046 93250 490102
rect 93306 490046 93374 490102
rect 93430 490046 93498 490102
rect 93554 490046 93622 490102
rect 93678 490046 111250 490102
rect 111306 490046 111374 490102
rect 111430 490046 111498 490102
rect 111554 490046 111622 490102
rect 111678 490046 129250 490102
rect 129306 490046 129374 490102
rect 129430 490046 129498 490102
rect 129554 490046 129622 490102
rect 129678 490046 147250 490102
rect 147306 490046 147374 490102
rect 147430 490046 147498 490102
rect 147554 490046 147622 490102
rect 147678 490046 165250 490102
rect 165306 490046 165374 490102
rect 165430 490046 165498 490102
rect 165554 490046 165622 490102
rect 165678 490046 183250 490102
rect 183306 490046 183374 490102
rect 183430 490046 183498 490102
rect 183554 490046 183622 490102
rect 183678 490046 201250 490102
rect 201306 490046 201374 490102
rect 201430 490046 201498 490102
rect 201554 490046 201622 490102
rect 201678 490046 204518 490102
rect 204574 490046 204642 490102
rect 204698 490046 235238 490102
rect 235294 490046 235362 490102
rect 235418 490046 265958 490102
rect 266014 490046 266082 490102
rect 266138 490046 296678 490102
rect 296734 490046 296802 490102
rect 296858 490046 327398 490102
rect 327454 490046 327522 490102
rect 327578 490046 358118 490102
rect 358174 490046 358242 490102
rect 358298 490046 388838 490102
rect 388894 490046 388962 490102
rect 389018 490046 419558 490102
rect 419614 490046 419682 490102
rect 419738 490046 450278 490102
rect 450334 490046 450402 490102
rect 450458 490046 480998 490102
rect 481054 490046 481122 490102
rect 481178 490046 507250 490102
rect 507306 490046 507374 490102
rect 507430 490046 507498 490102
rect 507554 490046 507622 490102
rect 507678 490046 525250 490102
rect 525306 490046 525374 490102
rect 525430 490046 525498 490102
rect 525554 490046 525622 490102
rect 525678 490046 543250 490102
rect 543306 490046 543374 490102
rect 543430 490046 543498 490102
rect 543554 490046 543622 490102
rect 543678 490046 561250 490102
rect 561306 490046 561374 490102
rect 561430 490046 561498 490102
rect 561554 490046 561622 490102
rect 561678 490046 579250 490102
rect 579306 490046 579374 490102
rect 579430 490046 579498 490102
rect 579554 490046 579622 490102
rect 579678 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 3250 489978
rect 3306 489922 3374 489978
rect 3430 489922 3498 489978
rect 3554 489922 3622 489978
rect 3678 489922 21250 489978
rect 21306 489922 21374 489978
rect 21430 489922 21498 489978
rect 21554 489922 21622 489978
rect 21678 489922 39250 489978
rect 39306 489922 39374 489978
rect 39430 489922 39498 489978
rect 39554 489922 39622 489978
rect 39678 489922 57250 489978
rect 57306 489922 57374 489978
rect 57430 489922 57498 489978
rect 57554 489922 57622 489978
rect 57678 489922 75250 489978
rect 75306 489922 75374 489978
rect 75430 489922 75498 489978
rect 75554 489922 75622 489978
rect 75678 489922 93250 489978
rect 93306 489922 93374 489978
rect 93430 489922 93498 489978
rect 93554 489922 93622 489978
rect 93678 489922 111250 489978
rect 111306 489922 111374 489978
rect 111430 489922 111498 489978
rect 111554 489922 111622 489978
rect 111678 489922 129250 489978
rect 129306 489922 129374 489978
rect 129430 489922 129498 489978
rect 129554 489922 129622 489978
rect 129678 489922 147250 489978
rect 147306 489922 147374 489978
rect 147430 489922 147498 489978
rect 147554 489922 147622 489978
rect 147678 489922 165250 489978
rect 165306 489922 165374 489978
rect 165430 489922 165498 489978
rect 165554 489922 165622 489978
rect 165678 489922 183250 489978
rect 183306 489922 183374 489978
rect 183430 489922 183498 489978
rect 183554 489922 183622 489978
rect 183678 489922 201250 489978
rect 201306 489922 201374 489978
rect 201430 489922 201498 489978
rect 201554 489922 201622 489978
rect 201678 489922 204518 489978
rect 204574 489922 204642 489978
rect 204698 489922 235238 489978
rect 235294 489922 235362 489978
rect 235418 489922 265958 489978
rect 266014 489922 266082 489978
rect 266138 489922 296678 489978
rect 296734 489922 296802 489978
rect 296858 489922 327398 489978
rect 327454 489922 327522 489978
rect 327578 489922 358118 489978
rect 358174 489922 358242 489978
rect 358298 489922 388838 489978
rect 388894 489922 388962 489978
rect 389018 489922 419558 489978
rect 419614 489922 419682 489978
rect 419738 489922 450278 489978
rect 450334 489922 450402 489978
rect 450458 489922 480998 489978
rect 481054 489922 481122 489978
rect 481178 489922 507250 489978
rect 507306 489922 507374 489978
rect 507430 489922 507498 489978
rect 507554 489922 507622 489978
rect 507678 489922 525250 489978
rect 525306 489922 525374 489978
rect 525430 489922 525498 489978
rect 525554 489922 525622 489978
rect 525678 489922 543250 489978
rect 543306 489922 543374 489978
rect 543430 489922 543498 489978
rect 543554 489922 543622 489978
rect 543678 489922 561250 489978
rect 561306 489922 561374 489978
rect 561430 489922 561498 489978
rect 561554 489922 561622 489978
rect 561678 489922 579250 489978
rect 579306 489922 579374 489978
rect 579430 489922 579498 489978
rect 579554 489922 579622 489978
rect 579678 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 6970 478350
rect 7026 478294 7094 478350
rect 7150 478294 7218 478350
rect 7274 478294 7342 478350
rect 7398 478294 24970 478350
rect 25026 478294 25094 478350
rect 25150 478294 25218 478350
rect 25274 478294 25342 478350
rect 25398 478294 42970 478350
rect 43026 478294 43094 478350
rect 43150 478294 43218 478350
rect 43274 478294 43342 478350
rect 43398 478294 60970 478350
rect 61026 478294 61094 478350
rect 61150 478294 61218 478350
rect 61274 478294 61342 478350
rect 61398 478294 78970 478350
rect 79026 478294 79094 478350
rect 79150 478294 79218 478350
rect 79274 478294 79342 478350
rect 79398 478294 96970 478350
rect 97026 478294 97094 478350
rect 97150 478294 97218 478350
rect 97274 478294 97342 478350
rect 97398 478294 114970 478350
rect 115026 478294 115094 478350
rect 115150 478294 115218 478350
rect 115274 478294 115342 478350
rect 115398 478294 132970 478350
rect 133026 478294 133094 478350
rect 133150 478294 133218 478350
rect 133274 478294 133342 478350
rect 133398 478294 150970 478350
rect 151026 478294 151094 478350
rect 151150 478294 151218 478350
rect 151274 478294 151342 478350
rect 151398 478294 168970 478350
rect 169026 478294 169094 478350
rect 169150 478294 169218 478350
rect 169274 478294 169342 478350
rect 169398 478294 186970 478350
rect 187026 478294 187094 478350
rect 187150 478294 187218 478350
rect 187274 478294 187342 478350
rect 187398 478294 219878 478350
rect 219934 478294 220002 478350
rect 220058 478294 250598 478350
rect 250654 478294 250722 478350
rect 250778 478294 281318 478350
rect 281374 478294 281442 478350
rect 281498 478294 312038 478350
rect 312094 478294 312162 478350
rect 312218 478294 342758 478350
rect 342814 478294 342882 478350
rect 342938 478294 373478 478350
rect 373534 478294 373602 478350
rect 373658 478294 404198 478350
rect 404254 478294 404322 478350
rect 404378 478294 434918 478350
rect 434974 478294 435042 478350
rect 435098 478294 465638 478350
rect 465694 478294 465762 478350
rect 465818 478294 496358 478350
rect 496414 478294 496482 478350
rect 496538 478294 510970 478350
rect 511026 478294 511094 478350
rect 511150 478294 511218 478350
rect 511274 478294 511342 478350
rect 511398 478294 528970 478350
rect 529026 478294 529094 478350
rect 529150 478294 529218 478350
rect 529274 478294 529342 478350
rect 529398 478294 546970 478350
rect 547026 478294 547094 478350
rect 547150 478294 547218 478350
rect 547274 478294 547342 478350
rect 547398 478294 564970 478350
rect 565026 478294 565094 478350
rect 565150 478294 565218 478350
rect 565274 478294 565342 478350
rect 565398 478294 582970 478350
rect 583026 478294 583094 478350
rect 583150 478294 583218 478350
rect 583274 478294 583342 478350
rect 583398 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 6970 478226
rect 7026 478170 7094 478226
rect 7150 478170 7218 478226
rect 7274 478170 7342 478226
rect 7398 478170 24970 478226
rect 25026 478170 25094 478226
rect 25150 478170 25218 478226
rect 25274 478170 25342 478226
rect 25398 478170 42970 478226
rect 43026 478170 43094 478226
rect 43150 478170 43218 478226
rect 43274 478170 43342 478226
rect 43398 478170 60970 478226
rect 61026 478170 61094 478226
rect 61150 478170 61218 478226
rect 61274 478170 61342 478226
rect 61398 478170 78970 478226
rect 79026 478170 79094 478226
rect 79150 478170 79218 478226
rect 79274 478170 79342 478226
rect 79398 478170 96970 478226
rect 97026 478170 97094 478226
rect 97150 478170 97218 478226
rect 97274 478170 97342 478226
rect 97398 478170 114970 478226
rect 115026 478170 115094 478226
rect 115150 478170 115218 478226
rect 115274 478170 115342 478226
rect 115398 478170 132970 478226
rect 133026 478170 133094 478226
rect 133150 478170 133218 478226
rect 133274 478170 133342 478226
rect 133398 478170 150970 478226
rect 151026 478170 151094 478226
rect 151150 478170 151218 478226
rect 151274 478170 151342 478226
rect 151398 478170 168970 478226
rect 169026 478170 169094 478226
rect 169150 478170 169218 478226
rect 169274 478170 169342 478226
rect 169398 478170 186970 478226
rect 187026 478170 187094 478226
rect 187150 478170 187218 478226
rect 187274 478170 187342 478226
rect 187398 478170 219878 478226
rect 219934 478170 220002 478226
rect 220058 478170 250598 478226
rect 250654 478170 250722 478226
rect 250778 478170 281318 478226
rect 281374 478170 281442 478226
rect 281498 478170 312038 478226
rect 312094 478170 312162 478226
rect 312218 478170 342758 478226
rect 342814 478170 342882 478226
rect 342938 478170 373478 478226
rect 373534 478170 373602 478226
rect 373658 478170 404198 478226
rect 404254 478170 404322 478226
rect 404378 478170 434918 478226
rect 434974 478170 435042 478226
rect 435098 478170 465638 478226
rect 465694 478170 465762 478226
rect 465818 478170 496358 478226
rect 496414 478170 496482 478226
rect 496538 478170 510970 478226
rect 511026 478170 511094 478226
rect 511150 478170 511218 478226
rect 511274 478170 511342 478226
rect 511398 478170 528970 478226
rect 529026 478170 529094 478226
rect 529150 478170 529218 478226
rect 529274 478170 529342 478226
rect 529398 478170 546970 478226
rect 547026 478170 547094 478226
rect 547150 478170 547218 478226
rect 547274 478170 547342 478226
rect 547398 478170 564970 478226
rect 565026 478170 565094 478226
rect 565150 478170 565218 478226
rect 565274 478170 565342 478226
rect 565398 478170 582970 478226
rect 583026 478170 583094 478226
rect 583150 478170 583218 478226
rect 583274 478170 583342 478226
rect 583398 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 6970 478102
rect 7026 478046 7094 478102
rect 7150 478046 7218 478102
rect 7274 478046 7342 478102
rect 7398 478046 24970 478102
rect 25026 478046 25094 478102
rect 25150 478046 25218 478102
rect 25274 478046 25342 478102
rect 25398 478046 42970 478102
rect 43026 478046 43094 478102
rect 43150 478046 43218 478102
rect 43274 478046 43342 478102
rect 43398 478046 60970 478102
rect 61026 478046 61094 478102
rect 61150 478046 61218 478102
rect 61274 478046 61342 478102
rect 61398 478046 78970 478102
rect 79026 478046 79094 478102
rect 79150 478046 79218 478102
rect 79274 478046 79342 478102
rect 79398 478046 96970 478102
rect 97026 478046 97094 478102
rect 97150 478046 97218 478102
rect 97274 478046 97342 478102
rect 97398 478046 114970 478102
rect 115026 478046 115094 478102
rect 115150 478046 115218 478102
rect 115274 478046 115342 478102
rect 115398 478046 132970 478102
rect 133026 478046 133094 478102
rect 133150 478046 133218 478102
rect 133274 478046 133342 478102
rect 133398 478046 150970 478102
rect 151026 478046 151094 478102
rect 151150 478046 151218 478102
rect 151274 478046 151342 478102
rect 151398 478046 168970 478102
rect 169026 478046 169094 478102
rect 169150 478046 169218 478102
rect 169274 478046 169342 478102
rect 169398 478046 186970 478102
rect 187026 478046 187094 478102
rect 187150 478046 187218 478102
rect 187274 478046 187342 478102
rect 187398 478046 219878 478102
rect 219934 478046 220002 478102
rect 220058 478046 250598 478102
rect 250654 478046 250722 478102
rect 250778 478046 281318 478102
rect 281374 478046 281442 478102
rect 281498 478046 312038 478102
rect 312094 478046 312162 478102
rect 312218 478046 342758 478102
rect 342814 478046 342882 478102
rect 342938 478046 373478 478102
rect 373534 478046 373602 478102
rect 373658 478046 404198 478102
rect 404254 478046 404322 478102
rect 404378 478046 434918 478102
rect 434974 478046 435042 478102
rect 435098 478046 465638 478102
rect 465694 478046 465762 478102
rect 465818 478046 496358 478102
rect 496414 478046 496482 478102
rect 496538 478046 510970 478102
rect 511026 478046 511094 478102
rect 511150 478046 511218 478102
rect 511274 478046 511342 478102
rect 511398 478046 528970 478102
rect 529026 478046 529094 478102
rect 529150 478046 529218 478102
rect 529274 478046 529342 478102
rect 529398 478046 546970 478102
rect 547026 478046 547094 478102
rect 547150 478046 547218 478102
rect 547274 478046 547342 478102
rect 547398 478046 564970 478102
rect 565026 478046 565094 478102
rect 565150 478046 565218 478102
rect 565274 478046 565342 478102
rect 565398 478046 582970 478102
rect 583026 478046 583094 478102
rect 583150 478046 583218 478102
rect 583274 478046 583342 478102
rect 583398 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 6970 477978
rect 7026 477922 7094 477978
rect 7150 477922 7218 477978
rect 7274 477922 7342 477978
rect 7398 477922 24970 477978
rect 25026 477922 25094 477978
rect 25150 477922 25218 477978
rect 25274 477922 25342 477978
rect 25398 477922 42970 477978
rect 43026 477922 43094 477978
rect 43150 477922 43218 477978
rect 43274 477922 43342 477978
rect 43398 477922 60970 477978
rect 61026 477922 61094 477978
rect 61150 477922 61218 477978
rect 61274 477922 61342 477978
rect 61398 477922 78970 477978
rect 79026 477922 79094 477978
rect 79150 477922 79218 477978
rect 79274 477922 79342 477978
rect 79398 477922 96970 477978
rect 97026 477922 97094 477978
rect 97150 477922 97218 477978
rect 97274 477922 97342 477978
rect 97398 477922 114970 477978
rect 115026 477922 115094 477978
rect 115150 477922 115218 477978
rect 115274 477922 115342 477978
rect 115398 477922 132970 477978
rect 133026 477922 133094 477978
rect 133150 477922 133218 477978
rect 133274 477922 133342 477978
rect 133398 477922 150970 477978
rect 151026 477922 151094 477978
rect 151150 477922 151218 477978
rect 151274 477922 151342 477978
rect 151398 477922 168970 477978
rect 169026 477922 169094 477978
rect 169150 477922 169218 477978
rect 169274 477922 169342 477978
rect 169398 477922 186970 477978
rect 187026 477922 187094 477978
rect 187150 477922 187218 477978
rect 187274 477922 187342 477978
rect 187398 477922 219878 477978
rect 219934 477922 220002 477978
rect 220058 477922 250598 477978
rect 250654 477922 250722 477978
rect 250778 477922 281318 477978
rect 281374 477922 281442 477978
rect 281498 477922 312038 477978
rect 312094 477922 312162 477978
rect 312218 477922 342758 477978
rect 342814 477922 342882 477978
rect 342938 477922 373478 477978
rect 373534 477922 373602 477978
rect 373658 477922 404198 477978
rect 404254 477922 404322 477978
rect 404378 477922 434918 477978
rect 434974 477922 435042 477978
rect 435098 477922 465638 477978
rect 465694 477922 465762 477978
rect 465818 477922 496358 477978
rect 496414 477922 496482 477978
rect 496538 477922 510970 477978
rect 511026 477922 511094 477978
rect 511150 477922 511218 477978
rect 511274 477922 511342 477978
rect 511398 477922 528970 477978
rect 529026 477922 529094 477978
rect 529150 477922 529218 477978
rect 529274 477922 529342 477978
rect 529398 477922 546970 477978
rect 547026 477922 547094 477978
rect 547150 477922 547218 477978
rect 547274 477922 547342 477978
rect 547398 477922 564970 477978
rect 565026 477922 565094 477978
rect 565150 477922 565218 477978
rect 565274 477922 565342 477978
rect 565398 477922 582970 477978
rect 583026 477922 583094 477978
rect 583150 477922 583218 477978
rect 583274 477922 583342 477978
rect 583398 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 3250 472350
rect 3306 472294 3374 472350
rect 3430 472294 3498 472350
rect 3554 472294 3622 472350
rect 3678 472294 21250 472350
rect 21306 472294 21374 472350
rect 21430 472294 21498 472350
rect 21554 472294 21622 472350
rect 21678 472294 39250 472350
rect 39306 472294 39374 472350
rect 39430 472294 39498 472350
rect 39554 472294 39622 472350
rect 39678 472294 57250 472350
rect 57306 472294 57374 472350
rect 57430 472294 57498 472350
rect 57554 472294 57622 472350
rect 57678 472294 75250 472350
rect 75306 472294 75374 472350
rect 75430 472294 75498 472350
rect 75554 472294 75622 472350
rect 75678 472294 93250 472350
rect 93306 472294 93374 472350
rect 93430 472294 93498 472350
rect 93554 472294 93622 472350
rect 93678 472294 111250 472350
rect 111306 472294 111374 472350
rect 111430 472294 111498 472350
rect 111554 472294 111622 472350
rect 111678 472294 129250 472350
rect 129306 472294 129374 472350
rect 129430 472294 129498 472350
rect 129554 472294 129622 472350
rect 129678 472294 147250 472350
rect 147306 472294 147374 472350
rect 147430 472294 147498 472350
rect 147554 472294 147622 472350
rect 147678 472294 165250 472350
rect 165306 472294 165374 472350
rect 165430 472294 165498 472350
rect 165554 472294 165622 472350
rect 165678 472294 183250 472350
rect 183306 472294 183374 472350
rect 183430 472294 183498 472350
rect 183554 472294 183622 472350
rect 183678 472294 201250 472350
rect 201306 472294 201374 472350
rect 201430 472294 201498 472350
rect 201554 472294 201622 472350
rect 201678 472294 204518 472350
rect 204574 472294 204642 472350
rect 204698 472294 235238 472350
rect 235294 472294 235362 472350
rect 235418 472294 265958 472350
rect 266014 472294 266082 472350
rect 266138 472294 296678 472350
rect 296734 472294 296802 472350
rect 296858 472294 327398 472350
rect 327454 472294 327522 472350
rect 327578 472294 358118 472350
rect 358174 472294 358242 472350
rect 358298 472294 388838 472350
rect 388894 472294 388962 472350
rect 389018 472294 419558 472350
rect 419614 472294 419682 472350
rect 419738 472294 450278 472350
rect 450334 472294 450402 472350
rect 450458 472294 480998 472350
rect 481054 472294 481122 472350
rect 481178 472294 507250 472350
rect 507306 472294 507374 472350
rect 507430 472294 507498 472350
rect 507554 472294 507622 472350
rect 507678 472294 525250 472350
rect 525306 472294 525374 472350
rect 525430 472294 525498 472350
rect 525554 472294 525622 472350
rect 525678 472294 543250 472350
rect 543306 472294 543374 472350
rect 543430 472294 543498 472350
rect 543554 472294 543622 472350
rect 543678 472294 561250 472350
rect 561306 472294 561374 472350
rect 561430 472294 561498 472350
rect 561554 472294 561622 472350
rect 561678 472294 579250 472350
rect 579306 472294 579374 472350
rect 579430 472294 579498 472350
rect 579554 472294 579622 472350
rect 579678 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 3250 472226
rect 3306 472170 3374 472226
rect 3430 472170 3498 472226
rect 3554 472170 3622 472226
rect 3678 472170 21250 472226
rect 21306 472170 21374 472226
rect 21430 472170 21498 472226
rect 21554 472170 21622 472226
rect 21678 472170 39250 472226
rect 39306 472170 39374 472226
rect 39430 472170 39498 472226
rect 39554 472170 39622 472226
rect 39678 472170 57250 472226
rect 57306 472170 57374 472226
rect 57430 472170 57498 472226
rect 57554 472170 57622 472226
rect 57678 472170 75250 472226
rect 75306 472170 75374 472226
rect 75430 472170 75498 472226
rect 75554 472170 75622 472226
rect 75678 472170 93250 472226
rect 93306 472170 93374 472226
rect 93430 472170 93498 472226
rect 93554 472170 93622 472226
rect 93678 472170 111250 472226
rect 111306 472170 111374 472226
rect 111430 472170 111498 472226
rect 111554 472170 111622 472226
rect 111678 472170 129250 472226
rect 129306 472170 129374 472226
rect 129430 472170 129498 472226
rect 129554 472170 129622 472226
rect 129678 472170 147250 472226
rect 147306 472170 147374 472226
rect 147430 472170 147498 472226
rect 147554 472170 147622 472226
rect 147678 472170 165250 472226
rect 165306 472170 165374 472226
rect 165430 472170 165498 472226
rect 165554 472170 165622 472226
rect 165678 472170 183250 472226
rect 183306 472170 183374 472226
rect 183430 472170 183498 472226
rect 183554 472170 183622 472226
rect 183678 472170 201250 472226
rect 201306 472170 201374 472226
rect 201430 472170 201498 472226
rect 201554 472170 201622 472226
rect 201678 472170 204518 472226
rect 204574 472170 204642 472226
rect 204698 472170 235238 472226
rect 235294 472170 235362 472226
rect 235418 472170 265958 472226
rect 266014 472170 266082 472226
rect 266138 472170 296678 472226
rect 296734 472170 296802 472226
rect 296858 472170 327398 472226
rect 327454 472170 327522 472226
rect 327578 472170 358118 472226
rect 358174 472170 358242 472226
rect 358298 472170 388838 472226
rect 388894 472170 388962 472226
rect 389018 472170 419558 472226
rect 419614 472170 419682 472226
rect 419738 472170 450278 472226
rect 450334 472170 450402 472226
rect 450458 472170 480998 472226
rect 481054 472170 481122 472226
rect 481178 472170 507250 472226
rect 507306 472170 507374 472226
rect 507430 472170 507498 472226
rect 507554 472170 507622 472226
rect 507678 472170 525250 472226
rect 525306 472170 525374 472226
rect 525430 472170 525498 472226
rect 525554 472170 525622 472226
rect 525678 472170 543250 472226
rect 543306 472170 543374 472226
rect 543430 472170 543498 472226
rect 543554 472170 543622 472226
rect 543678 472170 561250 472226
rect 561306 472170 561374 472226
rect 561430 472170 561498 472226
rect 561554 472170 561622 472226
rect 561678 472170 579250 472226
rect 579306 472170 579374 472226
rect 579430 472170 579498 472226
rect 579554 472170 579622 472226
rect 579678 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 3250 472102
rect 3306 472046 3374 472102
rect 3430 472046 3498 472102
rect 3554 472046 3622 472102
rect 3678 472046 21250 472102
rect 21306 472046 21374 472102
rect 21430 472046 21498 472102
rect 21554 472046 21622 472102
rect 21678 472046 39250 472102
rect 39306 472046 39374 472102
rect 39430 472046 39498 472102
rect 39554 472046 39622 472102
rect 39678 472046 57250 472102
rect 57306 472046 57374 472102
rect 57430 472046 57498 472102
rect 57554 472046 57622 472102
rect 57678 472046 75250 472102
rect 75306 472046 75374 472102
rect 75430 472046 75498 472102
rect 75554 472046 75622 472102
rect 75678 472046 93250 472102
rect 93306 472046 93374 472102
rect 93430 472046 93498 472102
rect 93554 472046 93622 472102
rect 93678 472046 111250 472102
rect 111306 472046 111374 472102
rect 111430 472046 111498 472102
rect 111554 472046 111622 472102
rect 111678 472046 129250 472102
rect 129306 472046 129374 472102
rect 129430 472046 129498 472102
rect 129554 472046 129622 472102
rect 129678 472046 147250 472102
rect 147306 472046 147374 472102
rect 147430 472046 147498 472102
rect 147554 472046 147622 472102
rect 147678 472046 165250 472102
rect 165306 472046 165374 472102
rect 165430 472046 165498 472102
rect 165554 472046 165622 472102
rect 165678 472046 183250 472102
rect 183306 472046 183374 472102
rect 183430 472046 183498 472102
rect 183554 472046 183622 472102
rect 183678 472046 201250 472102
rect 201306 472046 201374 472102
rect 201430 472046 201498 472102
rect 201554 472046 201622 472102
rect 201678 472046 204518 472102
rect 204574 472046 204642 472102
rect 204698 472046 235238 472102
rect 235294 472046 235362 472102
rect 235418 472046 265958 472102
rect 266014 472046 266082 472102
rect 266138 472046 296678 472102
rect 296734 472046 296802 472102
rect 296858 472046 327398 472102
rect 327454 472046 327522 472102
rect 327578 472046 358118 472102
rect 358174 472046 358242 472102
rect 358298 472046 388838 472102
rect 388894 472046 388962 472102
rect 389018 472046 419558 472102
rect 419614 472046 419682 472102
rect 419738 472046 450278 472102
rect 450334 472046 450402 472102
rect 450458 472046 480998 472102
rect 481054 472046 481122 472102
rect 481178 472046 507250 472102
rect 507306 472046 507374 472102
rect 507430 472046 507498 472102
rect 507554 472046 507622 472102
rect 507678 472046 525250 472102
rect 525306 472046 525374 472102
rect 525430 472046 525498 472102
rect 525554 472046 525622 472102
rect 525678 472046 543250 472102
rect 543306 472046 543374 472102
rect 543430 472046 543498 472102
rect 543554 472046 543622 472102
rect 543678 472046 561250 472102
rect 561306 472046 561374 472102
rect 561430 472046 561498 472102
rect 561554 472046 561622 472102
rect 561678 472046 579250 472102
rect 579306 472046 579374 472102
rect 579430 472046 579498 472102
rect 579554 472046 579622 472102
rect 579678 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 3250 471978
rect 3306 471922 3374 471978
rect 3430 471922 3498 471978
rect 3554 471922 3622 471978
rect 3678 471922 21250 471978
rect 21306 471922 21374 471978
rect 21430 471922 21498 471978
rect 21554 471922 21622 471978
rect 21678 471922 39250 471978
rect 39306 471922 39374 471978
rect 39430 471922 39498 471978
rect 39554 471922 39622 471978
rect 39678 471922 57250 471978
rect 57306 471922 57374 471978
rect 57430 471922 57498 471978
rect 57554 471922 57622 471978
rect 57678 471922 75250 471978
rect 75306 471922 75374 471978
rect 75430 471922 75498 471978
rect 75554 471922 75622 471978
rect 75678 471922 93250 471978
rect 93306 471922 93374 471978
rect 93430 471922 93498 471978
rect 93554 471922 93622 471978
rect 93678 471922 111250 471978
rect 111306 471922 111374 471978
rect 111430 471922 111498 471978
rect 111554 471922 111622 471978
rect 111678 471922 129250 471978
rect 129306 471922 129374 471978
rect 129430 471922 129498 471978
rect 129554 471922 129622 471978
rect 129678 471922 147250 471978
rect 147306 471922 147374 471978
rect 147430 471922 147498 471978
rect 147554 471922 147622 471978
rect 147678 471922 165250 471978
rect 165306 471922 165374 471978
rect 165430 471922 165498 471978
rect 165554 471922 165622 471978
rect 165678 471922 183250 471978
rect 183306 471922 183374 471978
rect 183430 471922 183498 471978
rect 183554 471922 183622 471978
rect 183678 471922 201250 471978
rect 201306 471922 201374 471978
rect 201430 471922 201498 471978
rect 201554 471922 201622 471978
rect 201678 471922 204518 471978
rect 204574 471922 204642 471978
rect 204698 471922 235238 471978
rect 235294 471922 235362 471978
rect 235418 471922 265958 471978
rect 266014 471922 266082 471978
rect 266138 471922 296678 471978
rect 296734 471922 296802 471978
rect 296858 471922 327398 471978
rect 327454 471922 327522 471978
rect 327578 471922 358118 471978
rect 358174 471922 358242 471978
rect 358298 471922 388838 471978
rect 388894 471922 388962 471978
rect 389018 471922 419558 471978
rect 419614 471922 419682 471978
rect 419738 471922 450278 471978
rect 450334 471922 450402 471978
rect 450458 471922 480998 471978
rect 481054 471922 481122 471978
rect 481178 471922 507250 471978
rect 507306 471922 507374 471978
rect 507430 471922 507498 471978
rect 507554 471922 507622 471978
rect 507678 471922 525250 471978
rect 525306 471922 525374 471978
rect 525430 471922 525498 471978
rect 525554 471922 525622 471978
rect 525678 471922 543250 471978
rect 543306 471922 543374 471978
rect 543430 471922 543498 471978
rect 543554 471922 543622 471978
rect 543678 471922 561250 471978
rect 561306 471922 561374 471978
rect 561430 471922 561498 471978
rect 561554 471922 561622 471978
rect 561678 471922 579250 471978
rect 579306 471922 579374 471978
rect 579430 471922 579498 471978
rect 579554 471922 579622 471978
rect 579678 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 6970 460350
rect 7026 460294 7094 460350
rect 7150 460294 7218 460350
rect 7274 460294 7342 460350
rect 7398 460294 24970 460350
rect 25026 460294 25094 460350
rect 25150 460294 25218 460350
rect 25274 460294 25342 460350
rect 25398 460294 42970 460350
rect 43026 460294 43094 460350
rect 43150 460294 43218 460350
rect 43274 460294 43342 460350
rect 43398 460294 60970 460350
rect 61026 460294 61094 460350
rect 61150 460294 61218 460350
rect 61274 460294 61342 460350
rect 61398 460294 78970 460350
rect 79026 460294 79094 460350
rect 79150 460294 79218 460350
rect 79274 460294 79342 460350
rect 79398 460294 96970 460350
rect 97026 460294 97094 460350
rect 97150 460294 97218 460350
rect 97274 460294 97342 460350
rect 97398 460294 114970 460350
rect 115026 460294 115094 460350
rect 115150 460294 115218 460350
rect 115274 460294 115342 460350
rect 115398 460294 132970 460350
rect 133026 460294 133094 460350
rect 133150 460294 133218 460350
rect 133274 460294 133342 460350
rect 133398 460294 150970 460350
rect 151026 460294 151094 460350
rect 151150 460294 151218 460350
rect 151274 460294 151342 460350
rect 151398 460294 168970 460350
rect 169026 460294 169094 460350
rect 169150 460294 169218 460350
rect 169274 460294 169342 460350
rect 169398 460294 186970 460350
rect 187026 460294 187094 460350
rect 187150 460294 187218 460350
rect 187274 460294 187342 460350
rect 187398 460294 219878 460350
rect 219934 460294 220002 460350
rect 220058 460294 250598 460350
rect 250654 460294 250722 460350
rect 250778 460294 281318 460350
rect 281374 460294 281442 460350
rect 281498 460294 312038 460350
rect 312094 460294 312162 460350
rect 312218 460294 342758 460350
rect 342814 460294 342882 460350
rect 342938 460294 373478 460350
rect 373534 460294 373602 460350
rect 373658 460294 404198 460350
rect 404254 460294 404322 460350
rect 404378 460294 434918 460350
rect 434974 460294 435042 460350
rect 435098 460294 465638 460350
rect 465694 460294 465762 460350
rect 465818 460294 496358 460350
rect 496414 460294 496482 460350
rect 496538 460294 510970 460350
rect 511026 460294 511094 460350
rect 511150 460294 511218 460350
rect 511274 460294 511342 460350
rect 511398 460294 528970 460350
rect 529026 460294 529094 460350
rect 529150 460294 529218 460350
rect 529274 460294 529342 460350
rect 529398 460294 546970 460350
rect 547026 460294 547094 460350
rect 547150 460294 547218 460350
rect 547274 460294 547342 460350
rect 547398 460294 564970 460350
rect 565026 460294 565094 460350
rect 565150 460294 565218 460350
rect 565274 460294 565342 460350
rect 565398 460294 582970 460350
rect 583026 460294 583094 460350
rect 583150 460294 583218 460350
rect 583274 460294 583342 460350
rect 583398 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 6970 460226
rect 7026 460170 7094 460226
rect 7150 460170 7218 460226
rect 7274 460170 7342 460226
rect 7398 460170 24970 460226
rect 25026 460170 25094 460226
rect 25150 460170 25218 460226
rect 25274 460170 25342 460226
rect 25398 460170 42970 460226
rect 43026 460170 43094 460226
rect 43150 460170 43218 460226
rect 43274 460170 43342 460226
rect 43398 460170 60970 460226
rect 61026 460170 61094 460226
rect 61150 460170 61218 460226
rect 61274 460170 61342 460226
rect 61398 460170 78970 460226
rect 79026 460170 79094 460226
rect 79150 460170 79218 460226
rect 79274 460170 79342 460226
rect 79398 460170 96970 460226
rect 97026 460170 97094 460226
rect 97150 460170 97218 460226
rect 97274 460170 97342 460226
rect 97398 460170 114970 460226
rect 115026 460170 115094 460226
rect 115150 460170 115218 460226
rect 115274 460170 115342 460226
rect 115398 460170 132970 460226
rect 133026 460170 133094 460226
rect 133150 460170 133218 460226
rect 133274 460170 133342 460226
rect 133398 460170 150970 460226
rect 151026 460170 151094 460226
rect 151150 460170 151218 460226
rect 151274 460170 151342 460226
rect 151398 460170 168970 460226
rect 169026 460170 169094 460226
rect 169150 460170 169218 460226
rect 169274 460170 169342 460226
rect 169398 460170 186970 460226
rect 187026 460170 187094 460226
rect 187150 460170 187218 460226
rect 187274 460170 187342 460226
rect 187398 460170 219878 460226
rect 219934 460170 220002 460226
rect 220058 460170 250598 460226
rect 250654 460170 250722 460226
rect 250778 460170 281318 460226
rect 281374 460170 281442 460226
rect 281498 460170 312038 460226
rect 312094 460170 312162 460226
rect 312218 460170 342758 460226
rect 342814 460170 342882 460226
rect 342938 460170 373478 460226
rect 373534 460170 373602 460226
rect 373658 460170 404198 460226
rect 404254 460170 404322 460226
rect 404378 460170 434918 460226
rect 434974 460170 435042 460226
rect 435098 460170 465638 460226
rect 465694 460170 465762 460226
rect 465818 460170 496358 460226
rect 496414 460170 496482 460226
rect 496538 460170 510970 460226
rect 511026 460170 511094 460226
rect 511150 460170 511218 460226
rect 511274 460170 511342 460226
rect 511398 460170 528970 460226
rect 529026 460170 529094 460226
rect 529150 460170 529218 460226
rect 529274 460170 529342 460226
rect 529398 460170 546970 460226
rect 547026 460170 547094 460226
rect 547150 460170 547218 460226
rect 547274 460170 547342 460226
rect 547398 460170 564970 460226
rect 565026 460170 565094 460226
rect 565150 460170 565218 460226
rect 565274 460170 565342 460226
rect 565398 460170 582970 460226
rect 583026 460170 583094 460226
rect 583150 460170 583218 460226
rect 583274 460170 583342 460226
rect 583398 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 6970 460102
rect 7026 460046 7094 460102
rect 7150 460046 7218 460102
rect 7274 460046 7342 460102
rect 7398 460046 24970 460102
rect 25026 460046 25094 460102
rect 25150 460046 25218 460102
rect 25274 460046 25342 460102
rect 25398 460046 42970 460102
rect 43026 460046 43094 460102
rect 43150 460046 43218 460102
rect 43274 460046 43342 460102
rect 43398 460046 60970 460102
rect 61026 460046 61094 460102
rect 61150 460046 61218 460102
rect 61274 460046 61342 460102
rect 61398 460046 78970 460102
rect 79026 460046 79094 460102
rect 79150 460046 79218 460102
rect 79274 460046 79342 460102
rect 79398 460046 96970 460102
rect 97026 460046 97094 460102
rect 97150 460046 97218 460102
rect 97274 460046 97342 460102
rect 97398 460046 114970 460102
rect 115026 460046 115094 460102
rect 115150 460046 115218 460102
rect 115274 460046 115342 460102
rect 115398 460046 132970 460102
rect 133026 460046 133094 460102
rect 133150 460046 133218 460102
rect 133274 460046 133342 460102
rect 133398 460046 150970 460102
rect 151026 460046 151094 460102
rect 151150 460046 151218 460102
rect 151274 460046 151342 460102
rect 151398 460046 168970 460102
rect 169026 460046 169094 460102
rect 169150 460046 169218 460102
rect 169274 460046 169342 460102
rect 169398 460046 186970 460102
rect 187026 460046 187094 460102
rect 187150 460046 187218 460102
rect 187274 460046 187342 460102
rect 187398 460046 219878 460102
rect 219934 460046 220002 460102
rect 220058 460046 250598 460102
rect 250654 460046 250722 460102
rect 250778 460046 281318 460102
rect 281374 460046 281442 460102
rect 281498 460046 312038 460102
rect 312094 460046 312162 460102
rect 312218 460046 342758 460102
rect 342814 460046 342882 460102
rect 342938 460046 373478 460102
rect 373534 460046 373602 460102
rect 373658 460046 404198 460102
rect 404254 460046 404322 460102
rect 404378 460046 434918 460102
rect 434974 460046 435042 460102
rect 435098 460046 465638 460102
rect 465694 460046 465762 460102
rect 465818 460046 496358 460102
rect 496414 460046 496482 460102
rect 496538 460046 510970 460102
rect 511026 460046 511094 460102
rect 511150 460046 511218 460102
rect 511274 460046 511342 460102
rect 511398 460046 528970 460102
rect 529026 460046 529094 460102
rect 529150 460046 529218 460102
rect 529274 460046 529342 460102
rect 529398 460046 546970 460102
rect 547026 460046 547094 460102
rect 547150 460046 547218 460102
rect 547274 460046 547342 460102
rect 547398 460046 564970 460102
rect 565026 460046 565094 460102
rect 565150 460046 565218 460102
rect 565274 460046 565342 460102
rect 565398 460046 582970 460102
rect 583026 460046 583094 460102
rect 583150 460046 583218 460102
rect 583274 460046 583342 460102
rect 583398 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 6970 459978
rect 7026 459922 7094 459978
rect 7150 459922 7218 459978
rect 7274 459922 7342 459978
rect 7398 459922 24970 459978
rect 25026 459922 25094 459978
rect 25150 459922 25218 459978
rect 25274 459922 25342 459978
rect 25398 459922 42970 459978
rect 43026 459922 43094 459978
rect 43150 459922 43218 459978
rect 43274 459922 43342 459978
rect 43398 459922 60970 459978
rect 61026 459922 61094 459978
rect 61150 459922 61218 459978
rect 61274 459922 61342 459978
rect 61398 459922 78970 459978
rect 79026 459922 79094 459978
rect 79150 459922 79218 459978
rect 79274 459922 79342 459978
rect 79398 459922 96970 459978
rect 97026 459922 97094 459978
rect 97150 459922 97218 459978
rect 97274 459922 97342 459978
rect 97398 459922 114970 459978
rect 115026 459922 115094 459978
rect 115150 459922 115218 459978
rect 115274 459922 115342 459978
rect 115398 459922 132970 459978
rect 133026 459922 133094 459978
rect 133150 459922 133218 459978
rect 133274 459922 133342 459978
rect 133398 459922 150970 459978
rect 151026 459922 151094 459978
rect 151150 459922 151218 459978
rect 151274 459922 151342 459978
rect 151398 459922 168970 459978
rect 169026 459922 169094 459978
rect 169150 459922 169218 459978
rect 169274 459922 169342 459978
rect 169398 459922 186970 459978
rect 187026 459922 187094 459978
rect 187150 459922 187218 459978
rect 187274 459922 187342 459978
rect 187398 459922 219878 459978
rect 219934 459922 220002 459978
rect 220058 459922 250598 459978
rect 250654 459922 250722 459978
rect 250778 459922 281318 459978
rect 281374 459922 281442 459978
rect 281498 459922 312038 459978
rect 312094 459922 312162 459978
rect 312218 459922 342758 459978
rect 342814 459922 342882 459978
rect 342938 459922 373478 459978
rect 373534 459922 373602 459978
rect 373658 459922 404198 459978
rect 404254 459922 404322 459978
rect 404378 459922 434918 459978
rect 434974 459922 435042 459978
rect 435098 459922 465638 459978
rect 465694 459922 465762 459978
rect 465818 459922 496358 459978
rect 496414 459922 496482 459978
rect 496538 459922 510970 459978
rect 511026 459922 511094 459978
rect 511150 459922 511218 459978
rect 511274 459922 511342 459978
rect 511398 459922 528970 459978
rect 529026 459922 529094 459978
rect 529150 459922 529218 459978
rect 529274 459922 529342 459978
rect 529398 459922 546970 459978
rect 547026 459922 547094 459978
rect 547150 459922 547218 459978
rect 547274 459922 547342 459978
rect 547398 459922 564970 459978
rect 565026 459922 565094 459978
rect 565150 459922 565218 459978
rect 565274 459922 565342 459978
rect 565398 459922 582970 459978
rect 583026 459922 583094 459978
rect 583150 459922 583218 459978
rect 583274 459922 583342 459978
rect 583398 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 3250 454350
rect 3306 454294 3374 454350
rect 3430 454294 3498 454350
rect 3554 454294 3622 454350
rect 3678 454294 21250 454350
rect 21306 454294 21374 454350
rect 21430 454294 21498 454350
rect 21554 454294 21622 454350
rect 21678 454294 39250 454350
rect 39306 454294 39374 454350
rect 39430 454294 39498 454350
rect 39554 454294 39622 454350
rect 39678 454294 57250 454350
rect 57306 454294 57374 454350
rect 57430 454294 57498 454350
rect 57554 454294 57622 454350
rect 57678 454294 75250 454350
rect 75306 454294 75374 454350
rect 75430 454294 75498 454350
rect 75554 454294 75622 454350
rect 75678 454294 93250 454350
rect 93306 454294 93374 454350
rect 93430 454294 93498 454350
rect 93554 454294 93622 454350
rect 93678 454294 111250 454350
rect 111306 454294 111374 454350
rect 111430 454294 111498 454350
rect 111554 454294 111622 454350
rect 111678 454294 129250 454350
rect 129306 454294 129374 454350
rect 129430 454294 129498 454350
rect 129554 454294 129622 454350
rect 129678 454294 147250 454350
rect 147306 454294 147374 454350
rect 147430 454294 147498 454350
rect 147554 454294 147622 454350
rect 147678 454294 165250 454350
rect 165306 454294 165374 454350
rect 165430 454294 165498 454350
rect 165554 454294 165622 454350
rect 165678 454294 183250 454350
rect 183306 454294 183374 454350
rect 183430 454294 183498 454350
rect 183554 454294 183622 454350
rect 183678 454294 201250 454350
rect 201306 454294 201374 454350
rect 201430 454294 201498 454350
rect 201554 454294 201622 454350
rect 201678 454294 204518 454350
rect 204574 454294 204642 454350
rect 204698 454294 235238 454350
rect 235294 454294 235362 454350
rect 235418 454294 265958 454350
rect 266014 454294 266082 454350
rect 266138 454294 296678 454350
rect 296734 454294 296802 454350
rect 296858 454294 327398 454350
rect 327454 454294 327522 454350
rect 327578 454294 358118 454350
rect 358174 454294 358242 454350
rect 358298 454294 388838 454350
rect 388894 454294 388962 454350
rect 389018 454294 419558 454350
rect 419614 454294 419682 454350
rect 419738 454294 450278 454350
rect 450334 454294 450402 454350
rect 450458 454294 480998 454350
rect 481054 454294 481122 454350
rect 481178 454294 507250 454350
rect 507306 454294 507374 454350
rect 507430 454294 507498 454350
rect 507554 454294 507622 454350
rect 507678 454294 525250 454350
rect 525306 454294 525374 454350
rect 525430 454294 525498 454350
rect 525554 454294 525622 454350
rect 525678 454294 543250 454350
rect 543306 454294 543374 454350
rect 543430 454294 543498 454350
rect 543554 454294 543622 454350
rect 543678 454294 561250 454350
rect 561306 454294 561374 454350
rect 561430 454294 561498 454350
rect 561554 454294 561622 454350
rect 561678 454294 579250 454350
rect 579306 454294 579374 454350
rect 579430 454294 579498 454350
rect 579554 454294 579622 454350
rect 579678 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 3250 454226
rect 3306 454170 3374 454226
rect 3430 454170 3498 454226
rect 3554 454170 3622 454226
rect 3678 454170 21250 454226
rect 21306 454170 21374 454226
rect 21430 454170 21498 454226
rect 21554 454170 21622 454226
rect 21678 454170 39250 454226
rect 39306 454170 39374 454226
rect 39430 454170 39498 454226
rect 39554 454170 39622 454226
rect 39678 454170 57250 454226
rect 57306 454170 57374 454226
rect 57430 454170 57498 454226
rect 57554 454170 57622 454226
rect 57678 454170 75250 454226
rect 75306 454170 75374 454226
rect 75430 454170 75498 454226
rect 75554 454170 75622 454226
rect 75678 454170 93250 454226
rect 93306 454170 93374 454226
rect 93430 454170 93498 454226
rect 93554 454170 93622 454226
rect 93678 454170 111250 454226
rect 111306 454170 111374 454226
rect 111430 454170 111498 454226
rect 111554 454170 111622 454226
rect 111678 454170 129250 454226
rect 129306 454170 129374 454226
rect 129430 454170 129498 454226
rect 129554 454170 129622 454226
rect 129678 454170 147250 454226
rect 147306 454170 147374 454226
rect 147430 454170 147498 454226
rect 147554 454170 147622 454226
rect 147678 454170 165250 454226
rect 165306 454170 165374 454226
rect 165430 454170 165498 454226
rect 165554 454170 165622 454226
rect 165678 454170 183250 454226
rect 183306 454170 183374 454226
rect 183430 454170 183498 454226
rect 183554 454170 183622 454226
rect 183678 454170 201250 454226
rect 201306 454170 201374 454226
rect 201430 454170 201498 454226
rect 201554 454170 201622 454226
rect 201678 454170 204518 454226
rect 204574 454170 204642 454226
rect 204698 454170 235238 454226
rect 235294 454170 235362 454226
rect 235418 454170 265958 454226
rect 266014 454170 266082 454226
rect 266138 454170 296678 454226
rect 296734 454170 296802 454226
rect 296858 454170 327398 454226
rect 327454 454170 327522 454226
rect 327578 454170 358118 454226
rect 358174 454170 358242 454226
rect 358298 454170 388838 454226
rect 388894 454170 388962 454226
rect 389018 454170 419558 454226
rect 419614 454170 419682 454226
rect 419738 454170 450278 454226
rect 450334 454170 450402 454226
rect 450458 454170 480998 454226
rect 481054 454170 481122 454226
rect 481178 454170 507250 454226
rect 507306 454170 507374 454226
rect 507430 454170 507498 454226
rect 507554 454170 507622 454226
rect 507678 454170 525250 454226
rect 525306 454170 525374 454226
rect 525430 454170 525498 454226
rect 525554 454170 525622 454226
rect 525678 454170 543250 454226
rect 543306 454170 543374 454226
rect 543430 454170 543498 454226
rect 543554 454170 543622 454226
rect 543678 454170 561250 454226
rect 561306 454170 561374 454226
rect 561430 454170 561498 454226
rect 561554 454170 561622 454226
rect 561678 454170 579250 454226
rect 579306 454170 579374 454226
rect 579430 454170 579498 454226
rect 579554 454170 579622 454226
rect 579678 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 3250 454102
rect 3306 454046 3374 454102
rect 3430 454046 3498 454102
rect 3554 454046 3622 454102
rect 3678 454046 21250 454102
rect 21306 454046 21374 454102
rect 21430 454046 21498 454102
rect 21554 454046 21622 454102
rect 21678 454046 39250 454102
rect 39306 454046 39374 454102
rect 39430 454046 39498 454102
rect 39554 454046 39622 454102
rect 39678 454046 57250 454102
rect 57306 454046 57374 454102
rect 57430 454046 57498 454102
rect 57554 454046 57622 454102
rect 57678 454046 75250 454102
rect 75306 454046 75374 454102
rect 75430 454046 75498 454102
rect 75554 454046 75622 454102
rect 75678 454046 93250 454102
rect 93306 454046 93374 454102
rect 93430 454046 93498 454102
rect 93554 454046 93622 454102
rect 93678 454046 111250 454102
rect 111306 454046 111374 454102
rect 111430 454046 111498 454102
rect 111554 454046 111622 454102
rect 111678 454046 129250 454102
rect 129306 454046 129374 454102
rect 129430 454046 129498 454102
rect 129554 454046 129622 454102
rect 129678 454046 147250 454102
rect 147306 454046 147374 454102
rect 147430 454046 147498 454102
rect 147554 454046 147622 454102
rect 147678 454046 165250 454102
rect 165306 454046 165374 454102
rect 165430 454046 165498 454102
rect 165554 454046 165622 454102
rect 165678 454046 183250 454102
rect 183306 454046 183374 454102
rect 183430 454046 183498 454102
rect 183554 454046 183622 454102
rect 183678 454046 201250 454102
rect 201306 454046 201374 454102
rect 201430 454046 201498 454102
rect 201554 454046 201622 454102
rect 201678 454046 204518 454102
rect 204574 454046 204642 454102
rect 204698 454046 235238 454102
rect 235294 454046 235362 454102
rect 235418 454046 265958 454102
rect 266014 454046 266082 454102
rect 266138 454046 296678 454102
rect 296734 454046 296802 454102
rect 296858 454046 327398 454102
rect 327454 454046 327522 454102
rect 327578 454046 358118 454102
rect 358174 454046 358242 454102
rect 358298 454046 388838 454102
rect 388894 454046 388962 454102
rect 389018 454046 419558 454102
rect 419614 454046 419682 454102
rect 419738 454046 450278 454102
rect 450334 454046 450402 454102
rect 450458 454046 480998 454102
rect 481054 454046 481122 454102
rect 481178 454046 507250 454102
rect 507306 454046 507374 454102
rect 507430 454046 507498 454102
rect 507554 454046 507622 454102
rect 507678 454046 525250 454102
rect 525306 454046 525374 454102
rect 525430 454046 525498 454102
rect 525554 454046 525622 454102
rect 525678 454046 543250 454102
rect 543306 454046 543374 454102
rect 543430 454046 543498 454102
rect 543554 454046 543622 454102
rect 543678 454046 561250 454102
rect 561306 454046 561374 454102
rect 561430 454046 561498 454102
rect 561554 454046 561622 454102
rect 561678 454046 579250 454102
rect 579306 454046 579374 454102
rect 579430 454046 579498 454102
rect 579554 454046 579622 454102
rect 579678 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 3250 453978
rect 3306 453922 3374 453978
rect 3430 453922 3498 453978
rect 3554 453922 3622 453978
rect 3678 453922 21250 453978
rect 21306 453922 21374 453978
rect 21430 453922 21498 453978
rect 21554 453922 21622 453978
rect 21678 453922 39250 453978
rect 39306 453922 39374 453978
rect 39430 453922 39498 453978
rect 39554 453922 39622 453978
rect 39678 453922 57250 453978
rect 57306 453922 57374 453978
rect 57430 453922 57498 453978
rect 57554 453922 57622 453978
rect 57678 453922 75250 453978
rect 75306 453922 75374 453978
rect 75430 453922 75498 453978
rect 75554 453922 75622 453978
rect 75678 453922 93250 453978
rect 93306 453922 93374 453978
rect 93430 453922 93498 453978
rect 93554 453922 93622 453978
rect 93678 453922 111250 453978
rect 111306 453922 111374 453978
rect 111430 453922 111498 453978
rect 111554 453922 111622 453978
rect 111678 453922 129250 453978
rect 129306 453922 129374 453978
rect 129430 453922 129498 453978
rect 129554 453922 129622 453978
rect 129678 453922 147250 453978
rect 147306 453922 147374 453978
rect 147430 453922 147498 453978
rect 147554 453922 147622 453978
rect 147678 453922 165250 453978
rect 165306 453922 165374 453978
rect 165430 453922 165498 453978
rect 165554 453922 165622 453978
rect 165678 453922 183250 453978
rect 183306 453922 183374 453978
rect 183430 453922 183498 453978
rect 183554 453922 183622 453978
rect 183678 453922 201250 453978
rect 201306 453922 201374 453978
rect 201430 453922 201498 453978
rect 201554 453922 201622 453978
rect 201678 453922 204518 453978
rect 204574 453922 204642 453978
rect 204698 453922 235238 453978
rect 235294 453922 235362 453978
rect 235418 453922 265958 453978
rect 266014 453922 266082 453978
rect 266138 453922 296678 453978
rect 296734 453922 296802 453978
rect 296858 453922 327398 453978
rect 327454 453922 327522 453978
rect 327578 453922 358118 453978
rect 358174 453922 358242 453978
rect 358298 453922 388838 453978
rect 388894 453922 388962 453978
rect 389018 453922 419558 453978
rect 419614 453922 419682 453978
rect 419738 453922 450278 453978
rect 450334 453922 450402 453978
rect 450458 453922 480998 453978
rect 481054 453922 481122 453978
rect 481178 453922 507250 453978
rect 507306 453922 507374 453978
rect 507430 453922 507498 453978
rect 507554 453922 507622 453978
rect 507678 453922 525250 453978
rect 525306 453922 525374 453978
rect 525430 453922 525498 453978
rect 525554 453922 525622 453978
rect 525678 453922 543250 453978
rect 543306 453922 543374 453978
rect 543430 453922 543498 453978
rect 543554 453922 543622 453978
rect 543678 453922 561250 453978
rect 561306 453922 561374 453978
rect 561430 453922 561498 453978
rect 561554 453922 561622 453978
rect 561678 453922 579250 453978
rect 579306 453922 579374 453978
rect 579430 453922 579498 453978
rect 579554 453922 579622 453978
rect 579678 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 6970 442350
rect 7026 442294 7094 442350
rect 7150 442294 7218 442350
rect 7274 442294 7342 442350
rect 7398 442294 24970 442350
rect 25026 442294 25094 442350
rect 25150 442294 25218 442350
rect 25274 442294 25342 442350
rect 25398 442294 42970 442350
rect 43026 442294 43094 442350
rect 43150 442294 43218 442350
rect 43274 442294 43342 442350
rect 43398 442294 60970 442350
rect 61026 442294 61094 442350
rect 61150 442294 61218 442350
rect 61274 442294 61342 442350
rect 61398 442294 78970 442350
rect 79026 442294 79094 442350
rect 79150 442294 79218 442350
rect 79274 442294 79342 442350
rect 79398 442294 96970 442350
rect 97026 442294 97094 442350
rect 97150 442294 97218 442350
rect 97274 442294 97342 442350
rect 97398 442294 114970 442350
rect 115026 442294 115094 442350
rect 115150 442294 115218 442350
rect 115274 442294 115342 442350
rect 115398 442294 132970 442350
rect 133026 442294 133094 442350
rect 133150 442294 133218 442350
rect 133274 442294 133342 442350
rect 133398 442294 150970 442350
rect 151026 442294 151094 442350
rect 151150 442294 151218 442350
rect 151274 442294 151342 442350
rect 151398 442294 168970 442350
rect 169026 442294 169094 442350
rect 169150 442294 169218 442350
rect 169274 442294 169342 442350
rect 169398 442294 186970 442350
rect 187026 442294 187094 442350
rect 187150 442294 187218 442350
rect 187274 442294 187342 442350
rect 187398 442294 219878 442350
rect 219934 442294 220002 442350
rect 220058 442294 250598 442350
rect 250654 442294 250722 442350
rect 250778 442294 281318 442350
rect 281374 442294 281442 442350
rect 281498 442294 312038 442350
rect 312094 442294 312162 442350
rect 312218 442294 342758 442350
rect 342814 442294 342882 442350
rect 342938 442294 373478 442350
rect 373534 442294 373602 442350
rect 373658 442294 404198 442350
rect 404254 442294 404322 442350
rect 404378 442294 434918 442350
rect 434974 442294 435042 442350
rect 435098 442294 465638 442350
rect 465694 442294 465762 442350
rect 465818 442294 496358 442350
rect 496414 442294 496482 442350
rect 496538 442294 510970 442350
rect 511026 442294 511094 442350
rect 511150 442294 511218 442350
rect 511274 442294 511342 442350
rect 511398 442294 528970 442350
rect 529026 442294 529094 442350
rect 529150 442294 529218 442350
rect 529274 442294 529342 442350
rect 529398 442294 546970 442350
rect 547026 442294 547094 442350
rect 547150 442294 547218 442350
rect 547274 442294 547342 442350
rect 547398 442294 564970 442350
rect 565026 442294 565094 442350
rect 565150 442294 565218 442350
rect 565274 442294 565342 442350
rect 565398 442294 582970 442350
rect 583026 442294 583094 442350
rect 583150 442294 583218 442350
rect 583274 442294 583342 442350
rect 583398 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 6970 442226
rect 7026 442170 7094 442226
rect 7150 442170 7218 442226
rect 7274 442170 7342 442226
rect 7398 442170 24970 442226
rect 25026 442170 25094 442226
rect 25150 442170 25218 442226
rect 25274 442170 25342 442226
rect 25398 442170 42970 442226
rect 43026 442170 43094 442226
rect 43150 442170 43218 442226
rect 43274 442170 43342 442226
rect 43398 442170 60970 442226
rect 61026 442170 61094 442226
rect 61150 442170 61218 442226
rect 61274 442170 61342 442226
rect 61398 442170 78970 442226
rect 79026 442170 79094 442226
rect 79150 442170 79218 442226
rect 79274 442170 79342 442226
rect 79398 442170 96970 442226
rect 97026 442170 97094 442226
rect 97150 442170 97218 442226
rect 97274 442170 97342 442226
rect 97398 442170 114970 442226
rect 115026 442170 115094 442226
rect 115150 442170 115218 442226
rect 115274 442170 115342 442226
rect 115398 442170 132970 442226
rect 133026 442170 133094 442226
rect 133150 442170 133218 442226
rect 133274 442170 133342 442226
rect 133398 442170 150970 442226
rect 151026 442170 151094 442226
rect 151150 442170 151218 442226
rect 151274 442170 151342 442226
rect 151398 442170 168970 442226
rect 169026 442170 169094 442226
rect 169150 442170 169218 442226
rect 169274 442170 169342 442226
rect 169398 442170 186970 442226
rect 187026 442170 187094 442226
rect 187150 442170 187218 442226
rect 187274 442170 187342 442226
rect 187398 442170 219878 442226
rect 219934 442170 220002 442226
rect 220058 442170 250598 442226
rect 250654 442170 250722 442226
rect 250778 442170 281318 442226
rect 281374 442170 281442 442226
rect 281498 442170 312038 442226
rect 312094 442170 312162 442226
rect 312218 442170 342758 442226
rect 342814 442170 342882 442226
rect 342938 442170 373478 442226
rect 373534 442170 373602 442226
rect 373658 442170 404198 442226
rect 404254 442170 404322 442226
rect 404378 442170 434918 442226
rect 434974 442170 435042 442226
rect 435098 442170 465638 442226
rect 465694 442170 465762 442226
rect 465818 442170 496358 442226
rect 496414 442170 496482 442226
rect 496538 442170 510970 442226
rect 511026 442170 511094 442226
rect 511150 442170 511218 442226
rect 511274 442170 511342 442226
rect 511398 442170 528970 442226
rect 529026 442170 529094 442226
rect 529150 442170 529218 442226
rect 529274 442170 529342 442226
rect 529398 442170 546970 442226
rect 547026 442170 547094 442226
rect 547150 442170 547218 442226
rect 547274 442170 547342 442226
rect 547398 442170 564970 442226
rect 565026 442170 565094 442226
rect 565150 442170 565218 442226
rect 565274 442170 565342 442226
rect 565398 442170 582970 442226
rect 583026 442170 583094 442226
rect 583150 442170 583218 442226
rect 583274 442170 583342 442226
rect 583398 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 6970 442102
rect 7026 442046 7094 442102
rect 7150 442046 7218 442102
rect 7274 442046 7342 442102
rect 7398 442046 24970 442102
rect 25026 442046 25094 442102
rect 25150 442046 25218 442102
rect 25274 442046 25342 442102
rect 25398 442046 42970 442102
rect 43026 442046 43094 442102
rect 43150 442046 43218 442102
rect 43274 442046 43342 442102
rect 43398 442046 60970 442102
rect 61026 442046 61094 442102
rect 61150 442046 61218 442102
rect 61274 442046 61342 442102
rect 61398 442046 78970 442102
rect 79026 442046 79094 442102
rect 79150 442046 79218 442102
rect 79274 442046 79342 442102
rect 79398 442046 96970 442102
rect 97026 442046 97094 442102
rect 97150 442046 97218 442102
rect 97274 442046 97342 442102
rect 97398 442046 114970 442102
rect 115026 442046 115094 442102
rect 115150 442046 115218 442102
rect 115274 442046 115342 442102
rect 115398 442046 132970 442102
rect 133026 442046 133094 442102
rect 133150 442046 133218 442102
rect 133274 442046 133342 442102
rect 133398 442046 150970 442102
rect 151026 442046 151094 442102
rect 151150 442046 151218 442102
rect 151274 442046 151342 442102
rect 151398 442046 168970 442102
rect 169026 442046 169094 442102
rect 169150 442046 169218 442102
rect 169274 442046 169342 442102
rect 169398 442046 186970 442102
rect 187026 442046 187094 442102
rect 187150 442046 187218 442102
rect 187274 442046 187342 442102
rect 187398 442046 219878 442102
rect 219934 442046 220002 442102
rect 220058 442046 250598 442102
rect 250654 442046 250722 442102
rect 250778 442046 281318 442102
rect 281374 442046 281442 442102
rect 281498 442046 312038 442102
rect 312094 442046 312162 442102
rect 312218 442046 342758 442102
rect 342814 442046 342882 442102
rect 342938 442046 373478 442102
rect 373534 442046 373602 442102
rect 373658 442046 404198 442102
rect 404254 442046 404322 442102
rect 404378 442046 434918 442102
rect 434974 442046 435042 442102
rect 435098 442046 465638 442102
rect 465694 442046 465762 442102
rect 465818 442046 496358 442102
rect 496414 442046 496482 442102
rect 496538 442046 510970 442102
rect 511026 442046 511094 442102
rect 511150 442046 511218 442102
rect 511274 442046 511342 442102
rect 511398 442046 528970 442102
rect 529026 442046 529094 442102
rect 529150 442046 529218 442102
rect 529274 442046 529342 442102
rect 529398 442046 546970 442102
rect 547026 442046 547094 442102
rect 547150 442046 547218 442102
rect 547274 442046 547342 442102
rect 547398 442046 564970 442102
rect 565026 442046 565094 442102
rect 565150 442046 565218 442102
rect 565274 442046 565342 442102
rect 565398 442046 582970 442102
rect 583026 442046 583094 442102
rect 583150 442046 583218 442102
rect 583274 442046 583342 442102
rect 583398 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 6970 441978
rect 7026 441922 7094 441978
rect 7150 441922 7218 441978
rect 7274 441922 7342 441978
rect 7398 441922 24970 441978
rect 25026 441922 25094 441978
rect 25150 441922 25218 441978
rect 25274 441922 25342 441978
rect 25398 441922 42970 441978
rect 43026 441922 43094 441978
rect 43150 441922 43218 441978
rect 43274 441922 43342 441978
rect 43398 441922 60970 441978
rect 61026 441922 61094 441978
rect 61150 441922 61218 441978
rect 61274 441922 61342 441978
rect 61398 441922 78970 441978
rect 79026 441922 79094 441978
rect 79150 441922 79218 441978
rect 79274 441922 79342 441978
rect 79398 441922 96970 441978
rect 97026 441922 97094 441978
rect 97150 441922 97218 441978
rect 97274 441922 97342 441978
rect 97398 441922 114970 441978
rect 115026 441922 115094 441978
rect 115150 441922 115218 441978
rect 115274 441922 115342 441978
rect 115398 441922 132970 441978
rect 133026 441922 133094 441978
rect 133150 441922 133218 441978
rect 133274 441922 133342 441978
rect 133398 441922 150970 441978
rect 151026 441922 151094 441978
rect 151150 441922 151218 441978
rect 151274 441922 151342 441978
rect 151398 441922 168970 441978
rect 169026 441922 169094 441978
rect 169150 441922 169218 441978
rect 169274 441922 169342 441978
rect 169398 441922 186970 441978
rect 187026 441922 187094 441978
rect 187150 441922 187218 441978
rect 187274 441922 187342 441978
rect 187398 441922 219878 441978
rect 219934 441922 220002 441978
rect 220058 441922 250598 441978
rect 250654 441922 250722 441978
rect 250778 441922 281318 441978
rect 281374 441922 281442 441978
rect 281498 441922 312038 441978
rect 312094 441922 312162 441978
rect 312218 441922 342758 441978
rect 342814 441922 342882 441978
rect 342938 441922 373478 441978
rect 373534 441922 373602 441978
rect 373658 441922 404198 441978
rect 404254 441922 404322 441978
rect 404378 441922 434918 441978
rect 434974 441922 435042 441978
rect 435098 441922 465638 441978
rect 465694 441922 465762 441978
rect 465818 441922 496358 441978
rect 496414 441922 496482 441978
rect 496538 441922 510970 441978
rect 511026 441922 511094 441978
rect 511150 441922 511218 441978
rect 511274 441922 511342 441978
rect 511398 441922 528970 441978
rect 529026 441922 529094 441978
rect 529150 441922 529218 441978
rect 529274 441922 529342 441978
rect 529398 441922 546970 441978
rect 547026 441922 547094 441978
rect 547150 441922 547218 441978
rect 547274 441922 547342 441978
rect 547398 441922 564970 441978
rect 565026 441922 565094 441978
rect 565150 441922 565218 441978
rect 565274 441922 565342 441978
rect 565398 441922 582970 441978
rect 583026 441922 583094 441978
rect 583150 441922 583218 441978
rect 583274 441922 583342 441978
rect 583398 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 3250 436350
rect 3306 436294 3374 436350
rect 3430 436294 3498 436350
rect 3554 436294 3622 436350
rect 3678 436294 21250 436350
rect 21306 436294 21374 436350
rect 21430 436294 21498 436350
rect 21554 436294 21622 436350
rect 21678 436294 39250 436350
rect 39306 436294 39374 436350
rect 39430 436294 39498 436350
rect 39554 436294 39622 436350
rect 39678 436294 57250 436350
rect 57306 436294 57374 436350
rect 57430 436294 57498 436350
rect 57554 436294 57622 436350
rect 57678 436294 75250 436350
rect 75306 436294 75374 436350
rect 75430 436294 75498 436350
rect 75554 436294 75622 436350
rect 75678 436294 93250 436350
rect 93306 436294 93374 436350
rect 93430 436294 93498 436350
rect 93554 436294 93622 436350
rect 93678 436294 111250 436350
rect 111306 436294 111374 436350
rect 111430 436294 111498 436350
rect 111554 436294 111622 436350
rect 111678 436294 129250 436350
rect 129306 436294 129374 436350
rect 129430 436294 129498 436350
rect 129554 436294 129622 436350
rect 129678 436294 147250 436350
rect 147306 436294 147374 436350
rect 147430 436294 147498 436350
rect 147554 436294 147622 436350
rect 147678 436294 165250 436350
rect 165306 436294 165374 436350
rect 165430 436294 165498 436350
rect 165554 436294 165622 436350
rect 165678 436294 183250 436350
rect 183306 436294 183374 436350
rect 183430 436294 183498 436350
rect 183554 436294 183622 436350
rect 183678 436294 201250 436350
rect 201306 436294 201374 436350
rect 201430 436294 201498 436350
rect 201554 436294 201622 436350
rect 201678 436294 204518 436350
rect 204574 436294 204642 436350
rect 204698 436294 235238 436350
rect 235294 436294 235362 436350
rect 235418 436294 265958 436350
rect 266014 436294 266082 436350
rect 266138 436294 296678 436350
rect 296734 436294 296802 436350
rect 296858 436294 327398 436350
rect 327454 436294 327522 436350
rect 327578 436294 358118 436350
rect 358174 436294 358242 436350
rect 358298 436294 388838 436350
rect 388894 436294 388962 436350
rect 389018 436294 419558 436350
rect 419614 436294 419682 436350
rect 419738 436294 450278 436350
rect 450334 436294 450402 436350
rect 450458 436294 480998 436350
rect 481054 436294 481122 436350
rect 481178 436294 507250 436350
rect 507306 436294 507374 436350
rect 507430 436294 507498 436350
rect 507554 436294 507622 436350
rect 507678 436294 525250 436350
rect 525306 436294 525374 436350
rect 525430 436294 525498 436350
rect 525554 436294 525622 436350
rect 525678 436294 543250 436350
rect 543306 436294 543374 436350
rect 543430 436294 543498 436350
rect 543554 436294 543622 436350
rect 543678 436294 561250 436350
rect 561306 436294 561374 436350
rect 561430 436294 561498 436350
rect 561554 436294 561622 436350
rect 561678 436294 579250 436350
rect 579306 436294 579374 436350
rect 579430 436294 579498 436350
rect 579554 436294 579622 436350
rect 579678 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 3250 436226
rect 3306 436170 3374 436226
rect 3430 436170 3498 436226
rect 3554 436170 3622 436226
rect 3678 436170 21250 436226
rect 21306 436170 21374 436226
rect 21430 436170 21498 436226
rect 21554 436170 21622 436226
rect 21678 436170 39250 436226
rect 39306 436170 39374 436226
rect 39430 436170 39498 436226
rect 39554 436170 39622 436226
rect 39678 436170 57250 436226
rect 57306 436170 57374 436226
rect 57430 436170 57498 436226
rect 57554 436170 57622 436226
rect 57678 436170 75250 436226
rect 75306 436170 75374 436226
rect 75430 436170 75498 436226
rect 75554 436170 75622 436226
rect 75678 436170 93250 436226
rect 93306 436170 93374 436226
rect 93430 436170 93498 436226
rect 93554 436170 93622 436226
rect 93678 436170 111250 436226
rect 111306 436170 111374 436226
rect 111430 436170 111498 436226
rect 111554 436170 111622 436226
rect 111678 436170 129250 436226
rect 129306 436170 129374 436226
rect 129430 436170 129498 436226
rect 129554 436170 129622 436226
rect 129678 436170 147250 436226
rect 147306 436170 147374 436226
rect 147430 436170 147498 436226
rect 147554 436170 147622 436226
rect 147678 436170 165250 436226
rect 165306 436170 165374 436226
rect 165430 436170 165498 436226
rect 165554 436170 165622 436226
rect 165678 436170 183250 436226
rect 183306 436170 183374 436226
rect 183430 436170 183498 436226
rect 183554 436170 183622 436226
rect 183678 436170 201250 436226
rect 201306 436170 201374 436226
rect 201430 436170 201498 436226
rect 201554 436170 201622 436226
rect 201678 436170 204518 436226
rect 204574 436170 204642 436226
rect 204698 436170 235238 436226
rect 235294 436170 235362 436226
rect 235418 436170 265958 436226
rect 266014 436170 266082 436226
rect 266138 436170 296678 436226
rect 296734 436170 296802 436226
rect 296858 436170 327398 436226
rect 327454 436170 327522 436226
rect 327578 436170 358118 436226
rect 358174 436170 358242 436226
rect 358298 436170 388838 436226
rect 388894 436170 388962 436226
rect 389018 436170 419558 436226
rect 419614 436170 419682 436226
rect 419738 436170 450278 436226
rect 450334 436170 450402 436226
rect 450458 436170 480998 436226
rect 481054 436170 481122 436226
rect 481178 436170 507250 436226
rect 507306 436170 507374 436226
rect 507430 436170 507498 436226
rect 507554 436170 507622 436226
rect 507678 436170 525250 436226
rect 525306 436170 525374 436226
rect 525430 436170 525498 436226
rect 525554 436170 525622 436226
rect 525678 436170 543250 436226
rect 543306 436170 543374 436226
rect 543430 436170 543498 436226
rect 543554 436170 543622 436226
rect 543678 436170 561250 436226
rect 561306 436170 561374 436226
rect 561430 436170 561498 436226
rect 561554 436170 561622 436226
rect 561678 436170 579250 436226
rect 579306 436170 579374 436226
rect 579430 436170 579498 436226
rect 579554 436170 579622 436226
rect 579678 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 3250 436102
rect 3306 436046 3374 436102
rect 3430 436046 3498 436102
rect 3554 436046 3622 436102
rect 3678 436046 21250 436102
rect 21306 436046 21374 436102
rect 21430 436046 21498 436102
rect 21554 436046 21622 436102
rect 21678 436046 39250 436102
rect 39306 436046 39374 436102
rect 39430 436046 39498 436102
rect 39554 436046 39622 436102
rect 39678 436046 57250 436102
rect 57306 436046 57374 436102
rect 57430 436046 57498 436102
rect 57554 436046 57622 436102
rect 57678 436046 75250 436102
rect 75306 436046 75374 436102
rect 75430 436046 75498 436102
rect 75554 436046 75622 436102
rect 75678 436046 93250 436102
rect 93306 436046 93374 436102
rect 93430 436046 93498 436102
rect 93554 436046 93622 436102
rect 93678 436046 111250 436102
rect 111306 436046 111374 436102
rect 111430 436046 111498 436102
rect 111554 436046 111622 436102
rect 111678 436046 129250 436102
rect 129306 436046 129374 436102
rect 129430 436046 129498 436102
rect 129554 436046 129622 436102
rect 129678 436046 147250 436102
rect 147306 436046 147374 436102
rect 147430 436046 147498 436102
rect 147554 436046 147622 436102
rect 147678 436046 165250 436102
rect 165306 436046 165374 436102
rect 165430 436046 165498 436102
rect 165554 436046 165622 436102
rect 165678 436046 183250 436102
rect 183306 436046 183374 436102
rect 183430 436046 183498 436102
rect 183554 436046 183622 436102
rect 183678 436046 201250 436102
rect 201306 436046 201374 436102
rect 201430 436046 201498 436102
rect 201554 436046 201622 436102
rect 201678 436046 204518 436102
rect 204574 436046 204642 436102
rect 204698 436046 235238 436102
rect 235294 436046 235362 436102
rect 235418 436046 265958 436102
rect 266014 436046 266082 436102
rect 266138 436046 296678 436102
rect 296734 436046 296802 436102
rect 296858 436046 327398 436102
rect 327454 436046 327522 436102
rect 327578 436046 358118 436102
rect 358174 436046 358242 436102
rect 358298 436046 388838 436102
rect 388894 436046 388962 436102
rect 389018 436046 419558 436102
rect 419614 436046 419682 436102
rect 419738 436046 450278 436102
rect 450334 436046 450402 436102
rect 450458 436046 480998 436102
rect 481054 436046 481122 436102
rect 481178 436046 507250 436102
rect 507306 436046 507374 436102
rect 507430 436046 507498 436102
rect 507554 436046 507622 436102
rect 507678 436046 525250 436102
rect 525306 436046 525374 436102
rect 525430 436046 525498 436102
rect 525554 436046 525622 436102
rect 525678 436046 543250 436102
rect 543306 436046 543374 436102
rect 543430 436046 543498 436102
rect 543554 436046 543622 436102
rect 543678 436046 561250 436102
rect 561306 436046 561374 436102
rect 561430 436046 561498 436102
rect 561554 436046 561622 436102
rect 561678 436046 579250 436102
rect 579306 436046 579374 436102
rect 579430 436046 579498 436102
rect 579554 436046 579622 436102
rect 579678 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 3250 435978
rect 3306 435922 3374 435978
rect 3430 435922 3498 435978
rect 3554 435922 3622 435978
rect 3678 435922 21250 435978
rect 21306 435922 21374 435978
rect 21430 435922 21498 435978
rect 21554 435922 21622 435978
rect 21678 435922 39250 435978
rect 39306 435922 39374 435978
rect 39430 435922 39498 435978
rect 39554 435922 39622 435978
rect 39678 435922 57250 435978
rect 57306 435922 57374 435978
rect 57430 435922 57498 435978
rect 57554 435922 57622 435978
rect 57678 435922 75250 435978
rect 75306 435922 75374 435978
rect 75430 435922 75498 435978
rect 75554 435922 75622 435978
rect 75678 435922 93250 435978
rect 93306 435922 93374 435978
rect 93430 435922 93498 435978
rect 93554 435922 93622 435978
rect 93678 435922 111250 435978
rect 111306 435922 111374 435978
rect 111430 435922 111498 435978
rect 111554 435922 111622 435978
rect 111678 435922 129250 435978
rect 129306 435922 129374 435978
rect 129430 435922 129498 435978
rect 129554 435922 129622 435978
rect 129678 435922 147250 435978
rect 147306 435922 147374 435978
rect 147430 435922 147498 435978
rect 147554 435922 147622 435978
rect 147678 435922 165250 435978
rect 165306 435922 165374 435978
rect 165430 435922 165498 435978
rect 165554 435922 165622 435978
rect 165678 435922 183250 435978
rect 183306 435922 183374 435978
rect 183430 435922 183498 435978
rect 183554 435922 183622 435978
rect 183678 435922 201250 435978
rect 201306 435922 201374 435978
rect 201430 435922 201498 435978
rect 201554 435922 201622 435978
rect 201678 435922 204518 435978
rect 204574 435922 204642 435978
rect 204698 435922 235238 435978
rect 235294 435922 235362 435978
rect 235418 435922 265958 435978
rect 266014 435922 266082 435978
rect 266138 435922 296678 435978
rect 296734 435922 296802 435978
rect 296858 435922 327398 435978
rect 327454 435922 327522 435978
rect 327578 435922 358118 435978
rect 358174 435922 358242 435978
rect 358298 435922 388838 435978
rect 388894 435922 388962 435978
rect 389018 435922 419558 435978
rect 419614 435922 419682 435978
rect 419738 435922 450278 435978
rect 450334 435922 450402 435978
rect 450458 435922 480998 435978
rect 481054 435922 481122 435978
rect 481178 435922 507250 435978
rect 507306 435922 507374 435978
rect 507430 435922 507498 435978
rect 507554 435922 507622 435978
rect 507678 435922 525250 435978
rect 525306 435922 525374 435978
rect 525430 435922 525498 435978
rect 525554 435922 525622 435978
rect 525678 435922 543250 435978
rect 543306 435922 543374 435978
rect 543430 435922 543498 435978
rect 543554 435922 543622 435978
rect 543678 435922 561250 435978
rect 561306 435922 561374 435978
rect 561430 435922 561498 435978
rect 561554 435922 561622 435978
rect 561678 435922 579250 435978
rect 579306 435922 579374 435978
rect 579430 435922 579498 435978
rect 579554 435922 579622 435978
rect 579678 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 6970 424350
rect 7026 424294 7094 424350
rect 7150 424294 7218 424350
rect 7274 424294 7342 424350
rect 7398 424294 24970 424350
rect 25026 424294 25094 424350
rect 25150 424294 25218 424350
rect 25274 424294 25342 424350
rect 25398 424294 42970 424350
rect 43026 424294 43094 424350
rect 43150 424294 43218 424350
rect 43274 424294 43342 424350
rect 43398 424294 60970 424350
rect 61026 424294 61094 424350
rect 61150 424294 61218 424350
rect 61274 424294 61342 424350
rect 61398 424294 78970 424350
rect 79026 424294 79094 424350
rect 79150 424294 79218 424350
rect 79274 424294 79342 424350
rect 79398 424294 96970 424350
rect 97026 424294 97094 424350
rect 97150 424294 97218 424350
rect 97274 424294 97342 424350
rect 97398 424294 114970 424350
rect 115026 424294 115094 424350
rect 115150 424294 115218 424350
rect 115274 424294 115342 424350
rect 115398 424294 132970 424350
rect 133026 424294 133094 424350
rect 133150 424294 133218 424350
rect 133274 424294 133342 424350
rect 133398 424294 150970 424350
rect 151026 424294 151094 424350
rect 151150 424294 151218 424350
rect 151274 424294 151342 424350
rect 151398 424294 168970 424350
rect 169026 424294 169094 424350
rect 169150 424294 169218 424350
rect 169274 424294 169342 424350
rect 169398 424294 186970 424350
rect 187026 424294 187094 424350
rect 187150 424294 187218 424350
rect 187274 424294 187342 424350
rect 187398 424294 219878 424350
rect 219934 424294 220002 424350
rect 220058 424294 250598 424350
rect 250654 424294 250722 424350
rect 250778 424294 281318 424350
rect 281374 424294 281442 424350
rect 281498 424294 312038 424350
rect 312094 424294 312162 424350
rect 312218 424294 342758 424350
rect 342814 424294 342882 424350
rect 342938 424294 373478 424350
rect 373534 424294 373602 424350
rect 373658 424294 404198 424350
rect 404254 424294 404322 424350
rect 404378 424294 434918 424350
rect 434974 424294 435042 424350
rect 435098 424294 465638 424350
rect 465694 424294 465762 424350
rect 465818 424294 496358 424350
rect 496414 424294 496482 424350
rect 496538 424294 510970 424350
rect 511026 424294 511094 424350
rect 511150 424294 511218 424350
rect 511274 424294 511342 424350
rect 511398 424294 528970 424350
rect 529026 424294 529094 424350
rect 529150 424294 529218 424350
rect 529274 424294 529342 424350
rect 529398 424294 546970 424350
rect 547026 424294 547094 424350
rect 547150 424294 547218 424350
rect 547274 424294 547342 424350
rect 547398 424294 564970 424350
rect 565026 424294 565094 424350
rect 565150 424294 565218 424350
rect 565274 424294 565342 424350
rect 565398 424294 582970 424350
rect 583026 424294 583094 424350
rect 583150 424294 583218 424350
rect 583274 424294 583342 424350
rect 583398 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 6970 424226
rect 7026 424170 7094 424226
rect 7150 424170 7218 424226
rect 7274 424170 7342 424226
rect 7398 424170 24970 424226
rect 25026 424170 25094 424226
rect 25150 424170 25218 424226
rect 25274 424170 25342 424226
rect 25398 424170 42970 424226
rect 43026 424170 43094 424226
rect 43150 424170 43218 424226
rect 43274 424170 43342 424226
rect 43398 424170 60970 424226
rect 61026 424170 61094 424226
rect 61150 424170 61218 424226
rect 61274 424170 61342 424226
rect 61398 424170 78970 424226
rect 79026 424170 79094 424226
rect 79150 424170 79218 424226
rect 79274 424170 79342 424226
rect 79398 424170 96970 424226
rect 97026 424170 97094 424226
rect 97150 424170 97218 424226
rect 97274 424170 97342 424226
rect 97398 424170 114970 424226
rect 115026 424170 115094 424226
rect 115150 424170 115218 424226
rect 115274 424170 115342 424226
rect 115398 424170 132970 424226
rect 133026 424170 133094 424226
rect 133150 424170 133218 424226
rect 133274 424170 133342 424226
rect 133398 424170 150970 424226
rect 151026 424170 151094 424226
rect 151150 424170 151218 424226
rect 151274 424170 151342 424226
rect 151398 424170 168970 424226
rect 169026 424170 169094 424226
rect 169150 424170 169218 424226
rect 169274 424170 169342 424226
rect 169398 424170 186970 424226
rect 187026 424170 187094 424226
rect 187150 424170 187218 424226
rect 187274 424170 187342 424226
rect 187398 424170 219878 424226
rect 219934 424170 220002 424226
rect 220058 424170 250598 424226
rect 250654 424170 250722 424226
rect 250778 424170 281318 424226
rect 281374 424170 281442 424226
rect 281498 424170 312038 424226
rect 312094 424170 312162 424226
rect 312218 424170 342758 424226
rect 342814 424170 342882 424226
rect 342938 424170 373478 424226
rect 373534 424170 373602 424226
rect 373658 424170 404198 424226
rect 404254 424170 404322 424226
rect 404378 424170 434918 424226
rect 434974 424170 435042 424226
rect 435098 424170 465638 424226
rect 465694 424170 465762 424226
rect 465818 424170 496358 424226
rect 496414 424170 496482 424226
rect 496538 424170 510970 424226
rect 511026 424170 511094 424226
rect 511150 424170 511218 424226
rect 511274 424170 511342 424226
rect 511398 424170 528970 424226
rect 529026 424170 529094 424226
rect 529150 424170 529218 424226
rect 529274 424170 529342 424226
rect 529398 424170 546970 424226
rect 547026 424170 547094 424226
rect 547150 424170 547218 424226
rect 547274 424170 547342 424226
rect 547398 424170 564970 424226
rect 565026 424170 565094 424226
rect 565150 424170 565218 424226
rect 565274 424170 565342 424226
rect 565398 424170 582970 424226
rect 583026 424170 583094 424226
rect 583150 424170 583218 424226
rect 583274 424170 583342 424226
rect 583398 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 6970 424102
rect 7026 424046 7094 424102
rect 7150 424046 7218 424102
rect 7274 424046 7342 424102
rect 7398 424046 24970 424102
rect 25026 424046 25094 424102
rect 25150 424046 25218 424102
rect 25274 424046 25342 424102
rect 25398 424046 42970 424102
rect 43026 424046 43094 424102
rect 43150 424046 43218 424102
rect 43274 424046 43342 424102
rect 43398 424046 60970 424102
rect 61026 424046 61094 424102
rect 61150 424046 61218 424102
rect 61274 424046 61342 424102
rect 61398 424046 78970 424102
rect 79026 424046 79094 424102
rect 79150 424046 79218 424102
rect 79274 424046 79342 424102
rect 79398 424046 96970 424102
rect 97026 424046 97094 424102
rect 97150 424046 97218 424102
rect 97274 424046 97342 424102
rect 97398 424046 114970 424102
rect 115026 424046 115094 424102
rect 115150 424046 115218 424102
rect 115274 424046 115342 424102
rect 115398 424046 132970 424102
rect 133026 424046 133094 424102
rect 133150 424046 133218 424102
rect 133274 424046 133342 424102
rect 133398 424046 150970 424102
rect 151026 424046 151094 424102
rect 151150 424046 151218 424102
rect 151274 424046 151342 424102
rect 151398 424046 168970 424102
rect 169026 424046 169094 424102
rect 169150 424046 169218 424102
rect 169274 424046 169342 424102
rect 169398 424046 186970 424102
rect 187026 424046 187094 424102
rect 187150 424046 187218 424102
rect 187274 424046 187342 424102
rect 187398 424046 219878 424102
rect 219934 424046 220002 424102
rect 220058 424046 250598 424102
rect 250654 424046 250722 424102
rect 250778 424046 281318 424102
rect 281374 424046 281442 424102
rect 281498 424046 312038 424102
rect 312094 424046 312162 424102
rect 312218 424046 342758 424102
rect 342814 424046 342882 424102
rect 342938 424046 373478 424102
rect 373534 424046 373602 424102
rect 373658 424046 404198 424102
rect 404254 424046 404322 424102
rect 404378 424046 434918 424102
rect 434974 424046 435042 424102
rect 435098 424046 465638 424102
rect 465694 424046 465762 424102
rect 465818 424046 496358 424102
rect 496414 424046 496482 424102
rect 496538 424046 510970 424102
rect 511026 424046 511094 424102
rect 511150 424046 511218 424102
rect 511274 424046 511342 424102
rect 511398 424046 528970 424102
rect 529026 424046 529094 424102
rect 529150 424046 529218 424102
rect 529274 424046 529342 424102
rect 529398 424046 546970 424102
rect 547026 424046 547094 424102
rect 547150 424046 547218 424102
rect 547274 424046 547342 424102
rect 547398 424046 564970 424102
rect 565026 424046 565094 424102
rect 565150 424046 565218 424102
rect 565274 424046 565342 424102
rect 565398 424046 582970 424102
rect 583026 424046 583094 424102
rect 583150 424046 583218 424102
rect 583274 424046 583342 424102
rect 583398 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 6970 423978
rect 7026 423922 7094 423978
rect 7150 423922 7218 423978
rect 7274 423922 7342 423978
rect 7398 423922 24970 423978
rect 25026 423922 25094 423978
rect 25150 423922 25218 423978
rect 25274 423922 25342 423978
rect 25398 423922 42970 423978
rect 43026 423922 43094 423978
rect 43150 423922 43218 423978
rect 43274 423922 43342 423978
rect 43398 423922 60970 423978
rect 61026 423922 61094 423978
rect 61150 423922 61218 423978
rect 61274 423922 61342 423978
rect 61398 423922 78970 423978
rect 79026 423922 79094 423978
rect 79150 423922 79218 423978
rect 79274 423922 79342 423978
rect 79398 423922 96970 423978
rect 97026 423922 97094 423978
rect 97150 423922 97218 423978
rect 97274 423922 97342 423978
rect 97398 423922 114970 423978
rect 115026 423922 115094 423978
rect 115150 423922 115218 423978
rect 115274 423922 115342 423978
rect 115398 423922 132970 423978
rect 133026 423922 133094 423978
rect 133150 423922 133218 423978
rect 133274 423922 133342 423978
rect 133398 423922 150970 423978
rect 151026 423922 151094 423978
rect 151150 423922 151218 423978
rect 151274 423922 151342 423978
rect 151398 423922 168970 423978
rect 169026 423922 169094 423978
rect 169150 423922 169218 423978
rect 169274 423922 169342 423978
rect 169398 423922 186970 423978
rect 187026 423922 187094 423978
rect 187150 423922 187218 423978
rect 187274 423922 187342 423978
rect 187398 423922 219878 423978
rect 219934 423922 220002 423978
rect 220058 423922 250598 423978
rect 250654 423922 250722 423978
rect 250778 423922 281318 423978
rect 281374 423922 281442 423978
rect 281498 423922 312038 423978
rect 312094 423922 312162 423978
rect 312218 423922 342758 423978
rect 342814 423922 342882 423978
rect 342938 423922 373478 423978
rect 373534 423922 373602 423978
rect 373658 423922 404198 423978
rect 404254 423922 404322 423978
rect 404378 423922 434918 423978
rect 434974 423922 435042 423978
rect 435098 423922 465638 423978
rect 465694 423922 465762 423978
rect 465818 423922 496358 423978
rect 496414 423922 496482 423978
rect 496538 423922 510970 423978
rect 511026 423922 511094 423978
rect 511150 423922 511218 423978
rect 511274 423922 511342 423978
rect 511398 423922 528970 423978
rect 529026 423922 529094 423978
rect 529150 423922 529218 423978
rect 529274 423922 529342 423978
rect 529398 423922 546970 423978
rect 547026 423922 547094 423978
rect 547150 423922 547218 423978
rect 547274 423922 547342 423978
rect 547398 423922 564970 423978
rect 565026 423922 565094 423978
rect 565150 423922 565218 423978
rect 565274 423922 565342 423978
rect 565398 423922 582970 423978
rect 583026 423922 583094 423978
rect 583150 423922 583218 423978
rect 583274 423922 583342 423978
rect 583398 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 3250 418350
rect 3306 418294 3374 418350
rect 3430 418294 3498 418350
rect 3554 418294 3622 418350
rect 3678 418294 21250 418350
rect 21306 418294 21374 418350
rect 21430 418294 21498 418350
rect 21554 418294 21622 418350
rect 21678 418294 39250 418350
rect 39306 418294 39374 418350
rect 39430 418294 39498 418350
rect 39554 418294 39622 418350
rect 39678 418294 57250 418350
rect 57306 418294 57374 418350
rect 57430 418294 57498 418350
rect 57554 418294 57622 418350
rect 57678 418294 75250 418350
rect 75306 418294 75374 418350
rect 75430 418294 75498 418350
rect 75554 418294 75622 418350
rect 75678 418294 93250 418350
rect 93306 418294 93374 418350
rect 93430 418294 93498 418350
rect 93554 418294 93622 418350
rect 93678 418294 111250 418350
rect 111306 418294 111374 418350
rect 111430 418294 111498 418350
rect 111554 418294 111622 418350
rect 111678 418294 129250 418350
rect 129306 418294 129374 418350
rect 129430 418294 129498 418350
rect 129554 418294 129622 418350
rect 129678 418294 147250 418350
rect 147306 418294 147374 418350
rect 147430 418294 147498 418350
rect 147554 418294 147622 418350
rect 147678 418294 165250 418350
rect 165306 418294 165374 418350
rect 165430 418294 165498 418350
rect 165554 418294 165622 418350
rect 165678 418294 183250 418350
rect 183306 418294 183374 418350
rect 183430 418294 183498 418350
rect 183554 418294 183622 418350
rect 183678 418294 201250 418350
rect 201306 418294 201374 418350
rect 201430 418294 201498 418350
rect 201554 418294 201622 418350
rect 201678 418294 204518 418350
rect 204574 418294 204642 418350
rect 204698 418294 235238 418350
rect 235294 418294 235362 418350
rect 235418 418294 265958 418350
rect 266014 418294 266082 418350
rect 266138 418294 296678 418350
rect 296734 418294 296802 418350
rect 296858 418294 327398 418350
rect 327454 418294 327522 418350
rect 327578 418294 358118 418350
rect 358174 418294 358242 418350
rect 358298 418294 388838 418350
rect 388894 418294 388962 418350
rect 389018 418294 419558 418350
rect 419614 418294 419682 418350
rect 419738 418294 450278 418350
rect 450334 418294 450402 418350
rect 450458 418294 480998 418350
rect 481054 418294 481122 418350
rect 481178 418294 507250 418350
rect 507306 418294 507374 418350
rect 507430 418294 507498 418350
rect 507554 418294 507622 418350
rect 507678 418294 525250 418350
rect 525306 418294 525374 418350
rect 525430 418294 525498 418350
rect 525554 418294 525622 418350
rect 525678 418294 543250 418350
rect 543306 418294 543374 418350
rect 543430 418294 543498 418350
rect 543554 418294 543622 418350
rect 543678 418294 561250 418350
rect 561306 418294 561374 418350
rect 561430 418294 561498 418350
rect 561554 418294 561622 418350
rect 561678 418294 579250 418350
rect 579306 418294 579374 418350
rect 579430 418294 579498 418350
rect 579554 418294 579622 418350
rect 579678 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 3250 418226
rect 3306 418170 3374 418226
rect 3430 418170 3498 418226
rect 3554 418170 3622 418226
rect 3678 418170 21250 418226
rect 21306 418170 21374 418226
rect 21430 418170 21498 418226
rect 21554 418170 21622 418226
rect 21678 418170 39250 418226
rect 39306 418170 39374 418226
rect 39430 418170 39498 418226
rect 39554 418170 39622 418226
rect 39678 418170 57250 418226
rect 57306 418170 57374 418226
rect 57430 418170 57498 418226
rect 57554 418170 57622 418226
rect 57678 418170 75250 418226
rect 75306 418170 75374 418226
rect 75430 418170 75498 418226
rect 75554 418170 75622 418226
rect 75678 418170 93250 418226
rect 93306 418170 93374 418226
rect 93430 418170 93498 418226
rect 93554 418170 93622 418226
rect 93678 418170 111250 418226
rect 111306 418170 111374 418226
rect 111430 418170 111498 418226
rect 111554 418170 111622 418226
rect 111678 418170 129250 418226
rect 129306 418170 129374 418226
rect 129430 418170 129498 418226
rect 129554 418170 129622 418226
rect 129678 418170 147250 418226
rect 147306 418170 147374 418226
rect 147430 418170 147498 418226
rect 147554 418170 147622 418226
rect 147678 418170 165250 418226
rect 165306 418170 165374 418226
rect 165430 418170 165498 418226
rect 165554 418170 165622 418226
rect 165678 418170 183250 418226
rect 183306 418170 183374 418226
rect 183430 418170 183498 418226
rect 183554 418170 183622 418226
rect 183678 418170 201250 418226
rect 201306 418170 201374 418226
rect 201430 418170 201498 418226
rect 201554 418170 201622 418226
rect 201678 418170 204518 418226
rect 204574 418170 204642 418226
rect 204698 418170 235238 418226
rect 235294 418170 235362 418226
rect 235418 418170 265958 418226
rect 266014 418170 266082 418226
rect 266138 418170 296678 418226
rect 296734 418170 296802 418226
rect 296858 418170 327398 418226
rect 327454 418170 327522 418226
rect 327578 418170 358118 418226
rect 358174 418170 358242 418226
rect 358298 418170 388838 418226
rect 388894 418170 388962 418226
rect 389018 418170 419558 418226
rect 419614 418170 419682 418226
rect 419738 418170 450278 418226
rect 450334 418170 450402 418226
rect 450458 418170 480998 418226
rect 481054 418170 481122 418226
rect 481178 418170 507250 418226
rect 507306 418170 507374 418226
rect 507430 418170 507498 418226
rect 507554 418170 507622 418226
rect 507678 418170 525250 418226
rect 525306 418170 525374 418226
rect 525430 418170 525498 418226
rect 525554 418170 525622 418226
rect 525678 418170 543250 418226
rect 543306 418170 543374 418226
rect 543430 418170 543498 418226
rect 543554 418170 543622 418226
rect 543678 418170 561250 418226
rect 561306 418170 561374 418226
rect 561430 418170 561498 418226
rect 561554 418170 561622 418226
rect 561678 418170 579250 418226
rect 579306 418170 579374 418226
rect 579430 418170 579498 418226
rect 579554 418170 579622 418226
rect 579678 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 3250 418102
rect 3306 418046 3374 418102
rect 3430 418046 3498 418102
rect 3554 418046 3622 418102
rect 3678 418046 21250 418102
rect 21306 418046 21374 418102
rect 21430 418046 21498 418102
rect 21554 418046 21622 418102
rect 21678 418046 39250 418102
rect 39306 418046 39374 418102
rect 39430 418046 39498 418102
rect 39554 418046 39622 418102
rect 39678 418046 57250 418102
rect 57306 418046 57374 418102
rect 57430 418046 57498 418102
rect 57554 418046 57622 418102
rect 57678 418046 75250 418102
rect 75306 418046 75374 418102
rect 75430 418046 75498 418102
rect 75554 418046 75622 418102
rect 75678 418046 93250 418102
rect 93306 418046 93374 418102
rect 93430 418046 93498 418102
rect 93554 418046 93622 418102
rect 93678 418046 111250 418102
rect 111306 418046 111374 418102
rect 111430 418046 111498 418102
rect 111554 418046 111622 418102
rect 111678 418046 129250 418102
rect 129306 418046 129374 418102
rect 129430 418046 129498 418102
rect 129554 418046 129622 418102
rect 129678 418046 147250 418102
rect 147306 418046 147374 418102
rect 147430 418046 147498 418102
rect 147554 418046 147622 418102
rect 147678 418046 165250 418102
rect 165306 418046 165374 418102
rect 165430 418046 165498 418102
rect 165554 418046 165622 418102
rect 165678 418046 183250 418102
rect 183306 418046 183374 418102
rect 183430 418046 183498 418102
rect 183554 418046 183622 418102
rect 183678 418046 201250 418102
rect 201306 418046 201374 418102
rect 201430 418046 201498 418102
rect 201554 418046 201622 418102
rect 201678 418046 204518 418102
rect 204574 418046 204642 418102
rect 204698 418046 235238 418102
rect 235294 418046 235362 418102
rect 235418 418046 265958 418102
rect 266014 418046 266082 418102
rect 266138 418046 296678 418102
rect 296734 418046 296802 418102
rect 296858 418046 327398 418102
rect 327454 418046 327522 418102
rect 327578 418046 358118 418102
rect 358174 418046 358242 418102
rect 358298 418046 388838 418102
rect 388894 418046 388962 418102
rect 389018 418046 419558 418102
rect 419614 418046 419682 418102
rect 419738 418046 450278 418102
rect 450334 418046 450402 418102
rect 450458 418046 480998 418102
rect 481054 418046 481122 418102
rect 481178 418046 507250 418102
rect 507306 418046 507374 418102
rect 507430 418046 507498 418102
rect 507554 418046 507622 418102
rect 507678 418046 525250 418102
rect 525306 418046 525374 418102
rect 525430 418046 525498 418102
rect 525554 418046 525622 418102
rect 525678 418046 543250 418102
rect 543306 418046 543374 418102
rect 543430 418046 543498 418102
rect 543554 418046 543622 418102
rect 543678 418046 561250 418102
rect 561306 418046 561374 418102
rect 561430 418046 561498 418102
rect 561554 418046 561622 418102
rect 561678 418046 579250 418102
rect 579306 418046 579374 418102
rect 579430 418046 579498 418102
rect 579554 418046 579622 418102
rect 579678 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 3250 417978
rect 3306 417922 3374 417978
rect 3430 417922 3498 417978
rect 3554 417922 3622 417978
rect 3678 417922 21250 417978
rect 21306 417922 21374 417978
rect 21430 417922 21498 417978
rect 21554 417922 21622 417978
rect 21678 417922 39250 417978
rect 39306 417922 39374 417978
rect 39430 417922 39498 417978
rect 39554 417922 39622 417978
rect 39678 417922 57250 417978
rect 57306 417922 57374 417978
rect 57430 417922 57498 417978
rect 57554 417922 57622 417978
rect 57678 417922 75250 417978
rect 75306 417922 75374 417978
rect 75430 417922 75498 417978
rect 75554 417922 75622 417978
rect 75678 417922 93250 417978
rect 93306 417922 93374 417978
rect 93430 417922 93498 417978
rect 93554 417922 93622 417978
rect 93678 417922 111250 417978
rect 111306 417922 111374 417978
rect 111430 417922 111498 417978
rect 111554 417922 111622 417978
rect 111678 417922 129250 417978
rect 129306 417922 129374 417978
rect 129430 417922 129498 417978
rect 129554 417922 129622 417978
rect 129678 417922 147250 417978
rect 147306 417922 147374 417978
rect 147430 417922 147498 417978
rect 147554 417922 147622 417978
rect 147678 417922 165250 417978
rect 165306 417922 165374 417978
rect 165430 417922 165498 417978
rect 165554 417922 165622 417978
rect 165678 417922 183250 417978
rect 183306 417922 183374 417978
rect 183430 417922 183498 417978
rect 183554 417922 183622 417978
rect 183678 417922 201250 417978
rect 201306 417922 201374 417978
rect 201430 417922 201498 417978
rect 201554 417922 201622 417978
rect 201678 417922 204518 417978
rect 204574 417922 204642 417978
rect 204698 417922 235238 417978
rect 235294 417922 235362 417978
rect 235418 417922 265958 417978
rect 266014 417922 266082 417978
rect 266138 417922 296678 417978
rect 296734 417922 296802 417978
rect 296858 417922 327398 417978
rect 327454 417922 327522 417978
rect 327578 417922 358118 417978
rect 358174 417922 358242 417978
rect 358298 417922 388838 417978
rect 388894 417922 388962 417978
rect 389018 417922 419558 417978
rect 419614 417922 419682 417978
rect 419738 417922 450278 417978
rect 450334 417922 450402 417978
rect 450458 417922 480998 417978
rect 481054 417922 481122 417978
rect 481178 417922 507250 417978
rect 507306 417922 507374 417978
rect 507430 417922 507498 417978
rect 507554 417922 507622 417978
rect 507678 417922 525250 417978
rect 525306 417922 525374 417978
rect 525430 417922 525498 417978
rect 525554 417922 525622 417978
rect 525678 417922 543250 417978
rect 543306 417922 543374 417978
rect 543430 417922 543498 417978
rect 543554 417922 543622 417978
rect 543678 417922 561250 417978
rect 561306 417922 561374 417978
rect 561430 417922 561498 417978
rect 561554 417922 561622 417978
rect 561678 417922 579250 417978
rect 579306 417922 579374 417978
rect 579430 417922 579498 417978
rect 579554 417922 579622 417978
rect 579678 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 6970 406350
rect 7026 406294 7094 406350
rect 7150 406294 7218 406350
rect 7274 406294 7342 406350
rect 7398 406294 24970 406350
rect 25026 406294 25094 406350
rect 25150 406294 25218 406350
rect 25274 406294 25342 406350
rect 25398 406294 42970 406350
rect 43026 406294 43094 406350
rect 43150 406294 43218 406350
rect 43274 406294 43342 406350
rect 43398 406294 60970 406350
rect 61026 406294 61094 406350
rect 61150 406294 61218 406350
rect 61274 406294 61342 406350
rect 61398 406294 78970 406350
rect 79026 406294 79094 406350
rect 79150 406294 79218 406350
rect 79274 406294 79342 406350
rect 79398 406294 96970 406350
rect 97026 406294 97094 406350
rect 97150 406294 97218 406350
rect 97274 406294 97342 406350
rect 97398 406294 114970 406350
rect 115026 406294 115094 406350
rect 115150 406294 115218 406350
rect 115274 406294 115342 406350
rect 115398 406294 132970 406350
rect 133026 406294 133094 406350
rect 133150 406294 133218 406350
rect 133274 406294 133342 406350
rect 133398 406294 150970 406350
rect 151026 406294 151094 406350
rect 151150 406294 151218 406350
rect 151274 406294 151342 406350
rect 151398 406294 168970 406350
rect 169026 406294 169094 406350
rect 169150 406294 169218 406350
rect 169274 406294 169342 406350
rect 169398 406294 186970 406350
rect 187026 406294 187094 406350
rect 187150 406294 187218 406350
rect 187274 406294 187342 406350
rect 187398 406294 219878 406350
rect 219934 406294 220002 406350
rect 220058 406294 250598 406350
rect 250654 406294 250722 406350
rect 250778 406294 281318 406350
rect 281374 406294 281442 406350
rect 281498 406294 312038 406350
rect 312094 406294 312162 406350
rect 312218 406294 342758 406350
rect 342814 406294 342882 406350
rect 342938 406294 373478 406350
rect 373534 406294 373602 406350
rect 373658 406294 404198 406350
rect 404254 406294 404322 406350
rect 404378 406294 434918 406350
rect 434974 406294 435042 406350
rect 435098 406294 465638 406350
rect 465694 406294 465762 406350
rect 465818 406294 496358 406350
rect 496414 406294 496482 406350
rect 496538 406294 510970 406350
rect 511026 406294 511094 406350
rect 511150 406294 511218 406350
rect 511274 406294 511342 406350
rect 511398 406294 528970 406350
rect 529026 406294 529094 406350
rect 529150 406294 529218 406350
rect 529274 406294 529342 406350
rect 529398 406294 546970 406350
rect 547026 406294 547094 406350
rect 547150 406294 547218 406350
rect 547274 406294 547342 406350
rect 547398 406294 564970 406350
rect 565026 406294 565094 406350
rect 565150 406294 565218 406350
rect 565274 406294 565342 406350
rect 565398 406294 582970 406350
rect 583026 406294 583094 406350
rect 583150 406294 583218 406350
rect 583274 406294 583342 406350
rect 583398 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 6970 406226
rect 7026 406170 7094 406226
rect 7150 406170 7218 406226
rect 7274 406170 7342 406226
rect 7398 406170 24970 406226
rect 25026 406170 25094 406226
rect 25150 406170 25218 406226
rect 25274 406170 25342 406226
rect 25398 406170 42970 406226
rect 43026 406170 43094 406226
rect 43150 406170 43218 406226
rect 43274 406170 43342 406226
rect 43398 406170 60970 406226
rect 61026 406170 61094 406226
rect 61150 406170 61218 406226
rect 61274 406170 61342 406226
rect 61398 406170 78970 406226
rect 79026 406170 79094 406226
rect 79150 406170 79218 406226
rect 79274 406170 79342 406226
rect 79398 406170 96970 406226
rect 97026 406170 97094 406226
rect 97150 406170 97218 406226
rect 97274 406170 97342 406226
rect 97398 406170 114970 406226
rect 115026 406170 115094 406226
rect 115150 406170 115218 406226
rect 115274 406170 115342 406226
rect 115398 406170 132970 406226
rect 133026 406170 133094 406226
rect 133150 406170 133218 406226
rect 133274 406170 133342 406226
rect 133398 406170 150970 406226
rect 151026 406170 151094 406226
rect 151150 406170 151218 406226
rect 151274 406170 151342 406226
rect 151398 406170 168970 406226
rect 169026 406170 169094 406226
rect 169150 406170 169218 406226
rect 169274 406170 169342 406226
rect 169398 406170 186970 406226
rect 187026 406170 187094 406226
rect 187150 406170 187218 406226
rect 187274 406170 187342 406226
rect 187398 406170 219878 406226
rect 219934 406170 220002 406226
rect 220058 406170 250598 406226
rect 250654 406170 250722 406226
rect 250778 406170 281318 406226
rect 281374 406170 281442 406226
rect 281498 406170 312038 406226
rect 312094 406170 312162 406226
rect 312218 406170 342758 406226
rect 342814 406170 342882 406226
rect 342938 406170 373478 406226
rect 373534 406170 373602 406226
rect 373658 406170 404198 406226
rect 404254 406170 404322 406226
rect 404378 406170 434918 406226
rect 434974 406170 435042 406226
rect 435098 406170 465638 406226
rect 465694 406170 465762 406226
rect 465818 406170 496358 406226
rect 496414 406170 496482 406226
rect 496538 406170 510970 406226
rect 511026 406170 511094 406226
rect 511150 406170 511218 406226
rect 511274 406170 511342 406226
rect 511398 406170 528970 406226
rect 529026 406170 529094 406226
rect 529150 406170 529218 406226
rect 529274 406170 529342 406226
rect 529398 406170 546970 406226
rect 547026 406170 547094 406226
rect 547150 406170 547218 406226
rect 547274 406170 547342 406226
rect 547398 406170 564970 406226
rect 565026 406170 565094 406226
rect 565150 406170 565218 406226
rect 565274 406170 565342 406226
rect 565398 406170 582970 406226
rect 583026 406170 583094 406226
rect 583150 406170 583218 406226
rect 583274 406170 583342 406226
rect 583398 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 6970 406102
rect 7026 406046 7094 406102
rect 7150 406046 7218 406102
rect 7274 406046 7342 406102
rect 7398 406046 24970 406102
rect 25026 406046 25094 406102
rect 25150 406046 25218 406102
rect 25274 406046 25342 406102
rect 25398 406046 42970 406102
rect 43026 406046 43094 406102
rect 43150 406046 43218 406102
rect 43274 406046 43342 406102
rect 43398 406046 60970 406102
rect 61026 406046 61094 406102
rect 61150 406046 61218 406102
rect 61274 406046 61342 406102
rect 61398 406046 78970 406102
rect 79026 406046 79094 406102
rect 79150 406046 79218 406102
rect 79274 406046 79342 406102
rect 79398 406046 96970 406102
rect 97026 406046 97094 406102
rect 97150 406046 97218 406102
rect 97274 406046 97342 406102
rect 97398 406046 114970 406102
rect 115026 406046 115094 406102
rect 115150 406046 115218 406102
rect 115274 406046 115342 406102
rect 115398 406046 132970 406102
rect 133026 406046 133094 406102
rect 133150 406046 133218 406102
rect 133274 406046 133342 406102
rect 133398 406046 150970 406102
rect 151026 406046 151094 406102
rect 151150 406046 151218 406102
rect 151274 406046 151342 406102
rect 151398 406046 168970 406102
rect 169026 406046 169094 406102
rect 169150 406046 169218 406102
rect 169274 406046 169342 406102
rect 169398 406046 186970 406102
rect 187026 406046 187094 406102
rect 187150 406046 187218 406102
rect 187274 406046 187342 406102
rect 187398 406046 219878 406102
rect 219934 406046 220002 406102
rect 220058 406046 250598 406102
rect 250654 406046 250722 406102
rect 250778 406046 281318 406102
rect 281374 406046 281442 406102
rect 281498 406046 312038 406102
rect 312094 406046 312162 406102
rect 312218 406046 342758 406102
rect 342814 406046 342882 406102
rect 342938 406046 373478 406102
rect 373534 406046 373602 406102
rect 373658 406046 404198 406102
rect 404254 406046 404322 406102
rect 404378 406046 434918 406102
rect 434974 406046 435042 406102
rect 435098 406046 465638 406102
rect 465694 406046 465762 406102
rect 465818 406046 496358 406102
rect 496414 406046 496482 406102
rect 496538 406046 510970 406102
rect 511026 406046 511094 406102
rect 511150 406046 511218 406102
rect 511274 406046 511342 406102
rect 511398 406046 528970 406102
rect 529026 406046 529094 406102
rect 529150 406046 529218 406102
rect 529274 406046 529342 406102
rect 529398 406046 546970 406102
rect 547026 406046 547094 406102
rect 547150 406046 547218 406102
rect 547274 406046 547342 406102
rect 547398 406046 564970 406102
rect 565026 406046 565094 406102
rect 565150 406046 565218 406102
rect 565274 406046 565342 406102
rect 565398 406046 582970 406102
rect 583026 406046 583094 406102
rect 583150 406046 583218 406102
rect 583274 406046 583342 406102
rect 583398 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 6970 405978
rect 7026 405922 7094 405978
rect 7150 405922 7218 405978
rect 7274 405922 7342 405978
rect 7398 405922 24970 405978
rect 25026 405922 25094 405978
rect 25150 405922 25218 405978
rect 25274 405922 25342 405978
rect 25398 405922 42970 405978
rect 43026 405922 43094 405978
rect 43150 405922 43218 405978
rect 43274 405922 43342 405978
rect 43398 405922 60970 405978
rect 61026 405922 61094 405978
rect 61150 405922 61218 405978
rect 61274 405922 61342 405978
rect 61398 405922 78970 405978
rect 79026 405922 79094 405978
rect 79150 405922 79218 405978
rect 79274 405922 79342 405978
rect 79398 405922 96970 405978
rect 97026 405922 97094 405978
rect 97150 405922 97218 405978
rect 97274 405922 97342 405978
rect 97398 405922 114970 405978
rect 115026 405922 115094 405978
rect 115150 405922 115218 405978
rect 115274 405922 115342 405978
rect 115398 405922 132970 405978
rect 133026 405922 133094 405978
rect 133150 405922 133218 405978
rect 133274 405922 133342 405978
rect 133398 405922 150970 405978
rect 151026 405922 151094 405978
rect 151150 405922 151218 405978
rect 151274 405922 151342 405978
rect 151398 405922 168970 405978
rect 169026 405922 169094 405978
rect 169150 405922 169218 405978
rect 169274 405922 169342 405978
rect 169398 405922 186970 405978
rect 187026 405922 187094 405978
rect 187150 405922 187218 405978
rect 187274 405922 187342 405978
rect 187398 405922 219878 405978
rect 219934 405922 220002 405978
rect 220058 405922 250598 405978
rect 250654 405922 250722 405978
rect 250778 405922 281318 405978
rect 281374 405922 281442 405978
rect 281498 405922 312038 405978
rect 312094 405922 312162 405978
rect 312218 405922 342758 405978
rect 342814 405922 342882 405978
rect 342938 405922 373478 405978
rect 373534 405922 373602 405978
rect 373658 405922 404198 405978
rect 404254 405922 404322 405978
rect 404378 405922 434918 405978
rect 434974 405922 435042 405978
rect 435098 405922 465638 405978
rect 465694 405922 465762 405978
rect 465818 405922 496358 405978
rect 496414 405922 496482 405978
rect 496538 405922 510970 405978
rect 511026 405922 511094 405978
rect 511150 405922 511218 405978
rect 511274 405922 511342 405978
rect 511398 405922 528970 405978
rect 529026 405922 529094 405978
rect 529150 405922 529218 405978
rect 529274 405922 529342 405978
rect 529398 405922 546970 405978
rect 547026 405922 547094 405978
rect 547150 405922 547218 405978
rect 547274 405922 547342 405978
rect 547398 405922 564970 405978
rect 565026 405922 565094 405978
rect 565150 405922 565218 405978
rect 565274 405922 565342 405978
rect 565398 405922 582970 405978
rect 583026 405922 583094 405978
rect 583150 405922 583218 405978
rect 583274 405922 583342 405978
rect 583398 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 3250 400350
rect 3306 400294 3374 400350
rect 3430 400294 3498 400350
rect 3554 400294 3622 400350
rect 3678 400294 21250 400350
rect 21306 400294 21374 400350
rect 21430 400294 21498 400350
rect 21554 400294 21622 400350
rect 21678 400294 39250 400350
rect 39306 400294 39374 400350
rect 39430 400294 39498 400350
rect 39554 400294 39622 400350
rect 39678 400294 57250 400350
rect 57306 400294 57374 400350
rect 57430 400294 57498 400350
rect 57554 400294 57622 400350
rect 57678 400294 75250 400350
rect 75306 400294 75374 400350
rect 75430 400294 75498 400350
rect 75554 400294 75622 400350
rect 75678 400294 93250 400350
rect 93306 400294 93374 400350
rect 93430 400294 93498 400350
rect 93554 400294 93622 400350
rect 93678 400294 111250 400350
rect 111306 400294 111374 400350
rect 111430 400294 111498 400350
rect 111554 400294 111622 400350
rect 111678 400294 129250 400350
rect 129306 400294 129374 400350
rect 129430 400294 129498 400350
rect 129554 400294 129622 400350
rect 129678 400294 147250 400350
rect 147306 400294 147374 400350
rect 147430 400294 147498 400350
rect 147554 400294 147622 400350
rect 147678 400294 165250 400350
rect 165306 400294 165374 400350
rect 165430 400294 165498 400350
rect 165554 400294 165622 400350
rect 165678 400294 183250 400350
rect 183306 400294 183374 400350
rect 183430 400294 183498 400350
rect 183554 400294 183622 400350
rect 183678 400294 201250 400350
rect 201306 400294 201374 400350
rect 201430 400294 201498 400350
rect 201554 400294 201622 400350
rect 201678 400294 204518 400350
rect 204574 400294 204642 400350
rect 204698 400294 235238 400350
rect 235294 400294 235362 400350
rect 235418 400294 265958 400350
rect 266014 400294 266082 400350
rect 266138 400294 296678 400350
rect 296734 400294 296802 400350
rect 296858 400294 327398 400350
rect 327454 400294 327522 400350
rect 327578 400294 358118 400350
rect 358174 400294 358242 400350
rect 358298 400294 388838 400350
rect 388894 400294 388962 400350
rect 389018 400294 419558 400350
rect 419614 400294 419682 400350
rect 419738 400294 450278 400350
rect 450334 400294 450402 400350
rect 450458 400294 480998 400350
rect 481054 400294 481122 400350
rect 481178 400294 507250 400350
rect 507306 400294 507374 400350
rect 507430 400294 507498 400350
rect 507554 400294 507622 400350
rect 507678 400294 525250 400350
rect 525306 400294 525374 400350
rect 525430 400294 525498 400350
rect 525554 400294 525622 400350
rect 525678 400294 543250 400350
rect 543306 400294 543374 400350
rect 543430 400294 543498 400350
rect 543554 400294 543622 400350
rect 543678 400294 561250 400350
rect 561306 400294 561374 400350
rect 561430 400294 561498 400350
rect 561554 400294 561622 400350
rect 561678 400294 579250 400350
rect 579306 400294 579374 400350
rect 579430 400294 579498 400350
rect 579554 400294 579622 400350
rect 579678 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 3250 400226
rect 3306 400170 3374 400226
rect 3430 400170 3498 400226
rect 3554 400170 3622 400226
rect 3678 400170 21250 400226
rect 21306 400170 21374 400226
rect 21430 400170 21498 400226
rect 21554 400170 21622 400226
rect 21678 400170 39250 400226
rect 39306 400170 39374 400226
rect 39430 400170 39498 400226
rect 39554 400170 39622 400226
rect 39678 400170 57250 400226
rect 57306 400170 57374 400226
rect 57430 400170 57498 400226
rect 57554 400170 57622 400226
rect 57678 400170 75250 400226
rect 75306 400170 75374 400226
rect 75430 400170 75498 400226
rect 75554 400170 75622 400226
rect 75678 400170 93250 400226
rect 93306 400170 93374 400226
rect 93430 400170 93498 400226
rect 93554 400170 93622 400226
rect 93678 400170 111250 400226
rect 111306 400170 111374 400226
rect 111430 400170 111498 400226
rect 111554 400170 111622 400226
rect 111678 400170 129250 400226
rect 129306 400170 129374 400226
rect 129430 400170 129498 400226
rect 129554 400170 129622 400226
rect 129678 400170 147250 400226
rect 147306 400170 147374 400226
rect 147430 400170 147498 400226
rect 147554 400170 147622 400226
rect 147678 400170 165250 400226
rect 165306 400170 165374 400226
rect 165430 400170 165498 400226
rect 165554 400170 165622 400226
rect 165678 400170 183250 400226
rect 183306 400170 183374 400226
rect 183430 400170 183498 400226
rect 183554 400170 183622 400226
rect 183678 400170 201250 400226
rect 201306 400170 201374 400226
rect 201430 400170 201498 400226
rect 201554 400170 201622 400226
rect 201678 400170 204518 400226
rect 204574 400170 204642 400226
rect 204698 400170 235238 400226
rect 235294 400170 235362 400226
rect 235418 400170 265958 400226
rect 266014 400170 266082 400226
rect 266138 400170 296678 400226
rect 296734 400170 296802 400226
rect 296858 400170 327398 400226
rect 327454 400170 327522 400226
rect 327578 400170 358118 400226
rect 358174 400170 358242 400226
rect 358298 400170 388838 400226
rect 388894 400170 388962 400226
rect 389018 400170 419558 400226
rect 419614 400170 419682 400226
rect 419738 400170 450278 400226
rect 450334 400170 450402 400226
rect 450458 400170 480998 400226
rect 481054 400170 481122 400226
rect 481178 400170 507250 400226
rect 507306 400170 507374 400226
rect 507430 400170 507498 400226
rect 507554 400170 507622 400226
rect 507678 400170 525250 400226
rect 525306 400170 525374 400226
rect 525430 400170 525498 400226
rect 525554 400170 525622 400226
rect 525678 400170 543250 400226
rect 543306 400170 543374 400226
rect 543430 400170 543498 400226
rect 543554 400170 543622 400226
rect 543678 400170 561250 400226
rect 561306 400170 561374 400226
rect 561430 400170 561498 400226
rect 561554 400170 561622 400226
rect 561678 400170 579250 400226
rect 579306 400170 579374 400226
rect 579430 400170 579498 400226
rect 579554 400170 579622 400226
rect 579678 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 3250 400102
rect 3306 400046 3374 400102
rect 3430 400046 3498 400102
rect 3554 400046 3622 400102
rect 3678 400046 21250 400102
rect 21306 400046 21374 400102
rect 21430 400046 21498 400102
rect 21554 400046 21622 400102
rect 21678 400046 39250 400102
rect 39306 400046 39374 400102
rect 39430 400046 39498 400102
rect 39554 400046 39622 400102
rect 39678 400046 57250 400102
rect 57306 400046 57374 400102
rect 57430 400046 57498 400102
rect 57554 400046 57622 400102
rect 57678 400046 75250 400102
rect 75306 400046 75374 400102
rect 75430 400046 75498 400102
rect 75554 400046 75622 400102
rect 75678 400046 93250 400102
rect 93306 400046 93374 400102
rect 93430 400046 93498 400102
rect 93554 400046 93622 400102
rect 93678 400046 111250 400102
rect 111306 400046 111374 400102
rect 111430 400046 111498 400102
rect 111554 400046 111622 400102
rect 111678 400046 129250 400102
rect 129306 400046 129374 400102
rect 129430 400046 129498 400102
rect 129554 400046 129622 400102
rect 129678 400046 147250 400102
rect 147306 400046 147374 400102
rect 147430 400046 147498 400102
rect 147554 400046 147622 400102
rect 147678 400046 165250 400102
rect 165306 400046 165374 400102
rect 165430 400046 165498 400102
rect 165554 400046 165622 400102
rect 165678 400046 183250 400102
rect 183306 400046 183374 400102
rect 183430 400046 183498 400102
rect 183554 400046 183622 400102
rect 183678 400046 201250 400102
rect 201306 400046 201374 400102
rect 201430 400046 201498 400102
rect 201554 400046 201622 400102
rect 201678 400046 204518 400102
rect 204574 400046 204642 400102
rect 204698 400046 235238 400102
rect 235294 400046 235362 400102
rect 235418 400046 265958 400102
rect 266014 400046 266082 400102
rect 266138 400046 296678 400102
rect 296734 400046 296802 400102
rect 296858 400046 327398 400102
rect 327454 400046 327522 400102
rect 327578 400046 358118 400102
rect 358174 400046 358242 400102
rect 358298 400046 388838 400102
rect 388894 400046 388962 400102
rect 389018 400046 419558 400102
rect 419614 400046 419682 400102
rect 419738 400046 450278 400102
rect 450334 400046 450402 400102
rect 450458 400046 480998 400102
rect 481054 400046 481122 400102
rect 481178 400046 507250 400102
rect 507306 400046 507374 400102
rect 507430 400046 507498 400102
rect 507554 400046 507622 400102
rect 507678 400046 525250 400102
rect 525306 400046 525374 400102
rect 525430 400046 525498 400102
rect 525554 400046 525622 400102
rect 525678 400046 543250 400102
rect 543306 400046 543374 400102
rect 543430 400046 543498 400102
rect 543554 400046 543622 400102
rect 543678 400046 561250 400102
rect 561306 400046 561374 400102
rect 561430 400046 561498 400102
rect 561554 400046 561622 400102
rect 561678 400046 579250 400102
rect 579306 400046 579374 400102
rect 579430 400046 579498 400102
rect 579554 400046 579622 400102
rect 579678 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 3250 399978
rect 3306 399922 3374 399978
rect 3430 399922 3498 399978
rect 3554 399922 3622 399978
rect 3678 399922 21250 399978
rect 21306 399922 21374 399978
rect 21430 399922 21498 399978
rect 21554 399922 21622 399978
rect 21678 399922 39250 399978
rect 39306 399922 39374 399978
rect 39430 399922 39498 399978
rect 39554 399922 39622 399978
rect 39678 399922 57250 399978
rect 57306 399922 57374 399978
rect 57430 399922 57498 399978
rect 57554 399922 57622 399978
rect 57678 399922 75250 399978
rect 75306 399922 75374 399978
rect 75430 399922 75498 399978
rect 75554 399922 75622 399978
rect 75678 399922 93250 399978
rect 93306 399922 93374 399978
rect 93430 399922 93498 399978
rect 93554 399922 93622 399978
rect 93678 399922 111250 399978
rect 111306 399922 111374 399978
rect 111430 399922 111498 399978
rect 111554 399922 111622 399978
rect 111678 399922 129250 399978
rect 129306 399922 129374 399978
rect 129430 399922 129498 399978
rect 129554 399922 129622 399978
rect 129678 399922 147250 399978
rect 147306 399922 147374 399978
rect 147430 399922 147498 399978
rect 147554 399922 147622 399978
rect 147678 399922 165250 399978
rect 165306 399922 165374 399978
rect 165430 399922 165498 399978
rect 165554 399922 165622 399978
rect 165678 399922 183250 399978
rect 183306 399922 183374 399978
rect 183430 399922 183498 399978
rect 183554 399922 183622 399978
rect 183678 399922 201250 399978
rect 201306 399922 201374 399978
rect 201430 399922 201498 399978
rect 201554 399922 201622 399978
rect 201678 399922 204518 399978
rect 204574 399922 204642 399978
rect 204698 399922 235238 399978
rect 235294 399922 235362 399978
rect 235418 399922 265958 399978
rect 266014 399922 266082 399978
rect 266138 399922 296678 399978
rect 296734 399922 296802 399978
rect 296858 399922 327398 399978
rect 327454 399922 327522 399978
rect 327578 399922 358118 399978
rect 358174 399922 358242 399978
rect 358298 399922 388838 399978
rect 388894 399922 388962 399978
rect 389018 399922 419558 399978
rect 419614 399922 419682 399978
rect 419738 399922 450278 399978
rect 450334 399922 450402 399978
rect 450458 399922 480998 399978
rect 481054 399922 481122 399978
rect 481178 399922 507250 399978
rect 507306 399922 507374 399978
rect 507430 399922 507498 399978
rect 507554 399922 507622 399978
rect 507678 399922 525250 399978
rect 525306 399922 525374 399978
rect 525430 399922 525498 399978
rect 525554 399922 525622 399978
rect 525678 399922 543250 399978
rect 543306 399922 543374 399978
rect 543430 399922 543498 399978
rect 543554 399922 543622 399978
rect 543678 399922 561250 399978
rect 561306 399922 561374 399978
rect 561430 399922 561498 399978
rect 561554 399922 561622 399978
rect 561678 399922 579250 399978
rect 579306 399922 579374 399978
rect 579430 399922 579498 399978
rect 579554 399922 579622 399978
rect 579678 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 6970 388350
rect 7026 388294 7094 388350
rect 7150 388294 7218 388350
rect 7274 388294 7342 388350
rect 7398 388294 24970 388350
rect 25026 388294 25094 388350
rect 25150 388294 25218 388350
rect 25274 388294 25342 388350
rect 25398 388294 42970 388350
rect 43026 388294 43094 388350
rect 43150 388294 43218 388350
rect 43274 388294 43342 388350
rect 43398 388294 60970 388350
rect 61026 388294 61094 388350
rect 61150 388294 61218 388350
rect 61274 388294 61342 388350
rect 61398 388294 78970 388350
rect 79026 388294 79094 388350
rect 79150 388294 79218 388350
rect 79274 388294 79342 388350
rect 79398 388294 96970 388350
rect 97026 388294 97094 388350
rect 97150 388294 97218 388350
rect 97274 388294 97342 388350
rect 97398 388294 114970 388350
rect 115026 388294 115094 388350
rect 115150 388294 115218 388350
rect 115274 388294 115342 388350
rect 115398 388294 132970 388350
rect 133026 388294 133094 388350
rect 133150 388294 133218 388350
rect 133274 388294 133342 388350
rect 133398 388294 150970 388350
rect 151026 388294 151094 388350
rect 151150 388294 151218 388350
rect 151274 388294 151342 388350
rect 151398 388294 168970 388350
rect 169026 388294 169094 388350
rect 169150 388294 169218 388350
rect 169274 388294 169342 388350
rect 169398 388294 186970 388350
rect 187026 388294 187094 388350
rect 187150 388294 187218 388350
rect 187274 388294 187342 388350
rect 187398 388294 219878 388350
rect 219934 388294 220002 388350
rect 220058 388294 250598 388350
rect 250654 388294 250722 388350
rect 250778 388294 281318 388350
rect 281374 388294 281442 388350
rect 281498 388294 312038 388350
rect 312094 388294 312162 388350
rect 312218 388294 342758 388350
rect 342814 388294 342882 388350
rect 342938 388294 373478 388350
rect 373534 388294 373602 388350
rect 373658 388294 404198 388350
rect 404254 388294 404322 388350
rect 404378 388294 434918 388350
rect 434974 388294 435042 388350
rect 435098 388294 465638 388350
rect 465694 388294 465762 388350
rect 465818 388294 496358 388350
rect 496414 388294 496482 388350
rect 496538 388294 510970 388350
rect 511026 388294 511094 388350
rect 511150 388294 511218 388350
rect 511274 388294 511342 388350
rect 511398 388294 528970 388350
rect 529026 388294 529094 388350
rect 529150 388294 529218 388350
rect 529274 388294 529342 388350
rect 529398 388294 546970 388350
rect 547026 388294 547094 388350
rect 547150 388294 547218 388350
rect 547274 388294 547342 388350
rect 547398 388294 564970 388350
rect 565026 388294 565094 388350
rect 565150 388294 565218 388350
rect 565274 388294 565342 388350
rect 565398 388294 582970 388350
rect 583026 388294 583094 388350
rect 583150 388294 583218 388350
rect 583274 388294 583342 388350
rect 583398 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 6970 388226
rect 7026 388170 7094 388226
rect 7150 388170 7218 388226
rect 7274 388170 7342 388226
rect 7398 388170 24970 388226
rect 25026 388170 25094 388226
rect 25150 388170 25218 388226
rect 25274 388170 25342 388226
rect 25398 388170 42970 388226
rect 43026 388170 43094 388226
rect 43150 388170 43218 388226
rect 43274 388170 43342 388226
rect 43398 388170 60970 388226
rect 61026 388170 61094 388226
rect 61150 388170 61218 388226
rect 61274 388170 61342 388226
rect 61398 388170 78970 388226
rect 79026 388170 79094 388226
rect 79150 388170 79218 388226
rect 79274 388170 79342 388226
rect 79398 388170 96970 388226
rect 97026 388170 97094 388226
rect 97150 388170 97218 388226
rect 97274 388170 97342 388226
rect 97398 388170 114970 388226
rect 115026 388170 115094 388226
rect 115150 388170 115218 388226
rect 115274 388170 115342 388226
rect 115398 388170 132970 388226
rect 133026 388170 133094 388226
rect 133150 388170 133218 388226
rect 133274 388170 133342 388226
rect 133398 388170 150970 388226
rect 151026 388170 151094 388226
rect 151150 388170 151218 388226
rect 151274 388170 151342 388226
rect 151398 388170 168970 388226
rect 169026 388170 169094 388226
rect 169150 388170 169218 388226
rect 169274 388170 169342 388226
rect 169398 388170 186970 388226
rect 187026 388170 187094 388226
rect 187150 388170 187218 388226
rect 187274 388170 187342 388226
rect 187398 388170 219878 388226
rect 219934 388170 220002 388226
rect 220058 388170 250598 388226
rect 250654 388170 250722 388226
rect 250778 388170 281318 388226
rect 281374 388170 281442 388226
rect 281498 388170 312038 388226
rect 312094 388170 312162 388226
rect 312218 388170 342758 388226
rect 342814 388170 342882 388226
rect 342938 388170 373478 388226
rect 373534 388170 373602 388226
rect 373658 388170 404198 388226
rect 404254 388170 404322 388226
rect 404378 388170 434918 388226
rect 434974 388170 435042 388226
rect 435098 388170 465638 388226
rect 465694 388170 465762 388226
rect 465818 388170 496358 388226
rect 496414 388170 496482 388226
rect 496538 388170 510970 388226
rect 511026 388170 511094 388226
rect 511150 388170 511218 388226
rect 511274 388170 511342 388226
rect 511398 388170 528970 388226
rect 529026 388170 529094 388226
rect 529150 388170 529218 388226
rect 529274 388170 529342 388226
rect 529398 388170 546970 388226
rect 547026 388170 547094 388226
rect 547150 388170 547218 388226
rect 547274 388170 547342 388226
rect 547398 388170 564970 388226
rect 565026 388170 565094 388226
rect 565150 388170 565218 388226
rect 565274 388170 565342 388226
rect 565398 388170 582970 388226
rect 583026 388170 583094 388226
rect 583150 388170 583218 388226
rect 583274 388170 583342 388226
rect 583398 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 6970 388102
rect 7026 388046 7094 388102
rect 7150 388046 7218 388102
rect 7274 388046 7342 388102
rect 7398 388046 24970 388102
rect 25026 388046 25094 388102
rect 25150 388046 25218 388102
rect 25274 388046 25342 388102
rect 25398 388046 42970 388102
rect 43026 388046 43094 388102
rect 43150 388046 43218 388102
rect 43274 388046 43342 388102
rect 43398 388046 60970 388102
rect 61026 388046 61094 388102
rect 61150 388046 61218 388102
rect 61274 388046 61342 388102
rect 61398 388046 78970 388102
rect 79026 388046 79094 388102
rect 79150 388046 79218 388102
rect 79274 388046 79342 388102
rect 79398 388046 96970 388102
rect 97026 388046 97094 388102
rect 97150 388046 97218 388102
rect 97274 388046 97342 388102
rect 97398 388046 114970 388102
rect 115026 388046 115094 388102
rect 115150 388046 115218 388102
rect 115274 388046 115342 388102
rect 115398 388046 132970 388102
rect 133026 388046 133094 388102
rect 133150 388046 133218 388102
rect 133274 388046 133342 388102
rect 133398 388046 150970 388102
rect 151026 388046 151094 388102
rect 151150 388046 151218 388102
rect 151274 388046 151342 388102
rect 151398 388046 168970 388102
rect 169026 388046 169094 388102
rect 169150 388046 169218 388102
rect 169274 388046 169342 388102
rect 169398 388046 186970 388102
rect 187026 388046 187094 388102
rect 187150 388046 187218 388102
rect 187274 388046 187342 388102
rect 187398 388046 219878 388102
rect 219934 388046 220002 388102
rect 220058 388046 250598 388102
rect 250654 388046 250722 388102
rect 250778 388046 281318 388102
rect 281374 388046 281442 388102
rect 281498 388046 312038 388102
rect 312094 388046 312162 388102
rect 312218 388046 342758 388102
rect 342814 388046 342882 388102
rect 342938 388046 373478 388102
rect 373534 388046 373602 388102
rect 373658 388046 404198 388102
rect 404254 388046 404322 388102
rect 404378 388046 434918 388102
rect 434974 388046 435042 388102
rect 435098 388046 465638 388102
rect 465694 388046 465762 388102
rect 465818 388046 496358 388102
rect 496414 388046 496482 388102
rect 496538 388046 510970 388102
rect 511026 388046 511094 388102
rect 511150 388046 511218 388102
rect 511274 388046 511342 388102
rect 511398 388046 528970 388102
rect 529026 388046 529094 388102
rect 529150 388046 529218 388102
rect 529274 388046 529342 388102
rect 529398 388046 546970 388102
rect 547026 388046 547094 388102
rect 547150 388046 547218 388102
rect 547274 388046 547342 388102
rect 547398 388046 564970 388102
rect 565026 388046 565094 388102
rect 565150 388046 565218 388102
rect 565274 388046 565342 388102
rect 565398 388046 582970 388102
rect 583026 388046 583094 388102
rect 583150 388046 583218 388102
rect 583274 388046 583342 388102
rect 583398 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 6970 387978
rect 7026 387922 7094 387978
rect 7150 387922 7218 387978
rect 7274 387922 7342 387978
rect 7398 387922 24970 387978
rect 25026 387922 25094 387978
rect 25150 387922 25218 387978
rect 25274 387922 25342 387978
rect 25398 387922 42970 387978
rect 43026 387922 43094 387978
rect 43150 387922 43218 387978
rect 43274 387922 43342 387978
rect 43398 387922 60970 387978
rect 61026 387922 61094 387978
rect 61150 387922 61218 387978
rect 61274 387922 61342 387978
rect 61398 387922 78970 387978
rect 79026 387922 79094 387978
rect 79150 387922 79218 387978
rect 79274 387922 79342 387978
rect 79398 387922 96970 387978
rect 97026 387922 97094 387978
rect 97150 387922 97218 387978
rect 97274 387922 97342 387978
rect 97398 387922 114970 387978
rect 115026 387922 115094 387978
rect 115150 387922 115218 387978
rect 115274 387922 115342 387978
rect 115398 387922 132970 387978
rect 133026 387922 133094 387978
rect 133150 387922 133218 387978
rect 133274 387922 133342 387978
rect 133398 387922 150970 387978
rect 151026 387922 151094 387978
rect 151150 387922 151218 387978
rect 151274 387922 151342 387978
rect 151398 387922 168970 387978
rect 169026 387922 169094 387978
rect 169150 387922 169218 387978
rect 169274 387922 169342 387978
rect 169398 387922 186970 387978
rect 187026 387922 187094 387978
rect 187150 387922 187218 387978
rect 187274 387922 187342 387978
rect 187398 387922 219878 387978
rect 219934 387922 220002 387978
rect 220058 387922 250598 387978
rect 250654 387922 250722 387978
rect 250778 387922 281318 387978
rect 281374 387922 281442 387978
rect 281498 387922 312038 387978
rect 312094 387922 312162 387978
rect 312218 387922 342758 387978
rect 342814 387922 342882 387978
rect 342938 387922 373478 387978
rect 373534 387922 373602 387978
rect 373658 387922 404198 387978
rect 404254 387922 404322 387978
rect 404378 387922 434918 387978
rect 434974 387922 435042 387978
rect 435098 387922 465638 387978
rect 465694 387922 465762 387978
rect 465818 387922 496358 387978
rect 496414 387922 496482 387978
rect 496538 387922 510970 387978
rect 511026 387922 511094 387978
rect 511150 387922 511218 387978
rect 511274 387922 511342 387978
rect 511398 387922 528970 387978
rect 529026 387922 529094 387978
rect 529150 387922 529218 387978
rect 529274 387922 529342 387978
rect 529398 387922 546970 387978
rect 547026 387922 547094 387978
rect 547150 387922 547218 387978
rect 547274 387922 547342 387978
rect 547398 387922 564970 387978
rect 565026 387922 565094 387978
rect 565150 387922 565218 387978
rect 565274 387922 565342 387978
rect 565398 387922 582970 387978
rect 583026 387922 583094 387978
rect 583150 387922 583218 387978
rect 583274 387922 583342 387978
rect 583398 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 3250 382350
rect 3306 382294 3374 382350
rect 3430 382294 3498 382350
rect 3554 382294 3622 382350
rect 3678 382294 21250 382350
rect 21306 382294 21374 382350
rect 21430 382294 21498 382350
rect 21554 382294 21622 382350
rect 21678 382294 39250 382350
rect 39306 382294 39374 382350
rect 39430 382294 39498 382350
rect 39554 382294 39622 382350
rect 39678 382294 57250 382350
rect 57306 382294 57374 382350
rect 57430 382294 57498 382350
rect 57554 382294 57622 382350
rect 57678 382294 75250 382350
rect 75306 382294 75374 382350
rect 75430 382294 75498 382350
rect 75554 382294 75622 382350
rect 75678 382294 93250 382350
rect 93306 382294 93374 382350
rect 93430 382294 93498 382350
rect 93554 382294 93622 382350
rect 93678 382294 111250 382350
rect 111306 382294 111374 382350
rect 111430 382294 111498 382350
rect 111554 382294 111622 382350
rect 111678 382294 129250 382350
rect 129306 382294 129374 382350
rect 129430 382294 129498 382350
rect 129554 382294 129622 382350
rect 129678 382294 147250 382350
rect 147306 382294 147374 382350
rect 147430 382294 147498 382350
rect 147554 382294 147622 382350
rect 147678 382294 165250 382350
rect 165306 382294 165374 382350
rect 165430 382294 165498 382350
rect 165554 382294 165622 382350
rect 165678 382294 183250 382350
rect 183306 382294 183374 382350
rect 183430 382294 183498 382350
rect 183554 382294 183622 382350
rect 183678 382294 201250 382350
rect 201306 382294 201374 382350
rect 201430 382294 201498 382350
rect 201554 382294 201622 382350
rect 201678 382294 204518 382350
rect 204574 382294 204642 382350
rect 204698 382294 235238 382350
rect 235294 382294 235362 382350
rect 235418 382294 265958 382350
rect 266014 382294 266082 382350
rect 266138 382294 296678 382350
rect 296734 382294 296802 382350
rect 296858 382294 327398 382350
rect 327454 382294 327522 382350
rect 327578 382294 358118 382350
rect 358174 382294 358242 382350
rect 358298 382294 388838 382350
rect 388894 382294 388962 382350
rect 389018 382294 419558 382350
rect 419614 382294 419682 382350
rect 419738 382294 450278 382350
rect 450334 382294 450402 382350
rect 450458 382294 480998 382350
rect 481054 382294 481122 382350
rect 481178 382294 507250 382350
rect 507306 382294 507374 382350
rect 507430 382294 507498 382350
rect 507554 382294 507622 382350
rect 507678 382294 525250 382350
rect 525306 382294 525374 382350
rect 525430 382294 525498 382350
rect 525554 382294 525622 382350
rect 525678 382294 543250 382350
rect 543306 382294 543374 382350
rect 543430 382294 543498 382350
rect 543554 382294 543622 382350
rect 543678 382294 561250 382350
rect 561306 382294 561374 382350
rect 561430 382294 561498 382350
rect 561554 382294 561622 382350
rect 561678 382294 579250 382350
rect 579306 382294 579374 382350
rect 579430 382294 579498 382350
rect 579554 382294 579622 382350
rect 579678 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 3250 382226
rect 3306 382170 3374 382226
rect 3430 382170 3498 382226
rect 3554 382170 3622 382226
rect 3678 382170 21250 382226
rect 21306 382170 21374 382226
rect 21430 382170 21498 382226
rect 21554 382170 21622 382226
rect 21678 382170 39250 382226
rect 39306 382170 39374 382226
rect 39430 382170 39498 382226
rect 39554 382170 39622 382226
rect 39678 382170 57250 382226
rect 57306 382170 57374 382226
rect 57430 382170 57498 382226
rect 57554 382170 57622 382226
rect 57678 382170 75250 382226
rect 75306 382170 75374 382226
rect 75430 382170 75498 382226
rect 75554 382170 75622 382226
rect 75678 382170 93250 382226
rect 93306 382170 93374 382226
rect 93430 382170 93498 382226
rect 93554 382170 93622 382226
rect 93678 382170 111250 382226
rect 111306 382170 111374 382226
rect 111430 382170 111498 382226
rect 111554 382170 111622 382226
rect 111678 382170 129250 382226
rect 129306 382170 129374 382226
rect 129430 382170 129498 382226
rect 129554 382170 129622 382226
rect 129678 382170 147250 382226
rect 147306 382170 147374 382226
rect 147430 382170 147498 382226
rect 147554 382170 147622 382226
rect 147678 382170 165250 382226
rect 165306 382170 165374 382226
rect 165430 382170 165498 382226
rect 165554 382170 165622 382226
rect 165678 382170 183250 382226
rect 183306 382170 183374 382226
rect 183430 382170 183498 382226
rect 183554 382170 183622 382226
rect 183678 382170 201250 382226
rect 201306 382170 201374 382226
rect 201430 382170 201498 382226
rect 201554 382170 201622 382226
rect 201678 382170 204518 382226
rect 204574 382170 204642 382226
rect 204698 382170 235238 382226
rect 235294 382170 235362 382226
rect 235418 382170 265958 382226
rect 266014 382170 266082 382226
rect 266138 382170 296678 382226
rect 296734 382170 296802 382226
rect 296858 382170 327398 382226
rect 327454 382170 327522 382226
rect 327578 382170 358118 382226
rect 358174 382170 358242 382226
rect 358298 382170 388838 382226
rect 388894 382170 388962 382226
rect 389018 382170 419558 382226
rect 419614 382170 419682 382226
rect 419738 382170 450278 382226
rect 450334 382170 450402 382226
rect 450458 382170 480998 382226
rect 481054 382170 481122 382226
rect 481178 382170 507250 382226
rect 507306 382170 507374 382226
rect 507430 382170 507498 382226
rect 507554 382170 507622 382226
rect 507678 382170 525250 382226
rect 525306 382170 525374 382226
rect 525430 382170 525498 382226
rect 525554 382170 525622 382226
rect 525678 382170 543250 382226
rect 543306 382170 543374 382226
rect 543430 382170 543498 382226
rect 543554 382170 543622 382226
rect 543678 382170 561250 382226
rect 561306 382170 561374 382226
rect 561430 382170 561498 382226
rect 561554 382170 561622 382226
rect 561678 382170 579250 382226
rect 579306 382170 579374 382226
rect 579430 382170 579498 382226
rect 579554 382170 579622 382226
rect 579678 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 3250 382102
rect 3306 382046 3374 382102
rect 3430 382046 3498 382102
rect 3554 382046 3622 382102
rect 3678 382046 21250 382102
rect 21306 382046 21374 382102
rect 21430 382046 21498 382102
rect 21554 382046 21622 382102
rect 21678 382046 39250 382102
rect 39306 382046 39374 382102
rect 39430 382046 39498 382102
rect 39554 382046 39622 382102
rect 39678 382046 57250 382102
rect 57306 382046 57374 382102
rect 57430 382046 57498 382102
rect 57554 382046 57622 382102
rect 57678 382046 75250 382102
rect 75306 382046 75374 382102
rect 75430 382046 75498 382102
rect 75554 382046 75622 382102
rect 75678 382046 93250 382102
rect 93306 382046 93374 382102
rect 93430 382046 93498 382102
rect 93554 382046 93622 382102
rect 93678 382046 111250 382102
rect 111306 382046 111374 382102
rect 111430 382046 111498 382102
rect 111554 382046 111622 382102
rect 111678 382046 129250 382102
rect 129306 382046 129374 382102
rect 129430 382046 129498 382102
rect 129554 382046 129622 382102
rect 129678 382046 147250 382102
rect 147306 382046 147374 382102
rect 147430 382046 147498 382102
rect 147554 382046 147622 382102
rect 147678 382046 165250 382102
rect 165306 382046 165374 382102
rect 165430 382046 165498 382102
rect 165554 382046 165622 382102
rect 165678 382046 183250 382102
rect 183306 382046 183374 382102
rect 183430 382046 183498 382102
rect 183554 382046 183622 382102
rect 183678 382046 201250 382102
rect 201306 382046 201374 382102
rect 201430 382046 201498 382102
rect 201554 382046 201622 382102
rect 201678 382046 204518 382102
rect 204574 382046 204642 382102
rect 204698 382046 235238 382102
rect 235294 382046 235362 382102
rect 235418 382046 265958 382102
rect 266014 382046 266082 382102
rect 266138 382046 296678 382102
rect 296734 382046 296802 382102
rect 296858 382046 327398 382102
rect 327454 382046 327522 382102
rect 327578 382046 358118 382102
rect 358174 382046 358242 382102
rect 358298 382046 388838 382102
rect 388894 382046 388962 382102
rect 389018 382046 419558 382102
rect 419614 382046 419682 382102
rect 419738 382046 450278 382102
rect 450334 382046 450402 382102
rect 450458 382046 480998 382102
rect 481054 382046 481122 382102
rect 481178 382046 507250 382102
rect 507306 382046 507374 382102
rect 507430 382046 507498 382102
rect 507554 382046 507622 382102
rect 507678 382046 525250 382102
rect 525306 382046 525374 382102
rect 525430 382046 525498 382102
rect 525554 382046 525622 382102
rect 525678 382046 543250 382102
rect 543306 382046 543374 382102
rect 543430 382046 543498 382102
rect 543554 382046 543622 382102
rect 543678 382046 561250 382102
rect 561306 382046 561374 382102
rect 561430 382046 561498 382102
rect 561554 382046 561622 382102
rect 561678 382046 579250 382102
rect 579306 382046 579374 382102
rect 579430 382046 579498 382102
rect 579554 382046 579622 382102
rect 579678 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 3250 381978
rect 3306 381922 3374 381978
rect 3430 381922 3498 381978
rect 3554 381922 3622 381978
rect 3678 381922 21250 381978
rect 21306 381922 21374 381978
rect 21430 381922 21498 381978
rect 21554 381922 21622 381978
rect 21678 381922 39250 381978
rect 39306 381922 39374 381978
rect 39430 381922 39498 381978
rect 39554 381922 39622 381978
rect 39678 381922 57250 381978
rect 57306 381922 57374 381978
rect 57430 381922 57498 381978
rect 57554 381922 57622 381978
rect 57678 381922 75250 381978
rect 75306 381922 75374 381978
rect 75430 381922 75498 381978
rect 75554 381922 75622 381978
rect 75678 381922 93250 381978
rect 93306 381922 93374 381978
rect 93430 381922 93498 381978
rect 93554 381922 93622 381978
rect 93678 381922 111250 381978
rect 111306 381922 111374 381978
rect 111430 381922 111498 381978
rect 111554 381922 111622 381978
rect 111678 381922 129250 381978
rect 129306 381922 129374 381978
rect 129430 381922 129498 381978
rect 129554 381922 129622 381978
rect 129678 381922 147250 381978
rect 147306 381922 147374 381978
rect 147430 381922 147498 381978
rect 147554 381922 147622 381978
rect 147678 381922 165250 381978
rect 165306 381922 165374 381978
rect 165430 381922 165498 381978
rect 165554 381922 165622 381978
rect 165678 381922 183250 381978
rect 183306 381922 183374 381978
rect 183430 381922 183498 381978
rect 183554 381922 183622 381978
rect 183678 381922 201250 381978
rect 201306 381922 201374 381978
rect 201430 381922 201498 381978
rect 201554 381922 201622 381978
rect 201678 381922 204518 381978
rect 204574 381922 204642 381978
rect 204698 381922 235238 381978
rect 235294 381922 235362 381978
rect 235418 381922 265958 381978
rect 266014 381922 266082 381978
rect 266138 381922 296678 381978
rect 296734 381922 296802 381978
rect 296858 381922 327398 381978
rect 327454 381922 327522 381978
rect 327578 381922 358118 381978
rect 358174 381922 358242 381978
rect 358298 381922 388838 381978
rect 388894 381922 388962 381978
rect 389018 381922 419558 381978
rect 419614 381922 419682 381978
rect 419738 381922 450278 381978
rect 450334 381922 450402 381978
rect 450458 381922 480998 381978
rect 481054 381922 481122 381978
rect 481178 381922 507250 381978
rect 507306 381922 507374 381978
rect 507430 381922 507498 381978
rect 507554 381922 507622 381978
rect 507678 381922 525250 381978
rect 525306 381922 525374 381978
rect 525430 381922 525498 381978
rect 525554 381922 525622 381978
rect 525678 381922 543250 381978
rect 543306 381922 543374 381978
rect 543430 381922 543498 381978
rect 543554 381922 543622 381978
rect 543678 381922 561250 381978
rect 561306 381922 561374 381978
rect 561430 381922 561498 381978
rect 561554 381922 561622 381978
rect 561678 381922 579250 381978
rect 579306 381922 579374 381978
rect 579430 381922 579498 381978
rect 579554 381922 579622 381978
rect 579678 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 6970 370350
rect 7026 370294 7094 370350
rect 7150 370294 7218 370350
rect 7274 370294 7342 370350
rect 7398 370294 24970 370350
rect 25026 370294 25094 370350
rect 25150 370294 25218 370350
rect 25274 370294 25342 370350
rect 25398 370294 42970 370350
rect 43026 370294 43094 370350
rect 43150 370294 43218 370350
rect 43274 370294 43342 370350
rect 43398 370294 60970 370350
rect 61026 370294 61094 370350
rect 61150 370294 61218 370350
rect 61274 370294 61342 370350
rect 61398 370294 78970 370350
rect 79026 370294 79094 370350
rect 79150 370294 79218 370350
rect 79274 370294 79342 370350
rect 79398 370294 96970 370350
rect 97026 370294 97094 370350
rect 97150 370294 97218 370350
rect 97274 370294 97342 370350
rect 97398 370294 114970 370350
rect 115026 370294 115094 370350
rect 115150 370294 115218 370350
rect 115274 370294 115342 370350
rect 115398 370294 132970 370350
rect 133026 370294 133094 370350
rect 133150 370294 133218 370350
rect 133274 370294 133342 370350
rect 133398 370294 150970 370350
rect 151026 370294 151094 370350
rect 151150 370294 151218 370350
rect 151274 370294 151342 370350
rect 151398 370294 168970 370350
rect 169026 370294 169094 370350
rect 169150 370294 169218 370350
rect 169274 370294 169342 370350
rect 169398 370294 186970 370350
rect 187026 370294 187094 370350
rect 187150 370294 187218 370350
rect 187274 370294 187342 370350
rect 187398 370294 219878 370350
rect 219934 370294 220002 370350
rect 220058 370294 250598 370350
rect 250654 370294 250722 370350
rect 250778 370294 281318 370350
rect 281374 370294 281442 370350
rect 281498 370294 312038 370350
rect 312094 370294 312162 370350
rect 312218 370294 342758 370350
rect 342814 370294 342882 370350
rect 342938 370294 373478 370350
rect 373534 370294 373602 370350
rect 373658 370294 404198 370350
rect 404254 370294 404322 370350
rect 404378 370294 434918 370350
rect 434974 370294 435042 370350
rect 435098 370294 465638 370350
rect 465694 370294 465762 370350
rect 465818 370294 496358 370350
rect 496414 370294 496482 370350
rect 496538 370294 510970 370350
rect 511026 370294 511094 370350
rect 511150 370294 511218 370350
rect 511274 370294 511342 370350
rect 511398 370294 528970 370350
rect 529026 370294 529094 370350
rect 529150 370294 529218 370350
rect 529274 370294 529342 370350
rect 529398 370294 546970 370350
rect 547026 370294 547094 370350
rect 547150 370294 547218 370350
rect 547274 370294 547342 370350
rect 547398 370294 564970 370350
rect 565026 370294 565094 370350
rect 565150 370294 565218 370350
rect 565274 370294 565342 370350
rect 565398 370294 582970 370350
rect 583026 370294 583094 370350
rect 583150 370294 583218 370350
rect 583274 370294 583342 370350
rect 583398 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 6970 370226
rect 7026 370170 7094 370226
rect 7150 370170 7218 370226
rect 7274 370170 7342 370226
rect 7398 370170 24970 370226
rect 25026 370170 25094 370226
rect 25150 370170 25218 370226
rect 25274 370170 25342 370226
rect 25398 370170 42970 370226
rect 43026 370170 43094 370226
rect 43150 370170 43218 370226
rect 43274 370170 43342 370226
rect 43398 370170 60970 370226
rect 61026 370170 61094 370226
rect 61150 370170 61218 370226
rect 61274 370170 61342 370226
rect 61398 370170 78970 370226
rect 79026 370170 79094 370226
rect 79150 370170 79218 370226
rect 79274 370170 79342 370226
rect 79398 370170 96970 370226
rect 97026 370170 97094 370226
rect 97150 370170 97218 370226
rect 97274 370170 97342 370226
rect 97398 370170 114970 370226
rect 115026 370170 115094 370226
rect 115150 370170 115218 370226
rect 115274 370170 115342 370226
rect 115398 370170 132970 370226
rect 133026 370170 133094 370226
rect 133150 370170 133218 370226
rect 133274 370170 133342 370226
rect 133398 370170 150970 370226
rect 151026 370170 151094 370226
rect 151150 370170 151218 370226
rect 151274 370170 151342 370226
rect 151398 370170 168970 370226
rect 169026 370170 169094 370226
rect 169150 370170 169218 370226
rect 169274 370170 169342 370226
rect 169398 370170 186970 370226
rect 187026 370170 187094 370226
rect 187150 370170 187218 370226
rect 187274 370170 187342 370226
rect 187398 370170 219878 370226
rect 219934 370170 220002 370226
rect 220058 370170 250598 370226
rect 250654 370170 250722 370226
rect 250778 370170 281318 370226
rect 281374 370170 281442 370226
rect 281498 370170 312038 370226
rect 312094 370170 312162 370226
rect 312218 370170 342758 370226
rect 342814 370170 342882 370226
rect 342938 370170 373478 370226
rect 373534 370170 373602 370226
rect 373658 370170 404198 370226
rect 404254 370170 404322 370226
rect 404378 370170 434918 370226
rect 434974 370170 435042 370226
rect 435098 370170 465638 370226
rect 465694 370170 465762 370226
rect 465818 370170 496358 370226
rect 496414 370170 496482 370226
rect 496538 370170 510970 370226
rect 511026 370170 511094 370226
rect 511150 370170 511218 370226
rect 511274 370170 511342 370226
rect 511398 370170 528970 370226
rect 529026 370170 529094 370226
rect 529150 370170 529218 370226
rect 529274 370170 529342 370226
rect 529398 370170 546970 370226
rect 547026 370170 547094 370226
rect 547150 370170 547218 370226
rect 547274 370170 547342 370226
rect 547398 370170 564970 370226
rect 565026 370170 565094 370226
rect 565150 370170 565218 370226
rect 565274 370170 565342 370226
rect 565398 370170 582970 370226
rect 583026 370170 583094 370226
rect 583150 370170 583218 370226
rect 583274 370170 583342 370226
rect 583398 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 6970 370102
rect 7026 370046 7094 370102
rect 7150 370046 7218 370102
rect 7274 370046 7342 370102
rect 7398 370046 24970 370102
rect 25026 370046 25094 370102
rect 25150 370046 25218 370102
rect 25274 370046 25342 370102
rect 25398 370046 42970 370102
rect 43026 370046 43094 370102
rect 43150 370046 43218 370102
rect 43274 370046 43342 370102
rect 43398 370046 60970 370102
rect 61026 370046 61094 370102
rect 61150 370046 61218 370102
rect 61274 370046 61342 370102
rect 61398 370046 78970 370102
rect 79026 370046 79094 370102
rect 79150 370046 79218 370102
rect 79274 370046 79342 370102
rect 79398 370046 96970 370102
rect 97026 370046 97094 370102
rect 97150 370046 97218 370102
rect 97274 370046 97342 370102
rect 97398 370046 114970 370102
rect 115026 370046 115094 370102
rect 115150 370046 115218 370102
rect 115274 370046 115342 370102
rect 115398 370046 132970 370102
rect 133026 370046 133094 370102
rect 133150 370046 133218 370102
rect 133274 370046 133342 370102
rect 133398 370046 150970 370102
rect 151026 370046 151094 370102
rect 151150 370046 151218 370102
rect 151274 370046 151342 370102
rect 151398 370046 168970 370102
rect 169026 370046 169094 370102
rect 169150 370046 169218 370102
rect 169274 370046 169342 370102
rect 169398 370046 186970 370102
rect 187026 370046 187094 370102
rect 187150 370046 187218 370102
rect 187274 370046 187342 370102
rect 187398 370046 219878 370102
rect 219934 370046 220002 370102
rect 220058 370046 250598 370102
rect 250654 370046 250722 370102
rect 250778 370046 281318 370102
rect 281374 370046 281442 370102
rect 281498 370046 312038 370102
rect 312094 370046 312162 370102
rect 312218 370046 342758 370102
rect 342814 370046 342882 370102
rect 342938 370046 373478 370102
rect 373534 370046 373602 370102
rect 373658 370046 404198 370102
rect 404254 370046 404322 370102
rect 404378 370046 434918 370102
rect 434974 370046 435042 370102
rect 435098 370046 465638 370102
rect 465694 370046 465762 370102
rect 465818 370046 496358 370102
rect 496414 370046 496482 370102
rect 496538 370046 510970 370102
rect 511026 370046 511094 370102
rect 511150 370046 511218 370102
rect 511274 370046 511342 370102
rect 511398 370046 528970 370102
rect 529026 370046 529094 370102
rect 529150 370046 529218 370102
rect 529274 370046 529342 370102
rect 529398 370046 546970 370102
rect 547026 370046 547094 370102
rect 547150 370046 547218 370102
rect 547274 370046 547342 370102
rect 547398 370046 564970 370102
rect 565026 370046 565094 370102
rect 565150 370046 565218 370102
rect 565274 370046 565342 370102
rect 565398 370046 582970 370102
rect 583026 370046 583094 370102
rect 583150 370046 583218 370102
rect 583274 370046 583342 370102
rect 583398 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 6970 369978
rect 7026 369922 7094 369978
rect 7150 369922 7218 369978
rect 7274 369922 7342 369978
rect 7398 369922 24970 369978
rect 25026 369922 25094 369978
rect 25150 369922 25218 369978
rect 25274 369922 25342 369978
rect 25398 369922 42970 369978
rect 43026 369922 43094 369978
rect 43150 369922 43218 369978
rect 43274 369922 43342 369978
rect 43398 369922 60970 369978
rect 61026 369922 61094 369978
rect 61150 369922 61218 369978
rect 61274 369922 61342 369978
rect 61398 369922 78970 369978
rect 79026 369922 79094 369978
rect 79150 369922 79218 369978
rect 79274 369922 79342 369978
rect 79398 369922 96970 369978
rect 97026 369922 97094 369978
rect 97150 369922 97218 369978
rect 97274 369922 97342 369978
rect 97398 369922 114970 369978
rect 115026 369922 115094 369978
rect 115150 369922 115218 369978
rect 115274 369922 115342 369978
rect 115398 369922 132970 369978
rect 133026 369922 133094 369978
rect 133150 369922 133218 369978
rect 133274 369922 133342 369978
rect 133398 369922 150970 369978
rect 151026 369922 151094 369978
rect 151150 369922 151218 369978
rect 151274 369922 151342 369978
rect 151398 369922 168970 369978
rect 169026 369922 169094 369978
rect 169150 369922 169218 369978
rect 169274 369922 169342 369978
rect 169398 369922 186970 369978
rect 187026 369922 187094 369978
rect 187150 369922 187218 369978
rect 187274 369922 187342 369978
rect 187398 369922 219878 369978
rect 219934 369922 220002 369978
rect 220058 369922 250598 369978
rect 250654 369922 250722 369978
rect 250778 369922 281318 369978
rect 281374 369922 281442 369978
rect 281498 369922 312038 369978
rect 312094 369922 312162 369978
rect 312218 369922 342758 369978
rect 342814 369922 342882 369978
rect 342938 369922 373478 369978
rect 373534 369922 373602 369978
rect 373658 369922 404198 369978
rect 404254 369922 404322 369978
rect 404378 369922 434918 369978
rect 434974 369922 435042 369978
rect 435098 369922 465638 369978
rect 465694 369922 465762 369978
rect 465818 369922 496358 369978
rect 496414 369922 496482 369978
rect 496538 369922 510970 369978
rect 511026 369922 511094 369978
rect 511150 369922 511218 369978
rect 511274 369922 511342 369978
rect 511398 369922 528970 369978
rect 529026 369922 529094 369978
rect 529150 369922 529218 369978
rect 529274 369922 529342 369978
rect 529398 369922 546970 369978
rect 547026 369922 547094 369978
rect 547150 369922 547218 369978
rect 547274 369922 547342 369978
rect 547398 369922 564970 369978
rect 565026 369922 565094 369978
rect 565150 369922 565218 369978
rect 565274 369922 565342 369978
rect 565398 369922 582970 369978
rect 583026 369922 583094 369978
rect 583150 369922 583218 369978
rect 583274 369922 583342 369978
rect 583398 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 3250 364350
rect 3306 364294 3374 364350
rect 3430 364294 3498 364350
rect 3554 364294 3622 364350
rect 3678 364294 21250 364350
rect 21306 364294 21374 364350
rect 21430 364294 21498 364350
rect 21554 364294 21622 364350
rect 21678 364294 39250 364350
rect 39306 364294 39374 364350
rect 39430 364294 39498 364350
rect 39554 364294 39622 364350
rect 39678 364294 57250 364350
rect 57306 364294 57374 364350
rect 57430 364294 57498 364350
rect 57554 364294 57622 364350
rect 57678 364294 75250 364350
rect 75306 364294 75374 364350
rect 75430 364294 75498 364350
rect 75554 364294 75622 364350
rect 75678 364294 93250 364350
rect 93306 364294 93374 364350
rect 93430 364294 93498 364350
rect 93554 364294 93622 364350
rect 93678 364294 111250 364350
rect 111306 364294 111374 364350
rect 111430 364294 111498 364350
rect 111554 364294 111622 364350
rect 111678 364294 129250 364350
rect 129306 364294 129374 364350
rect 129430 364294 129498 364350
rect 129554 364294 129622 364350
rect 129678 364294 147250 364350
rect 147306 364294 147374 364350
rect 147430 364294 147498 364350
rect 147554 364294 147622 364350
rect 147678 364294 165250 364350
rect 165306 364294 165374 364350
rect 165430 364294 165498 364350
rect 165554 364294 165622 364350
rect 165678 364294 183250 364350
rect 183306 364294 183374 364350
rect 183430 364294 183498 364350
rect 183554 364294 183622 364350
rect 183678 364294 201250 364350
rect 201306 364294 201374 364350
rect 201430 364294 201498 364350
rect 201554 364294 201622 364350
rect 201678 364294 204518 364350
rect 204574 364294 204642 364350
rect 204698 364294 235238 364350
rect 235294 364294 235362 364350
rect 235418 364294 265958 364350
rect 266014 364294 266082 364350
rect 266138 364294 296678 364350
rect 296734 364294 296802 364350
rect 296858 364294 327398 364350
rect 327454 364294 327522 364350
rect 327578 364294 358118 364350
rect 358174 364294 358242 364350
rect 358298 364294 388838 364350
rect 388894 364294 388962 364350
rect 389018 364294 419558 364350
rect 419614 364294 419682 364350
rect 419738 364294 450278 364350
rect 450334 364294 450402 364350
rect 450458 364294 480998 364350
rect 481054 364294 481122 364350
rect 481178 364294 507250 364350
rect 507306 364294 507374 364350
rect 507430 364294 507498 364350
rect 507554 364294 507622 364350
rect 507678 364294 525250 364350
rect 525306 364294 525374 364350
rect 525430 364294 525498 364350
rect 525554 364294 525622 364350
rect 525678 364294 543250 364350
rect 543306 364294 543374 364350
rect 543430 364294 543498 364350
rect 543554 364294 543622 364350
rect 543678 364294 561250 364350
rect 561306 364294 561374 364350
rect 561430 364294 561498 364350
rect 561554 364294 561622 364350
rect 561678 364294 579250 364350
rect 579306 364294 579374 364350
rect 579430 364294 579498 364350
rect 579554 364294 579622 364350
rect 579678 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 3250 364226
rect 3306 364170 3374 364226
rect 3430 364170 3498 364226
rect 3554 364170 3622 364226
rect 3678 364170 21250 364226
rect 21306 364170 21374 364226
rect 21430 364170 21498 364226
rect 21554 364170 21622 364226
rect 21678 364170 39250 364226
rect 39306 364170 39374 364226
rect 39430 364170 39498 364226
rect 39554 364170 39622 364226
rect 39678 364170 57250 364226
rect 57306 364170 57374 364226
rect 57430 364170 57498 364226
rect 57554 364170 57622 364226
rect 57678 364170 75250 364226
rect 75306 364170 75374 364226
rect 75430 364170 75498 364226
rect 75554 364170 75622 364226
rect 75678 364170 93250 364226
rect 93306 364170 93374 364226
rect 93430 364170 93498 364226
rect 93554 364170 93622 364226
rect 93678 364170 111250 364226
rect 111306 364170 111374 364226
rect 111430 364170 111498 364226
rect 111554 364170 111622 364226
rect 111678 364170 129250 364226
rect 129306 364170 129374 364226
rect 129430 364170 129498 364226
rect 129554 364170 129622 364226
rect 129678 364170 147250 364226
rect 147306 364170 147374 364226
rect 147430 364170 147498 364226
rect 147554 364170 147622 364226
rect 147678 364170 165250 364226
rect 165306 364170 165374 364226
rect 165430 364170 165498 364226
rect 165554 364170 165622 364226
rect 165678 364170 183250 364226
rect 183306 364170 183374 364226
rect 183430 364170 183498 364226
rect 183554 364170 183622 364226
rect 183678 364170 201250 364226
rect 201306 364170 201374 364226
rect 201430 364170 201498 364226
rect 201554 364170 201622 364226
rect 201678 364170 204518 364226
rect 204574 364170 204642 364226
rect 204698 364170 235238 364226
rect 235294 364170 235362 364226
rect 235418 364170 265958 364226
rect 266014 364170 266082 364226
rect 266138 364170 296678 364226
rect 296734 364170 296802 364226
rect 296858 364170 327398 364226
rect 327454 364170 327522 364226
rect 327578 364170 358118 364226
rect 358174 364170 358242 364226
rect 358298 364170 388838 364226
rect 388894 364170 388962 364226
rect 389018 364170 419558 364226
rect 419614 364170 419682 364226
rect 419738 364170 450278 364226
rect 450334 364170 450402 364226
rect 450458 364170 480998 364226
rect 481054 364170 481122 364226
rect 481178 364170 507250 364226
rect 507306 364170 507374 364226
rect 507430 364170 507498 364226
rect 507554 364170 507622 364226
rect 507678 364170 525250 364226
rect 525306 364170 525374 364226
rect 525430 364170 525498 364226
rect 525554 364170 525622 364226
rect 525678 364170 543250 364226
rect 543306 364170 543374 364226
rect 543430 364170 543498 364226
rect 543554 364170 543622 364226
rect 543678 364170 561250 364226
rect 561306 364170 561374 364226
rect 561430 364170 561498 364226
rect 561554 364170 561622 364226
rect 561678 364170 579250 364226
rect 579306 364170 579374 364226
rect 579430 364170 579498 364226
rect 579554 364170 579622 364226
rect 579678 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 3250 364102
rect 3306 364046 3374 364102
rect 3430 364046 3498 364102
rect 3554 364046 3622 364102
rect 3678 364046 21250 364102
rect 21306 364046 21374 364102
rect 21430 364046 21498 364102
rect 21554 364046 21622 364102
rect 21678 364046 39250 364102
rect 39306 364046 39374 364102
rect 39430 364046 39498 364102
rect 39554 364046 39622 364102
rect 39678 364046 57250 364102
rect 57306 364046 57374 364102
rect 57430 364046 57498 364102
rect 57554 364046 57622 364102
rect 57678 364046 75250 364102
rect 75306 364046 75374 364102
rect 75430 364046 75498 364102
rect 75554 364046 75622 364102
rect 75678 364046 93250 364102
rect 93306 364046 93374 364102
rect 93430 364046 93498 364102
rect 93554 364046 93622 364102
rect 93678 364046 111250 364102
rect 111306 364046 111374 364102
rect 111430 364046 111498 364102
rect 111554 364046 111622 364102
rect 111678 364046 129250 364102
rect 129306 364046 129374 364102
rect 129430 364046 129498 364102
rect 129554 364046 129622 364102
rect 129678 364046 147250 364102
rect 147306 364046 147374 364102
rect 147430 364046 147498 364102
rect 147554 364046 147622 364102
rect 147678 364046 165250 364102
rect 165306 364046 165374 364102
rect 165430 364046 165498 364102
rect 165554 364046 165622 364102
rect 165678 364046 183250 364102
rect 183306 364046 183374 364102
rect 183430 364046 183498 364102
rect 183554 364046 183622 364102
rect 183678 364046 201250 364102
rect 201306 364046 201374 364102
rect 201430 364046 201498 364102
rect 201554 364046 201622 364102
rect 201678 364046 204518 364102
rect 204574 364046 204642 364102
rect 204698 364046 235238 364102
rect 235294 364046 235362 364102
rect 235418 364046 265958 364102
rect 266014 364046 266082 364102
rect 266138 364046 296678 364102
rect 296734 364046 296802 364102
rect 296858 364046 327398 364102
rect 327454 364046 327522 364102
rect 327578 364046 358118 364102
rect 358174 364046 358242 364102
rect 358298 364046 388838 364102
rect 388894 364046 388962 364102
rect 389018 364046 419558 364102
rect 419614 364046 419682 364102
rect 419738 364046 450278 364102
rect 450334 364046 450402 364102
rect 450458 364046 480998 364102
rect 481054 364046 481122 364102
rect 481178 364046 507250 364102
rect 507306 364046 507374 364102
rect 507430 364046 507498 364102
rect 507554 364046 507622 364102
rect 507678 364046 525250 364102
rect 525306 364046 525374 364102
rect 525430 364046 525498 364102
rect 525554 364046 525622 364102
rect 525678 364046 543250 364102
rect 543306 364046 543374 364102
rect 543430 364046 543498 364102
rect 543554 364046 543622 364102
rect 543678 364046 561250 364102
rect 561306 364046 561374 364102
rect 561430 364046 561498 364102
rect 561554 364046 561622 364102
rect 561678 364046 579250 364102
rect 579306 364046 579374 364102
rect 579430 364046 579498 364102
rect 579554 364046 579622 364102
rect 579678 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 3250 363978
rect 3306 363922 3374 363978
rect 3430 363922 3498 363978
rect 3554 363922 3622 363978
rect 3678 363922 21250 363978
rect 21306 363922 21374 363978
rect 21430 363922 21498 363978
rect 21554 363922 21622 363978
rect 21678 363922 39250 363978
rect 39306 363922 39374 363978
rect 39430 363922 39498 363978
rect 39554 363922 39622 363978
rect 39678 363922 57250 363978
rect 57306 363922 57374 363978
rect 57430 363922 57498 363978
rect 57554 363922 57622 363978
rect 57678 363922 75250 363978
rect 75306 363922 75374 363978
rect 75430 363922 75498 363978
rect 75554 363922 75622 363978
rect 75678 363922 93250 363978
rect 93306 363922 93374 363978
rect 93430 363922 93498 363978
rect 93554 363922 93622 363978
rect 93678 363922 111250 363978
rect 111306 363922 111374 363978
rect 111430 363922 111498 363978
rect 111554 363922 111622 363978
rect 111678 363922 129250 363978
rect 129306 363922 129374 363978
rect 129430 363922 129498 363978
rect 129554 363922 129622 363978
rect 129678 363922 147250 363978
rect 147306 363922 147374 363978
rect 147430 363922 147498 363978
rect 147554 363922 147622 363978
rect 147678 363922 165250 363978
rect 165306 363922 165374 363978
rect 165430 363922 165498 363978
rect 165554 363922 165622 363978
rect 165678 363922 183250 363978
rect 183306 363922 183374 363978
rect 183430 363922 183498 363978
rect 183554 363922 183622 363978
rect 183678 363922 201250 363978
rect 201306 363922 201374 363978
rect 201430 363922 201498 363978
rect 201554 363922 201622 363978
rect 201678 363922 204518 363978
rect 204574 363922 204642 363978
rect 204698 363922 235238 363978
rect 235294 363922 235362 363978
rect 235418 363922 265958 363978
rect 266014 363922 266082 363978
rect 266138 363922 296678 363978
rect 296734 363922 296802 363978
rect 296858 363922 327398 363978
rect 327454 363922 327522 363978
rect 327578 363922 358118 363978
rect 358174 363922 358242 363978
rect 358298 363922 388838 363978
rect 388894 363922 388962 363978
rect 389018 363922 419558 363978
rect 419614 363922 419682 363978
rect 419738 363922 450278 363978
rect 450334 363922 450402 363978
rect 450458 363922 480998 363978
rect 481054 363922 481122 363978
rect 481178 363922 507250 363978
rect 507306 363922 507374 363978
rect 507430 363922 507498 363978
rect 507554 363922 507622 363978
rect 507678 363922 525250 363978
rect 525306 363922 525374 363978
rect 525430 363922 525498 363978
rect 525554 363922 525622 363978
rect 525678 363922 543250 363978
rect 543306 363922 543374 363978
rect 543430 363922 543498 363978
rect 543554 363922 543622 363978
rect 543678 363922 561250 363978
rect 561306 363922 561374 363978
rect 561430 363922 561498 363978
rect 561554 363922 561622 363978
rect 561678 363922 579250 363978
rect 579306 363922 579374 363978
rect 579430 363922 579498 363978
rect 579554 363922 579622 363978
rect 579678 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 6970 352350
rect 7026 352294 7094 352350
rect 7150 352294 7218 352350
rect 7274 352294 7342 352350
rect 7398 352294 24970 352350
rect 25026 352294 25094 352350
rect 25150 352294 25218 352350
rect 25274 352294 25342 352350
rect 25398 352294 42970 352350
rect 43026 352294 43094 352350
rect 43150 352294 43218 352350
rect 43274 352294 43342 352350
rect 43398 352294 60970 352350
rect 61026 352294 61094 352350
rect 61150 352294 61218 352350
rect 61274 352294 61342 352350
rect 61398 352294 78970 352350
rect 79026 352294 79094 352350
rect 79150 352294 79218 352350
rect 79274 352294 79342 352350
rect 79398 352294 96970 352350
rect 97026 352294 97094 352350
rect 97150 352294 97218 352350
rect 97274 352294 97342 352350
rect 97398 352294 114970 352350
rect 115026 352294 115094 352350
rect 115150 352294 115218 352350
rect 115274 352294 115342 352350
rect 115398 352294 132970 352350
rect 133026 352294 133094 352350
rect 133150 352294 133218 352350
rect 133274 352294 133342 352350
rect 133398 352294 150970 352350
rect 151026 352294 151094 352350
rect 151150 352294 151218 352350
rect 151274 352294 151342 352350
rect 151398 352294 168970 352350
rect 169026 352294 169094 352350
rect 169150 352294 169218 352350
rect 169274 352294 169342 352350
rect 169398 352294 186970 352350
rect 187026 352294 187094 352350
rect 187150 352294 187218 352350
rect 187274 352294 187342 352350
rect 187398 352294 219878 352350
rect 219934 352294 220002 352350
rect 220058 352294 250598 352350
rect 250654 352294 250722 352350
rect 250778 352294 281318 352350
rect 281374 352294 281442 352350
rect 281498 352294 312038 352350
rect 312094 352294 312162 352350
rect 312218 352294 342758 352350
rect 342814 352294 342882 352350
rect 342938 352294 373478 352350
rect 373534 352294 373602 352350
rect 373658 352294 404198 352350
rect 404254 352294 404322 352350
rect 404378 352294 434918 352350
rect 434974 352294 435042 352350
rect 435098 352294 465638 352350
rect 465694 352294 465762 352350
rect 465818 352294 496358 352350
rect 496414 352294 496482 352350
rect 496538 352294 510970 352350
rect 511026 352294 511094 352350
rect 511150 352294 511218 352350
rect 511274 352294 511342 352350
rect 511398 352294 528970 352350
rect 529026 352294 529094 352350
rect 529150 352294 529218 352350
rect 529274 352294 529342 352350
rect 529398 352294 546970 352350
rect 547026 352294 547094 352350
rect 547150 352294 547218 352350
rect 547274 352294 547342 352350
rect 547398 352294 564970 352350
rect 565026 352294 565094 352350
rect 565150 352294 565218 352350
rect 565274 352294 565342 352350
rect 565398 352294 582970 352350
rect 583026 352294 583094 352350
rect 583150 352294 583218 352350
rect 583274 352294 583342 352350
rect 583398 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 6970 352226
rect 7026 352170 7094 352226
rect 7150 352170 7218 352226
rect 7274 352170 7342 352226
rect 7398 352170 24970 352226
rect 25026 352170 25094 352226
rect 25150 352170 25218 352226
rect 25274 352170 25342 352226
rect 25398 352170 42970 352226
rect 43026 352170 43094 352226
rect 43150 352170 43218 352226
rect 43274 352170 43342 352226
rect 43398 352170 60970 352226
rect 61026 352170 61094 352226
rect 61150 352170 61218 352226
rect 61274 352170 61342 352226
rect 61398 352170 78970 352226
rect 79026 352170 79094 352226
rect 79150 352170 79218 352226
rect 79274 352170 79342 352226
rect 79398 352170 96970 352226
rect 97026 352170 97094 352226
rect 97150 352170 97218 352226
rect 97274 352170 97342 352226
rect 97398 352170 114970 352226
rect 115026 352170 115094 352226
rect 115150 352170 115218 352226
rect 115274 352170 115342 352226
rect 115398 352170 132970 352226
rect 133026 352170 133094 352226
rect 133150 352170 133218 352226
rect 133274 352170 133342 352226
rect 133398 352170 150970 352226
rect 151026 352170 151094 352226
rect 151150 352170 151218 352226
rect 151274 352170 151342 352226
rect 151398 352170 168970 352226
rect 169026 352170 169094 352226
rect 169150 352170 169218 352226
rect 169274 352170 169342 352226
rect 169398 352170 186970 352226
rect 187026 352170 187094 352226
rect 187150 352170 187218 352226
rect 187274 352170 187342 352226
rect 187398 352170 219878 352226
rect 219934 352170 220002 352226
rect 220058 352170 250598 352226
rect 250654 352170 250722 352226
rect 250778 352170 281318 352226
rect 281374 352170 281442 352226
rect 281498 352170 312038 352226
rect 312094 352170 312162 352226
rect 312218 352170 342758 352226
rect 342814 352170 342882 352226
rect 342938 352170 373478 352226
rect 373534 352170 373602 352226
rect 373658 352170 404198 352226
rect 404254 352170 404322 352226
rect 404378 352170 434918 352226
rect 434974 352170 435042 352226
rect 435098 352170 465638 352226
rect 465694 352170 465762 352226
rect 465818 352170 496358 352226
rect 496414 352170 496482 352226
rect 496538 352170 510970 352226
rect 511026 352170 511094 352226
rect 511150 352170 511218 352226
rect 511274 352170 511342 352226
rect 511398 352170 528970 352226
rect 529026 352170 529094 352226
rect 529150 352170 529218 352226
rect 529274 352170 529342 352226
rect 529398 352170 546970 352226
rect 547026 352170 547094 352226
rect 547150 352170 547218 352226
rect 547274 352170 547342 352226
rect 547398 352170 564970 352226
rect 565026 352170 565094 352226
rect 565150 352170 565218 352226
rect 565274 352170 565342 352226
rect 565398 352170 582970 352226
rect 583026 352170 583094 352226
rect 583150 352170 583218 352226
rect 583274 352170 583342 352226
rect 583398 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 6970 352102
rect 7026 352046 7094 352102
rect 7150 352046 7218 352102
rect 7274 352046 7342 352102
rect 7398 352046 24970 352102
rect 25026 352046 25094 352102
rect 25150 352046 25218 352102
rect 25274 352046 25342 352102
rect 25398 352046 42970 352102
rect 43026 352046 43094 352102
rect 43150 352046 43218 352102
rect 43274 352046 43342 352102
rect 43398 352046 60970 352102
rect 61026 352046 61094 352102
rect 61150 352046 61218 352102
rect 61274 352046 61342 352102
rect 61398 352046 78970 352102
rect 79026 352046 79094 352102
rect 79150 352046 79218 352102
rect 79274 352046 79342 352102
rect 79398 352046 96970 352102
rect 97026 352046 97094 352102
rect 97150 352046 97218 352102
rect 97274 352046 97342 352102
rect 97398 352046 114970 352102
rect 115026 352046 115094 352102
rect 115150 352046 115218 352102
rect 115274 352046 115342 352102
rect 115398 352046 132970 352102
rect 133026 352046 133094 352102
rect 133150 352046 133218 352102
rect 133274 352046 133342 352102
rect 133398 352046 150970 352102
rect 151026 352046 151094 352102
rect 151150 352046 151218 352102
rect 151274 352046 151342 352102
rect 151398 352046 168970 352102
rect 169026 352046 169094 352102
rect 169150 352046 169218 352102
rect 169274 352046 169342 352102
rect 169398 352046 186970 352102
rect 187026 352046 187094 352102
rect 187150 352046 187218 352102
rect 187274 352046 187342 352102
rect 187398 352046 219878 352102
rect 219934 352046 220002 352102
rect 220058 352046 250598 352102
rect 250654 352046 250722 352102
rect 250778 352046 281318 352102
rect 281374 352046 281442 352102
rect 281498 352046 312038 352102
rect 312094 352046 312162 352102
rect 312218 352046 342758 352102
rect 342814 352046 342882 352102
rect 342938 352046 373478 352102
rect 373534 352046 373602 352102
rect 373658 352046 404198 352102
rect 404254 352046 404322 352102
rect 404378 352046 434918 352102
rect 434974 352046 435042 352102
rect 435098 352046 465638 352102
rect 465694 352046 465762 352102
rect 465818 352046 496358 352102
rect 496414 352046 496482 352102
rect 496538 352046 510970 352102
rect 511026 352046 511094 352102
rect 511150 352046 511218 352102
rect 511274 352046 511342 352102
rect 511398 352046 528970 352102
rect 529026 352046 529094 352102
rect 529150 352046 529218 352102
rect 529274 352046 529342 352102
rect 529398 352046 546970 352102
rect 547026 352046 547094 352102
rect 547150 352046 547218 352102
rect 547274 352046 547342 352102
rect 547398 352046 564970 352102
rect 565026 352046 565094 352102
rect 565150 352046 565218 352102
rect 565274 352046 565342 352102
rect 565398 352046 582970 352102
rect 583026 352046 583094 352102
rect 583150 352046 583218 352102
rect 583274 352046 583342 352102
rect 583398 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 6970 351978
rect 7026 351922 7094 351978
rect 7150 351922 7218 351978
rect 7274 351922 7342 351978
rect 7398 351922 24970 351978
rect 25026 351922 25094 351978
rect 25150 351922 25218 351978
rect 25274 351922 25342 351978
rect 25398 351922 42970 351978
rect 43026 351922 43094 351978
rect 43150 351922 43218 351978
rect 43274 351922 43342 351978
rect 43398 351922 60970 351978
rect 61026 351922 61094 351978
rect 61150 351922 61218 351978
rect 61274 351922 61342 351978
rect 61398 351922 78970 351978
rect 79026 351922 79094 351978
rect 79150 351922 79218 351978
rect 79274 351922 79342 351978
rect 79398 351922 96970 351978
rect 97026 351922 97094 351978
rect 97150 351922 97218 351978
rect 97274 351922 97342 351978
rect 97398 351922 114970 351978
rect 115026 351922 115094 351978
rect 115150 351922 115218 351978
rect 115274 351922 115342 351978
rect 115398 351922 132970 351978
rect 133026 351922 133094 351978
rect 133150 351922 133218 351978
rect 133274 351922 133342 351978
rect 133398 351922 150970 351978
rect 151026 351922 151094 351978
rect 151150 351922 151218 351978
rect 151274 351922 151342 351978
rect 151398 351922 168970 351978
rect 169026 351922 169094 351978
rect 169150 351922 169218 351978
rect 169274 351922 169342 351978
rect 169398 351922 186970 351978
rect 187026 351922 187094 351978
rect 187150 351922 187218 351978
rect 187274 351922 187342 351978
rect 187398 351922 219878 351978
rect 219934 351922 220002 351978
rect 220058 351922 250598 351978
rect 250654 351922 250722 351978
rect 250778 351922 281318 351978
rect 281374 351922 281442 351978
rect 281498 351922 312038 351978
rect 312094 351922 312162 351978
rect 312218 351922 342758 351978
rect 342814 351922 342882 351978
rect 342938 351922 373478 351978
rect 373534 351922 373602 351978
rect 373658 351922 404198 351978
rect 404254 351922 404322 351978
rect 404378 351922 434918 351978
rect 434974 351922 435042 351978
rect 435098 351922 465638 351978
rect 465694 351922 465762 351978
rect 465818 351922 496358 351978
rect 496414 351922 496482 351978
rect 496538 351922 510970 351978
rect 511026 351922 511094 351978
rect 511150 351922 511218 351978
rect 511274 351922 511342 351978
rect 511398 351922 528970 351978
rect 529026 351922 529094 351978
rect 529150 351922 529218 351978
rect 529274 351922 529342 351978
rect 529398 351922 546970 351978
rect 547026 351922 547094 351978
rect 547150 351922 547218 351978
rect 547274 351922 547342 351978
rect 547398 351922 564970 351978
rect 565026 351922 565094 351978
rect 565150 351922 565218 351978
rect 565274 351922 565342 351978
rect 565398 351922 582970 351978
rect 583026 351922 583094 351978
rect 583150 351922 583218 351978
rect 583274 351922 583342 351978
rect 583398 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 3250 346350
rect 3306 346294 3374 346350
rect 3430 346294 3498 346350
rect 3554 346294 3622 346350
rect 3678 346294 21250 346350
rect 21306 346294 21374 346350
rect 21430 346294 21498 346350
rect 21554 346294 21622 346350
rect 21678 346294 39250 346350
rect 39306 346294 39374 346350
rect 39430 346294 39498 346350
rect 39554 346294 39622 346350
rect 39678 346294 57250 346350
rect 57306 346294 57374 346350
rect 57430 346294 57498 346350
rect 57554 346294 57622 346350
rect 57678 346294 75250 346350
rect 75306 346294 75374 346350
rect 75430 346294 75498 346350
rect 75554 346294 75622 346350
rect 75678 346294 93250 346350
rect 93306 346294 93374 346350
rect 93430 346294 93498 346350
rect 93554 346294 93622 346350
rect 93678 346294 111250 346350
rect 111306 346294 111374 346350
rect 111430 346294 111498 346350
rect 111554 346294 111622 346350
rect 111678 346294 129250 346350
rect 129306 346294 129374 346350
rect 129430 346294 129498 346350
rect 129554 346294 129622 346350
rect 129678 346294 147250 346350
rect 147306 346294 147374 346350
rect 147430 346294 147498 346350
rect 147554 346294 147622 346350
rect 147678 346294 165250 346350
rect 165306 346294 165374 346350
rect 165430 346294 165498 346350
rect 165554 346294 165622 346350
rect 165678 346294 183250 346350
rect 183306 346294 183374 346350
rect 183430 346294 183498 346350
rect 183554 346294 183622 346350
rect 183678 346294 201250 346350
rect 201306 346294 201374 346350
rect 201430 346294 201498 346350
rect 201554 346294 201622 346350
rect 201678 346294 204518 346350
rect 204574 346294 204642 346350
rect 204698 346294 235238 346350
rect 235294 346294 235362 346350
rect 235418 346294 265958 346350
rect 266014 346294 266082 346350
rect 266138 346294 296678 346350
rect 296734 346294 296802 346350
rect 296858 346294 327398 346350
rect 327454 346294 327522 346350
rect 327578 346294 358118 346350
rect 358174 346294 358242 346350
rect 358298 346294 388838 346350
rect 388894 346294 388962 346350
rect 389018 346294 419558 346350
rect 419614 346294 419682 346350
rect 419738 346294 450278 346350
rect 450334 346294 450402 346350
rect 450458 346294 480998 346350
rect 481054 346294 481122 346350
rect 481178 346294 507250 346350
rect 507306 346294 507374 346350
rect 507430 346294 507498 346350
rect 507554 346294 507622 346350
rect 507678 346294 525250 346350
rect 525306 346294 525374 346350
rect 525430 346294 525498 346350
rect 525554 346294 525622 346350
rect 525678 346294 543250 346350
rect 543306 346294 543374 346350
rect 543430 346294 543498 346350
rect 543554 346294 543622 346350
rect 543678 346294 561250 346350
rect 561306 346294 561374 346350
rect 561430 346294 561498 346350
rect 561554 346294 561622 346350
rect 561678 346294 579250 346350
rect 579306 346294 579374 346350
rect 579430 346294 579498 346350
rect 579554 346294 579622 346350
rect 579678 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 3250 346226
rect 3306 346170 3374 346226
rect 3430 346170 3498 346226
rect 3554 346170 3622 346226
rect 3678 346170 21250 346226
rect 21306 346170 21374 346226
rect 21430 346170 21498 346226
rect 21554 346170 21622 346226
rect 21678 346170 39250 346226
rect 39306 346170 39374 346226
rect 39430 346170 39498 346226
rect 39554 346170 39622 346226
rect 39678 346170 57250 346226
rect 57306 346170 57374 346226
rect 57430 346170 57498 346226
rect 57554 346170 57622 346226
rect 57678 346170 75250 346226
rect 75306 346170 75374 346226
rect 75430 346170 75498 346226
rect 75554 346170 75622 346226
rect 75678 346170 93250 346226
rect 93306 346170 93374 346226
rect 93430 346170 93498 346226
rect 93554 346170 93622 346226
rect 93678 346170 111250 346226
rect 111306 346170 111374 346226
rect 111430 346170 111498 346226
rect 111554 346170 111622 346226
rect 111678 346170 129250 346226
rect 129306 346170 129374 346226
rect 129430 346170 129498 346226
rect 129554 346170 129622 346226
rect 129678 346170 147250 346226
rect 147306 346170 147374 346226
rect 147430 346170 147498 346226
rect 147554 346170 147622 346226
rect 147678 346170 165250 346226
rect 165306 346170 165374 346226
rect 165430 346170 165498 346226
rect 165554 346170 165622 346226
rect 165678 346170 183250 346226
rect 183306 346170 183374 346226
rect 183430 346170 183498 346226
rect 183554 346170 183622 346226
rect 183678 346170 201250 346226
rect 201306 346170 201374 346226
rect 201430 346170 201498 346226
rect 201554 346170 201622 346226
rect 201678 346170 204518 346226
rect 204574 346170 204642 346226
rect 204698 346170 235238 346226
rect 235294 346170 235362 346226
rect 235418 346170 265958 346226
rect 266014 346170 266082 346226
rect 266138 346170 296678 346226
rect 296734 346170 296802 346226
rect 296858 346170 327398 346226
rect 327454 346170 327522 346226
rect 327578 346170 358118 346226
rect 358174 346170 358242 346226
rect 358298 346170 388838 346226
rect 388894 346170 388962 346226
rect 389018 346170 419558 346226
rect 419614 346170 419682 346226
rect 419738 346170 450278 346226
rect 450334 346170 450402 346226
rect 450458 346170 480998 346226
rect 481054 346170 481122 346226
rect 481178 346170 507250 346226
rect 507306 346170 507374 346226
rect 507430 346170 507498 346226
rect 507554 346170 507622 346226
rect 507678 346170 525250 346226
rect 525306 346170 525374 346226
rect 525430 346170 525498 346226
rect 525554 346170 525622 346226
rect 525678 346170 543250 346226
rect 543306 346170 543374 346226
rect 543430 346170 543498 346226
rect 543554 346170 543622 346226
rect 543678 346170 561250 346226
rect 561306 346170 561374 346226
rect 561430 346170 561498 346226
rect 561554 346170 561622 346226
rect 561678 346170 579250 346226
rect 579306 346170 579374 346226
rect 579430 346170 579498 346226
rect 579554 346170 579622 346226
rect 579678 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 3250 346102
rect 3306 346046 3374 346102
rect 3430 346046 3498 346102
rect 3554 346046 3622 346102
rect 3678 346046 21250 346102
rect 21306 346046 21374 346102
rect 21430 346046 21498 346102
rect 21554 346046 21622 346102
rect 21678 346046 39250 346102
rect 39306 346046 39374 346102
rect 39430 346046 39498 346102
rect 39554 346046 39622 346102
rect 39678 346046 57250 346102
rect 57306 346046 57374 346102
rect 57430 346046 57498 346102
rect 57554 346046 57622 346102
rect 57678 346046 75250 346102
rect 75306 346046 75374 346102
rect 75430 346046 75498 346102
rect 75554 346046 75622 346102
rect 75678 346046 93250 346102
rect 93306 346046 93374 346102
rect 93430 346046 93498 346102
rect 93554 346046 93622 346102
rect 93678 346046 111250 346102
rect 111306 346046 111374 346102
rect 111430 346046 111498 346102
rect 111554 346046 111622 346102
rect 111678 346046 129250 346102
rect 129306 346046 129374 346102
rect 129430 346046 129498 346102
rect 129554 346046 129622 346102
rect 129678 346046 147250 346102
rect 147306 346046 147374 346102
rect 147430 346046 147498 346102
rect 147554 346046 147622 346102
rect 147678 346046 165250 346102
rect 165306 346046 165374 346102
rect 165430 346046 165498 346102
rect 165554 346046 165622 346102
rect 165678 346046 183250 346102
rect 183306 346046 183374 346102
rect 183430 346046 183498 346102
rect 183554 346046 183622 346102
rect 183678 346046 201250 346102
rect 201306 346046 201374 346102
rect 201430 346046 201498 346102
rect 201554 346046 201622 346102
rect 201678 346046 204518 346102
rect 204574 346046 204642 346102
rect 204698 346046 235238 346102
rect 235294 346046 235362 346102
rect 235418 346046 265958 346102
rect 266014 346046 266082 346102
rect 266138 346046 296678 346102
rect 296734 346046 296802 346102
rect 296858 346046 327398 346102
rect 327454 346046 327522 346102
rect 327578 346046 358118 346102
rect 358174 346046 358242 346102
rect 358298 346046 388838 346102
rect 388894 346046 388962 346102
rect 389018 346046 419558 346102
rect 419614 346046 419682 346102
rect 419738 346046 450278 346102
rect 450334 346046 450402 346102
rect 450458 346046 480998 346102
rect 481054 346046 481122 346102
rect 481178 346046 507250 346102
rect 507306 346046 507374 346102
rect 507430 346046 507498 346102
rect 507554 346046 507622 346102
rect 507678 346046 525250 346102
rect 525306 346046 525374 346102
rect 525430 346046 525498 346102
rect 525554 346046 525622 346102
rect 525678 346046 543250 346102
rect 543306 346046 543374 346102
rect 543430 346046 543498 346102
rect 543554 346046 543622 346102
rect 543678 346046 561250 346102
rect 561306 346046 561374 346102
rect 561430 346046 561498 346102
rect 561554 346046 561622 346102
rect 561678 346046 579250 346102
rect 579306 346046 579374 346102
rect 579430 346046 579498 346102
rect 579554 346046 579622 346102
rect 579678 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 3250 345978
rect 3306 345922 3374 345978
rect 3430 345922 3498 345978
rect 3554 345922 3622 345978
rect 3678 345922 21250 345978
rect 21306 345922 21374 345978
rect 21430 345922 21498 345978
rect 21554 345922 21622 345978
rect 21678 345922 39250 345978
rect 39306 345922 39374 345978
rect 39430 345922 39498 345978
rect 39554 345922 39622 345978
rect 39678 345922 57250 345978
rect 57306 345922 57374 345978
rect 57430 345922 57498 345978
rect 57554 345922 57622 345978
rect 57678 345922 75250 345978
rect 75306 345922 75374 345978
rect 75430 345922 75498 345978
rect 75554 345922 75622 345978
rect 75678 345922 93250 345978
rect 93306 345922 93374 345978
rect 93430 345922 93498 345978
rect 93554 345922 93622 345978
rect 93678 345922 111250 345978
rect 111306 345922 111374 345978
rect 111430 345922 111498 345978
rect 111554 345922 111622 345978
rect 111678 345922 129250 345978
rect 129306 345922 129374 345978
rect 129430 345922 129498 345978
rect 129554 345922 129622 345978
rect 129678 345922 147250 345978
rect 147306 345922 147374 345978
rect 147430 345922 147498 345978
rect 147554 345922 147622 345978
rect 147678 345922 165250 345978
rect 165306 345922 165374 345978
rect 165430 345922 165498 345978
rect 165554 345922 165622 345978
rect 165678 345922 183250 345978
rect 183306 345922 183374 345978
rect 183430 345922 183498 345978
rect 183554 345922 183622 345978
rect 183678 345922 201250 345978
rect 201306 345922 201374 345978
rect 201430 345922 201498 345978
rect 201554 345922 201622 345978
rect 201678 345922 204518 345978
rect 204574 345922 204642 345978
rect 204698 345922 235238 345978
rect 235294 345922 235362 345978
rect 235418 345922 265958 345978
rect 266014 345922 266082 345978
rect 266138 345922 296678 345978
rect 296734 345922 296802 345978
rect 296858 345922 327398 345978
rect 327454 345922 327522 345978
rect 327578 345922 358118 345978
rect 358174 345922 358242 345978
rect 358298 345922 388838 345978
rect 388894 345922 388962 345978
rect 389018 345922 419558 345978
rect 419614 345922 419682 345978
rect 419738 345922 450278 345978
rect 450334 345922 450402 345978
rect 450458 345922 480998 345978
rect 481054 345922 481122 345978
rect 481178 345922 507250 345978
rect 507306 345922 507374 345978
rect 507430 345922 507498 345978
rect 507554 345922 507622 345978
rect 507678 345922 525250 345978
rect 525306 345922 525374 345978
rect 525430 345922 525498 345978
rect 525554 345922 525622 345978
rect 525678 345922 543250 345978
rect 543306 345922 543374 345978
rect 543430 345922 543498 345978
rect 543554 345922 543622 345978
rect 543678 345922 561250 345978
rect 561306 345922 561374 345978
rect 561430 345922 561498 345978
rect 561554 345922 561622 345978
rect 561678 345922 579250 345978
rect 579306 345922 579374 345978
rect 579430 345922 579498 345978
rect 579554 345922 579622 345978
rect 579678 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 6970 334350
rect 7026 334294 7094 334350
rect 7150 334294 7218 334350
rect 7274 334294 7342 334350
rect 7398 334294 24970 334350
rect 25026 334294 25094 334350
rect 25150 334294 25218 334350
rect 25274 334294 25342 334350
rect 25398 334294 42970 334350
rect 43026 334294 43094 334350
rect 43150 334294 43218 334350
rect 43274 334294 43342 334350
rect 43398 334294 60970 334350
rect 61026 334294 61094 334350
rect 61150 334294 61218 334350
rect 61274 334294 61342 334350
rect 61398 334294 78970 334350
rect 79026 334294 79094 334350
rect 79150 334294 79218 334350
rect 79274 334294 79342 334350
rect 79398 334294 96970 334350
rect 97026 334294 97094 334350
rect 97150 334294 97218 334350
rect 97274 334294 97342 334350
rect 97398 334294 114970 334350
rect 115026 334294 115094 334350
rect 115150 334294 115218 334350
rect 115274 334294 115342 334350
rect 115398 334294 132970 334350
rect 133026 334294 133094 334350
rect 133150 334294 133218 334350
rect 133274 334294 133342 334350
rect 133398 334294 150970 334350
rect 151026 334294 151094 334350
rect 151150 334294 151218 334350
rect 151274 334294 151342 334350
rect 151398 334294 168970 334350
rect 169026 334294 169094 334350
rect 169150 334294 169218 334350
rect 169274 334294 169342 334350
rect 169398 334294 186970 334350
rect 187026 334294 187094 334350
rect 187150 334294 187218 334350
rect 187274 334294 187342 334350
rect 187398 334294 219878 334350
rect 219934 334294 220002 334350
rect 220058 334294 250598 334350
rect 250654 334294 250722 334350
rect 250778 334294 281318 334350
rect 281374 334294 281442 334350
rect 281498 334294 312038 334350
rect 312094 334294 312162 334350
rect 312218 334294 342758 334350
rect 342814 334294 342882 334350
rect 342938 334294 373478 334350
rect 373534 334294 373602 334350
rect 373658 334294 404198 334350
rect 404254 334294 404322 334350
rect 404378 334294 434918 334350
rect 434974 334294 435042 334350
rect 435098 334294 465638 334350
rect 465694 334294 465762 334350
rect 465818 334294 496358 334350
rect 496414 334294 496482 334350
rect 496538 334294 510970 334350
rect 511026 334294 511094 334350
rect 511150 334294 511218 334350
rect 511274 334294 511342 334350
rect 511398 334294 528970 334350
rect 529026 334294 529094 334350
rect 529150 334294 529218 334350
rect 529274 334294 529342 334350
rect 529398 334294 546970 334350
rect 547026 334294 547094 334350
rect 547150 334294 547218 334350
rect 547274 334294 547342 334350
rect 547398 334294 564970 334350
rect 565026 334294 565094 334350
rect 565150 334294 565218 334350
rect 565274 334294 565342 334350
rect 565398 334294 582970 334350
rect 583026 334294 583094 334350
rect 583150 334294 583218 334350
rect 583274 334294 583342 334350
rect 583398 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 6970 334226
rect 7026 334170 7094 334226
rect 7150 334170 7218 334226
rect 7274 334170 7342 334226
rect 7398 334170 24970 334226
rect 25026 334170 25094 334226
rect 25150 334170 25218 334226
rect 25274 334170 25342 334226
rect 25398 334170 42970 334226
rect 43026 334170 43094 334226
rect 43150 334170 43218 334226
rect 43274 334170 43342 334226
rect 43398 334170 60970 334226
rect 61026 334170 61094 334226
rect 61150 334170 61218 334226
rect 61274 334170 61342 334226
rect 61398 334170 78970 334226
rect 79026 334170 79094 334226
rect 79150 334170 79218 334226
rect 79274 334170 79342 334226
rect 79398 334170 96970 334226
rect 97026 334170 97094 334226
rect 97150 334170 97218 334226
rect 97274 334170 97342 334226
rect 97398 334170 114970 334226
rect 115026 334170 115094 334226
rect 115150 334170 115218 334226
rect 115274 334170 115342 334226
rect 115398 334170 132970 334226
rect 133026 334170 133094 334226
rect 133150 334170 133218 334226
rect 133274 334170 133342 334226
rect 133398 334170 150970 334226
rect 151026 334170 151094 334226
rect 151150 334170 151218 334226
rect 151274 334170 151342 334226
rect 151398 334170 168970 334226
rect 169026 334170 169094 334226
rect 169150 334170 169218 334226
rect 169274 334170 169342 334226
rect 169398 334170 186970 334226
rect 187026 334170 187094 334226
rect 187150 334170 187218 334226
rect 187274 334170 187342 334226
rect 187398 334170 219878 334226
rect 219934 334170 220002 334226
rect 220058 334170 250598 334226
rect 250654 334170 250722 334226
rect 250778 334170 281318 334226
rect 281374 334170 281442 334226
rect 281498 334170 312038 334226
rect 312094 334170 312162 334226
rect 312218 334170 342758 334226
rect 342814 334170 342882 334226
rect 342938 334170 373478 334226
rect 373534 334170 373602 334226
rect 373658 334170 404198 334226
rect 404254 334170 404322 334226
rect 404378 334170 434918 334226
rect 434974 334170 435042 334226
rect 435098 334170 465638 334226
rect 465694 334170 465762 334226
rect 465818 334170 496358 334226
rect 496414 334170 496482 334226
rect 496538 334170 510970 334226
rect 511026 334170 511094 334226
rect 511150 334170 511218 334226
rect 511274 334170 511342 334226
rect 511398 334170 528970 334226
rect 529026 334170 529094 334226
rect 529150 334170 529218 334226
rect 529274 334170 529342 334226
rect 529398 334170 546970 334226
rect 547026 334170 547094 334226
rect 547150 334170 547218 334226
rect 547274 334170 547342 334226
rect 547398 334170 564970 334226
rect 565026 334170 565094 334226
rect 565150 334170 565218 334226
rect 565274 334170 565342 334226
rect 565398 334170 582970 334226
rect 583026 334170 583094 334226
rect 583150 334170 583218 334226
rect 583274 334170 583342 334226
rect 583398 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 6970 334102
rect 7026 334046 7094 334102
rect 7150 334046 7218 334102
rect 7274 334046 7342 334102
rect 7398 334046 24970 334102
rect 25026 334046 25094 334102
rect 25150 334046 25218 334102
rect 25274 334046 25342 334102
rect 25398 334046 42970 334102
rect 43026 334046 43094 334102
rect 43150 334046 43218 334102
rect 43274 334046 43342 334102
rect 43398 334046 60970 334102
rect 61026 334046 61094 334102
rect 61150 334046 61218 334102
rect 61274 334046 61342 334102
rect 61398 334046 78970 334102
rect 79026 334046 79094 334102
rect 79150 334046 79218 334102
rect 79274 334046 79342 334102
rect 79398 334046 96970 334102
rect 97026 334046 97094 334102
rect 97150 334046 97218 334102
rect 97274 334046 97342 334102
rect 97398 334046 114970 334102
rect 115026 334046 115094 334102
rect 115150 334046 115218 334102
rect 115274 334046 115342 334102
rect 115398 334046 132970 334102
rect 133026 334046 133094 334102
rect 133150 334046 133218 334102
rect 133274 334046 133342 334102
rect 133398 334046 150970 334102
rect 151026 334046 151094 334102
rect 151150 334046 151218 334102
rect 151274 334046 151342 334102
rect 151398 334046 168970 334102
rect 169026 334046 169094 334102
rect 169150 334046 169218 334102
rect 169274 334046 169342 334102
rect 169398 334046 186970 334102
rect 187026 334046 187094 334102
rect 187150 334046 187218 334102
rect 187274 334046 187342 334102
rect 187398 334046 219878 334102
rect 219934 334046 220002 334102
rect 220058 334046 250598 334102
rect 250654 334046 250722 334102
rect 250778 334046 281318 334102
rect 281374 334046 281442 334102
rect 281498 334046 312038 334102
rect 312094 334046 312162 334102
rect 312218 334046 342758 334102
rect 342814 334046 342882 334102
rect 342938 334046 373478 334102
rect 373534 334046 373602 334102
rect 373658 334046 404198 334102
rect 404254 334046 404322 334102
rect 404378 334046 434918 334102
rect 434974 334046 435042 334102
rect 435098 334046 465638 334102
rect 465694 334046 465762 334102
rect 465818 334046 496358 334102
rect 496414 334046 496482 334102
rect 496538 334046 510970 334102
rect 511026 334046 511094 334102
rect 511150 334046 511218 334102
rect 511274 334046 511342 334102
rect 511398 334046 528970 334102
rect 529026 334046 529094 334102
rect 529150 334046 529218 334102
rect 529274 334046 529342 334102
rect 529398 334046 546970 334102
rect 547026 334046 547094 334102
rect 547150 334046 547218 334102
rect 547274 334046 547342 334102
rect 547398 334046 564970 334102
rect 565026 334046 565094 334102
rect 565150 334046 565218 334102
rect 565274 334046 565342 334102
rect 565398 334046 582970 334102
rect 583026 334046 583094 334102
rect 583150 334046 583218 334102
rect 583274 334046 583342 334102
rect 583398 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 6970 333978
rect 7026 333922 7094 333978
rect 7150 333922 7218 333978
rect 7274 333922 7342 333978
rect 7398 333922 24970 333978
rect 25026 333922 25094 333978
rect 25150 333922 25218 333978
rect 25274 333922 25342 333978
rect 25398 333922 42970 333978
rect 43026 333922 43094 333978
rect 43150 333922 43218 333978
rect 43274 333922 43342 333978
rect 43398 333922 60970 333978
rect 61026 333922 61094 333978
rect 61150 333922 61218 333978
rect 61274 333922 61342 333978
rect 61398 333922 78970 333978
rect 79026 333922 79094 333978
rect 79150 333922 79218 333978
rect 79274 333922 79342 333978
rect 79398 333922 96970 333978
rect 97026 333922 97094 333978
rect 97150 333922 97218 333978
rect 97274 333922 97342 333978
rect 97398 333922 114970 333978
rect 115026 333922 115094 333978
rect 115150 333922 115218 333978
rect 115274 333922 115342 333978
rect 115398 333922 132970 333978
rect 133026 333922 133094 333978
rect 133150 333922 133218 333978
rect 133274 333922 133342 333978
rect 133398 333922 150970 333978
rect 151026 333922 151094 333978
rect 151150 333922 151218 333978
rect 151274 333922 151342 333978
rect 151398 333922 168970 333978
rect 169026 333922 169094 333978
rect 169150 333922 169218 333978
rect 169274 333922 169342 333978
rect 169398 333922 186970 333978
rect 187026 333922 187094 333978
rect 187150 333922 187218 333978
rect 187274 333922 187342 333978
rect 187398 333922 219878 333978
rect 219934 333922 220002 333978
rect 220058 333922 250598 333978
rect 250654 333922 250722 333978
rect 250778 333922 281318 333978
rect 281374 333922 281442 333978
rect 281498 333922 312038 333978
rect 312094 333922 312162 333978
rect 312218 333922 342758 333978
rect 342814 333922 342882 333978
rect 342938 333922 373478 333978
rect 373534 333922 373602 333978
rect 373658 333922 404198 333978
rect 404254 333922 404322 333978
rect 404378 333922 434918 333978
rect 434974 333922 435042 333978
rect 435098 333922 465638 333978
rect 465694 333922 465762 333978
rect 465818 333922 496358 333978
rect 496414 333922 496482 333978
rect 496538 333922 510970 333978
rect 511026 333922 511094 333978
rect 511150 333922 511218 333978
rect 511274 333922 511342 333978
rect 511398 333922 528970 333978
rect 529026 333922 529094 333978
rect 529150 333922 529218 333978
rect 529274 333922 529342 333978
rect 529398 333922 546970 333978
rect 547026 333922 547094 333978
rect 547150 333922 547218 333978
rect 547274 333922 547342 333978
rect 547398 333922 564970 333978
rect 565026 333922 565094 333978
rect 565150 333922 565218 333978
rect 565274 333922 565342 333978
rect 565398 333922 582970 333978
rect 583026 333922 583094 333978
rect 583150 333922 583218 333978
rect 583274 333922 583342 333978
rect 583398 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 3250 328350
rect 3306 328294 3374 328350
rect 3430 328294 3498 328350
rect 3554 328294 3622 328350
rect 3678 328294 21250 328350
rect 21306 328294 21374 328350
rect 21430 328294 21498 328350
rect 21554 328294 21622 328350
rect 21678 328294 39250 328350
rect 39306 328294 39374 328350
rect 39430 328294 39498 328350
rect 39554 328294 39622 328350
rect 39678 328294 57250 328350
rect 57306 328294 57374 328350
rect 57430 328294 57498 328350
rect 57554 328294 57622 328350
rect 57678 328294 75250 328350
rect 75306 328294 75374 328350
rect 75430 328294 75498 328350
rect 75554 328294 75622 328350
rect 75678 328294 93250 328350
rect 93306 328294 93374 328350
rect 93430 328294 93498 328350
rect 93554 328294 93622 328350
rect 93678 328294 111250 328350
rect 111306 328294 111374 328350
rect 111430 328294 111498 328350
rect 111554 328294 111622 328350
rect 111678 328294 129250 328350
rect 129306 328294 129374 328350
rect 129430 328294 129498 328350
rect 129554 328294 129622 328350
rect 129678 328294 147250 328350
rect 147306 328294 147374 328350
rect 147430 328294 147498 328350
rect 147554 328294 147622 328350
rect 147678 328294 165250 328350
rect 165306 328294 165374 328350
rect 165430 328294 165498 328350
rect 165554 328294 165622 328350
rect 165678 328294 183250 328350
rect 183306 328294 183374 328350
rect 183430 328294 183498 328350
rect 183554 328294 183622 328350
rect 183678 328294 201250 328350
rect 201306 328294 201374 328350
rect 201430 328294 201498 328350
rect 201554 328294 201622 328350
rect 201678 328294 204518 328350
rect 204574 328294 204642 328350
rect 204698 328294 235238 328350
rect 235294 328294 235362 328350
rect 235418 328294 265958 328350
rect 266014 328294 266082 328350
rect 266138 328294 296678 328350
rect 296734 328294 296802 328350
rect 296858 328294 327398 328350
rect 327454 328294 327522 328350
rect 327578 328294 358118 328350
rect 358174 328294 358242 328350
rect 358298 328294 388838 328350
rect 388894 328294 388962 328350
rect 389018 328294 419558 328350
rect 419614 328294 419682 328350
rect 419738 328294 450278 328350
rect 450334 328294 450402 328350
rect 450458 328294 480998 328350
rect 481054 328294 481122 328350
rect 481178 328294 507250 328350
rect 507306 328294 507374 328350
rect 507430 328294 507498 328350
rect 507554 328294 507622 328350
rect 507678 328294 525250 328350
rect 525306 328294 525374 328350
rect 525430 328294 525498 328350
rect 525554 328294 525622 328350
rect 525678 328294 543250 328350
rect 543306 328294 543374 328350
rect 543430 328294 543498 328350
rect 543554 328294 543622 328350
rect 543678 328294 561250 328350
rect 561306 328294 561374 328350
rect 561430 328294 561498 328350
rect 561554 328294 561622 328350
rect 561678 328294 579250 328350
rect 579306 328294 579374 328350
rect 579430 328294 579498 328350
rect 579554 328294 579622 328350
rect 579678 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 3250 328226
rect 3306 328170 3374 328226
rect 3430 328170 3498 328226
rect 3554 328170 3622 328226
rect 3678 328170 21250 328226
rect 21306 328170 21374 328226
rect 21430 328170 21498 328226
rect 21554 328170 21622 328226
rect 21678 328170 39250 328226
rect 39306 328170 39374 328226
rect 39430 328170 39498 328226
rect 39554 328170 39622 328226
rect 39678 328170 57250 328226
rect 57306 328170 57374 328226
rect 57430 328170 57498 328226
rect 57554 328170 57622 328226
rect 57678 328170 75250 328226
rect 75306 328170 75374 328226
rect 75430 328170 75498 328226
rect 75554 328170 75622 328226
rect 75678 328170 93250 328226
rect 93306 328170 93374 328226
rect 93430 328170 93498 328226
rect 93554 328170 93622 328226
rect 93678 328170 111250 328226
rect 111306 328170 111374 328226
rect 111430 328170 111498 328226
rect 111554 328170 111622 328226
rect 111678 328170 129250 328226
rect 129306 328170 129374 328226
rect 129430 328170 129498 328226
rect 129554 328170 129622 328226
rect 129678 328170 147250 328226
rect 147306 328170 147374 328226
rect 147430 328170 147498 328226
rect 147554 328170 147622 328226
rect 147678 328170 165250 328226
rect 165306 328170 165374 328226
rect 165430 328170 165498 328226
rect 165554 328170 165622 328226
rect 165678 328170 183250 328226
rect 183306 328170 183374 328226
rect 183430 328170 183498 328226
rect 183554 328170 183622 328226
rect 183678 328170 201250 328226
rect 201306 328170 201374 328226
rect 201430 328170 201498 328226
rect 201554 328170 201622 328226
rect 201678 328170 204518 328226
rect 204574 328170 204642 328226
rect 204698 328170 235238 328226
rect 235294 328170 235362 328226
rect 235418 328170 265958 328226
rect 266014 328170 266082 328226
rect 266138 328170 296678 328226
rect 296734 328170 296802 328226
rect 296858 328170 327398 328226
rect 327454 328170 327522 328226
rect 327578 328170 358118 328226
rect 358174 328170 358242 328226
rect 358298 328170 388838 328226
rect 388894 328170 388962 328226
rect 389018 328170 419558 328226
rect 419614 328170 419682 328226
rect 419738 328170 450278 328226
rect 450334 328170 450402 328226
rect 450458 328170 480998 328226
rect 481054 328170 481122 328226
rect 481178 328170 507250 328226
rect 507306 328170 507374 328226
rect 507430 328170 507498 328226
rect 507554 328170 507622 328226
rect 507678 328170 525250 328226
rect 525306 328170 525374 328226
rect 525430 328170 525498 328226
rect 525554 328170 525622 328226
rect 525678 328170 543250 328226
rect 543306 328170 543374 328226
rect 543430 328170 543498 328226
rect 543554 328170 543622 328226
rect 543678 328170 561250 328226
rect 561306 328170 561374 328226
rect 561430 328170 561498 328226
rect 561554 328170 561622 328226
rect 561678 328170 579250 328226
rect 579306 328170 579374 328226
rect 579430 328170 579498 328226
rect 579554 328170 579622 328226
rect 579678 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 3250 328102
rect 3306 328046 3374 328102
rect 3430 328046 3498 328102
rect 3554 328046 3622 328102
rect 3678 328046 21250 328102
rect 21306 328046 21374 328102
rect 21430 328046 21498 328102
rect 21554 328046 21622 328102
rect 21678 328046 39250 328102
rect 39306 328046 39374 328102
rect 39430 328046 39498 328102
rect 39554 328046 39622 328102
rect 39678 328046 57250 328102
rect 57306 328046 57374 328102
rect 57430 328046 57498 328102
rect 57554 328046 57622 328102
rect 57678 328046 75250 328102
rect 75306 328046 75374 328102
rect 75430 328046 75498 328102
rect 75554 328046 75622 328102
rect 75678 328046 93250 328102
rect 93306 328046 93374 328102
rect 93430 328046 93498 328102
rect 93554 328046 93622 328102
rect 93678 328046 111250 328102
rect 111306 328046 111374 328102
rect 111430 328046 111498 328102
rect 111554 328046 111622 328102
rect 111678 328046 129250 328102
rect 129306 328046 129374 328102
rect 129430 328046 129498 328102
rect 129554 328046 129622 328102
rect 129678 328046 147250 328102
rect 147306 328046 147374 328102
rect 147430 328046 147498 328102
rect 147554 328046 147622 328102
rect 147678 328046 165250 328102
rect 165306 328046 165374 328102
rect 165430 328046 165498 328102
rect 165554 328046 165622 328102
rect 165678 328046 183250 328102
rect 183306 328046 183374 328102
rect 183430 328046 183498 328102
rect 183554 328046 183622 328102
rect 183678 328046 201250 328102
rect 201306 328046 201374 328102
rect 201430 328046 201498 328102
rect 201554 328046 201622 328102
rect 201678 328046 204518 328102
rect 204574 328046 204642 328102
rect 204698 328046 235238 328102
rect 235294 328046 235362 328102
rect 235418 328046 265958 328102
rect 266014 328046 266082 328102
rect 266138 328046 296678 328102
rect 296734 328046 296802 328102
rect 296858 328046 327398 328102
rect 327454 328046 327522 328102
rect 327578 328046 358118 328102
rect 358174 328046 358242 328102
rect 358298 328046 388838 328102
rect 388894 328046 388962 328102
rect 389018 328046 419558 328102
rect 419614 328046 419682 328102
rect 419738 328046 450278 328102
rect 450334 328046 450402 328102
rect 450458 328046 480998 328102
rect 481054 328046 481122 328102
rect 481178 328046 507250 328102
rect 507306 328046 507374 328102
rect 507430 328046 507498 328102
rect 507554 328046 507622 328102
rect 507678 328046 525250 328102
rect 525306 328046 525374 328102
rect 525430 328046 525498 328102
rect 525554 328046 525622 328102
rect 525678 328046 543250 328102
rect 543306 328046 543374 328102
rect 543430 328046 543498 328102
rect 543554 328046 543622 328102
rect 543678 328046 561250 328102
rect 561306 328046 561374 328102
rect 561430 328046 561498 328102
rect 561554 328046 561622 328102
rect 561678 328046 579250 328102
rect 579306 328046 579374 328102
rect 579430 328046 579498 328102
rect 579554 328046 579622 328102
rect 579678 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 3250 327978
rect 3306 327922 3374 327978
rect 3430 327922 3498 327978
rect 3554 327922 3622 327978
rect 3678 327922 21250 327978
rect 21306 327922 21374 327978
rect 21430 327922 21498 327978
rect 21554 327922 21622 327978
rect 21678 327922 39250 327978
rect 39306 327922 39374 327978
rect 39430 327922 39498 327978
rect 39554 327922 39622 327978
rect 39678 327922 57250 327978
rect 57306 327922 57374 327978
rect 57430 327922 57498 327978
rect 57554 327922 57622 327978
rect 57678 327922 75250 327978
rect 75306 327922 75374 327978
rect 75430 327922 75498 327978
rect 75554 327922 75622 327978
rect 75678 327922 93250 327978
rect 93306 327922 93374 327978
rect 93430 327922 93498 327978
rect 93554 327922 93622 327978
rect 93678 327922 111250 327978
rect 111306 327922 111374 327978
rect 111430 327922 111498 327978
rect 111554 327922 111622 327978
rect 111678 327922 129250 327978
rect 129306 327922 129374 327978
rect 129430 327922 129498 327978
rect 129554 327922 129622 327978
rect 129678 327922 147250 327978
rect 147306 327922 147374 327978
rect 147430 327922 147498 327978
rect 147554 327922 147622 327978
rect 147678 327922 165250 327978
rect 165306 327922 165374 327978
rect 165430 327922 165498 327978
rect 165554 327922 165622 327978
rect 165678 327922 183250 327978
rect 183306 327922 183374 327978
rect 183430 327922 183498 327978
rect 183554 327922 183622 327978
rect 183678 327922 201250 327978
rect 201306 327922 201374 327978
rect 201430 327922 201498 327978
rect 201554 327922 201622 327978
rect 201678 327922 204518 327978
rect 204574 327922 204642 327978
rect 204698 327922 235238 327978
rect 235294 327922 235362 327978
rect 235418 327922 265958 327978
rect 266014 327922 266082 327978
rect 266138 327922 296678 327978
rect 296734 327922 296802 327978
rect 296858 327922 327398 327978
rect 327454 327922 327522 327978
rect 327578 327922 358118 327978
rect 358174 327922 358242 327978
rect 358298 327922 388838 327978
rect 388894 327922 388962 327978
rect 389018 327922 419558 327978
rect 419614 327922 419682 327978
rect 419738 327922 450278 327978
rect 450334 327922 450402 327978
rect 450458 327922 480998 327978
rect 481054 327922 481122 327978
rect 481178 327922 507250 327978
rect 507306 327922 507374 327978
rect 507430 327922 507498 327978
rect 507554 327922 507622 327978
rect 507678 327922 525250 327978
rect 525306 327922 525374 327978
rect 525430 327922 525498 327978
rect 525554 327922 525622 327978
rect 525678 327922 543250 327978
rect 543306 327922 543374 327978
rect 543430 327922 543498 327978
rect 543554 327922 543622 327978
rect 543678 327922 561250 327978
rect 561306 327922 561374 327978
rect 561430 327922 561498 327978
rect 561554 327922 561622 327978
rect 561678 327922 579250 327978
rect 579306 327922 579374 327978
rect 579430 327922 579498 327978
rect 579554 327922 579622 327978
rect 579678 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 6970 316350
rect 7026 316294 7094 316350
rect 7150 316294 7218 316350
rect 7274 316294 7342 316350
rect 7398 316294 24970 316350
rect 25026 316294 25094 316350
rect 25150 316294 25218 316350
rect 25274 316294 25342 316350
rect 25398 316294 42970 316350
rect 43026 316294 43094 316350
rect 43150 316294 43218 316350
rect 43274 316294 43342 316350
rect 43398 316294 60970 316350
rect 61026 316294 61094 316350
rect 61150 316294 61218 316350
rect 61274 316294 61342 316350
rect 61398 316294 78970 316350
rect 79026 316294 79094 316350
rect 79150 316294 79218 316350
rect 79274 316294 79342 316350
rect 79398 316294 96970 316350
rect 97026 316294 97094 316350
rect 97150 316294 97218 316350
rect 97274 316294 97342 316350
rect 97398 316294 114970 316350
rect 115026 316294 115094 316350
rect 115150 316294 115218 316350
rect 115274 316294 115342 316350
rect 115398 316294 132970 316350
rect 133026 316294 133094 316350
rect 133150 316294 133218 316350
rect 133274 316294 133342 316350
rect 133398 316294 150970 316350
rect 151026 316294 151094 316350
rect 151150 316294 151218 316350
rect 151274 316294 151342 316350
rect 151398 316294 168970 316350
rect 169026 316294 169094 316350
rect 169150 316294 169218 316350
rect 169274 316294 169342 316350
rect 169398 316294 186970 316350
rect 187026 316294 187094 316350
rect 187150 316294 187218 316350
rect 187274 316294 187342 316350
rect 187398 316294 219878 316350
rect 219934 316294 220002 316350
rect 220058 316294 250598 316350
rect 250654 316294 250722 316350
rect 250778 316294 281318 316350
rect 281374 316294 281442 316350
rect 281498 316294 312038 316350
rect 312094 316294 312162 316350
rect 312218 316294 342758 316350
rect 342814 316294 342882 316350
rect 342938 316294 373478 316350
rect 373534 316294 373602 316350
rect 373658 316294 404198 316350
rect 404254 316294 404322 316350
rect 404378 316294 434918 316350
rect 434974 316294 435042 316350
rect 435098 316294 465638 316350
rect 465694 316294 465762 316350
rect 465818 316294 496358 316350
rect 496414 316294 496482 316350
rect 496538 316294 510970 316350
rect 511026 316294 511094 316350
rect 511150 316294 511218 316350
rect 511274 316294 511342 316350
rect 511398 316294 528970 316350
rect 529026 316294 529094 316350
rect 529150 316294 529218 316350
rect 529274 316294 529342 316350
rect 529398 316294 546970 316350
rect 547026 316294 547094 316350
rect 547150 316294 547218 316350
rect 547274 316294 547342 316350
rect 547398 316294 564970 316350
rect 565026 316294 565094 316350
rect 565150 316294 565218 316350
rect 565274 316294 565342 316350
rect 565398 316294 582970 316350
rect 583026 316294 583094 316350
rect 583150 316294 583218 316350
rect 583274 316294 583342 316350
rect 583398 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 6970 316226
rect 7026 316170 7094 316226
rect 7150 316170 7218 316226
rect 7274 316170 7342 316226
rect 7398 316170 24970 316226
rect 25026 316170 25094 316226
rect 25150 316170 25218 316226
rect 25274 316170 25342 316226
rect 25398 316170 42970 316226
rect 43026 316170 43094 316226
rect 43150 316170 43218 316226
rect 43274 316170 43342 316226
rect 43398 316170 60970 316226
rect 61026 316170 61094 316226
rect 61150 316170 61218 316226
rect 61274 316170 61342 316226
rect 61398 316170 78970 316226
rect 79026 316170 79094 316226
rect 79150 316170 79218 316226
rect 79274 316170 79342 316226
rect 79398 316170 96970 316226
rect 97026 316170 97094 316226
rect 97150 316170 97218 316226
rect 97274 316170 97342 316226
rect 97398 316170 114970 316226
rect 115026 316170 115094 316226
rect 115150 316170 115218 316226
rect 115274 316170 115342 316226
rect 115398 316170 132970 316226
rect 133026 316170 133094 316226
rect 133150 316170 133218 316226
rect 133274 316170 133342 316226
rect 133398 316170 150970 316226
rect 151026 316170 151094 316226
rect 151150 316170 151218 316226
rect 151274 316170 151342 316226
rect 151398 316170 168970 316226
rect 169026 316170 169094 316226
rect 169150 316170 169218 316226
rect 169274 316170 169342 316226
rect 169398 316170 186970 316226
rect 187026 316170 187094 316226
rect 187150 316170 187218 316226
rect 187274 316170 187342 316226
rect 187398 316170 219878 316226
rect 219934 316170 220002 316226
rect 220058 316170 250598 316226
rect 250654 316170 250722 316226
rect 250778 316170 281318 316226
rect 281374 316170 281442 316226
rect 281498 316170 312038 316226
rect 312094 316170 312162 316226
rect 312218 316170 342758 316226
rect 342814 316170 342882 316226
rect 342938 316170 373478 316226
rect 373534 316170 373602 316226
rect 373658 316170 404198 316226
rect 404254 316170 404322 316226
rect 404378 316170 434918 316226
rect 434974 316170 435042 316226
rect 435098 316170 465638 316226
rect 465694 316170 465762 316226
rect 465818 316170 496358 316226
rect 496414 316170 496482 316226
rect 496538 316170 510970 316226
rect 511026 316170 511094 316226
rect 511150 316170 511218 316226
rect 511274 316170 511342 316226
rect 511398 316170 528970 316226
rect 529026 316170 529094 316226
rect 529150 316170 529218 316226
rect 529274 316170 529342 316226
rect 529398 316170 546970 316226
rect 547026 316170 547094 316226
rect 547150 316170 547218 316226
rect 547274 316170 547342 316226
rect 547398 316170 564970 316226
rect 565026 316170 565094 316226
rect 565150 316170 565218 316226
rect 565274 316170 565342 316226
rect 565398 316170 582970 316226
rect 583026 316170 583094 316226
rect 583150 316170 583218 316226
rect 583274 316170 583342 316226
rect 583398 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 6970 316102
rect 7026 316046 7094 316102
rect 7150 316046 7218 316102
rect 7274 316046 7342 316102
rect 7398 316046 24970 316102
rect 25026 316046 25094 316102
rect 25150 316046 25218 316102
rect 25274 316046 25342 316102
rect 25398 316046 42970 316102
rect 43026 316046 43094 316102
rect 43150 316046 43218 316102
rect 43274 316046 43342 316102
rect 43398 316046 60970 316102
rect 61026 316046 61094 316102
rect 61150 316046 61218 316102
rect 61274 316046 61342 316102
rect 61398 316046 78970 316102
rect 79026 316046 79094 316102
rect 79150 316046 79218 316102
rect 79274 316046 79342 316102
rect 79398 316046 96970 316102
rect 97026 316046 97094 316102
rect 97150 316046 97218 316102
rect 97274 316046 97342 316102
rect 97398 316046 114970 316102
rect 115026 316046 115094 316102
rect 115150 316046 115218 316102
rect 115274 316046 115342 316102
rect 115398 316046 132970 316102
rect 133026 316046 133094 316102
rect 133150 316046 133218 316102
rect 133274 316046 133342 316102
rect 133398 316046 150970 316102
rect 151026 316046 151094 316102
rect 151150 316046 151218 316102
rect 151274 316046 151342 316102
rect 151398 316046 168970 316102
rect 169026 316046 169094 316102
rect 169150 316046 169218 316102
rect 169274 316046 169342 316102
rect 169398 316046 186970 316102
rect 187026 316046 187094 316102
rect 187150 316046 187218 316102
rect 187274 316046 187342 316102
rect 187398 316046 219878 316102
rect 219934 316046 220002 316102
rect 220058 316046 250598 316102
rect 250654 316046 250722 316102
rect 250778 316046 281318 316102
rect 281374 316046 281442 316102
rect 281498 316046 312038 316102
rect 312094 316046 312162 316102
rect 312218 316046 342758 316102
rect 342814 316046 342882 316102
rect 342938 316046 373478 316102
rect 373534 316046 373602 316102
rect 373658 316046 404198 316102
rect 404254 316046 404322 316102
rect 404378 316046 434918 316102
rect 434974 316046 435042 316102
rect 435098 316046 465638 316102
rect 465694 316046 465762 316102
rect 465818 316046 496358 316102
rect 496414 316046 496482 316102
rect 496538 316046 510970 316102
rect 511026 316046 511094 316102
rect 511150 316046 511218 316102
rect 511274 316046 511342 316102
rect 511398 316046 528970 316102
rect 529026 316046 529094 316102
rect 529150 316046 529218 316102
rect 529274 316046 529342 316102
rect 529398 316046 546970 316102
rect 547026 316046 547094 316102
rect 547150 316046 547218 316102
rect 547274 316046 547342 316102
rect 547398 316046 564970 316102
rect 565026 316046 565094 316102
rect 565150 316046 565218 316102
rect 565274 316046 565342 316102
rect 565398 316046 582970 316102
rect 583026 316046 583094 316102
rect 583150 316046 583218 316102
rect 583274 316046 583342 316102
rect 583398 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 6970 315978
rect 7026 315922 7094 315978
rect 7150 315922 7218 315978
rect 7274 315922 7342 315978
rect 7398 315922 24970 315978
rect 25026 315922 25094 315978
rect 25150 315922 25218 315978
rect 25274 315922 25342 315978
rect 25398 315922 42970 315978
rect 43026 315922 43094 315978
rect 43150 315922 43218 315978
rect 43274 315922 43342 315978
rect 43398 315922 60970 315978
rect 61026 315922 61094 315978
rect 61150 315922 61218 315978
rect 61274 315922 61342 315978
rect 61398 315922 78970 315978
rect 79026 315922 79094 315978
rect 79150 315922 79218 315978
rect 79274 315922 79342 315978
rect 79398 315922 96970 315978
rect 97026 315922 97094 315978
rect 97150 315922 97218 315978
rect 97274 315922 97342 315978
rect 97398 315922 114970 315978
rect 115026 315922 115094 315978
rect 115150 315922 115218 315978
rect 115274 315922 115342 315978
rect 115398 315922 132970 315978
rect 133026 315922 133094 315978
rect 133150 315922 133218 315978
rect 133274 315922 133342 315978
rect 133398 315922 150970 315978
rect 151026 315922 151094 315978
rect 151150 315922 151218 315978
rect 151274 315922 151342 315978
rect 151398 315922 168970 315978
rect 169026 315922 169094 315978
rect 169150 315922 169218 315978
rect 169274 315922 169342 315978
rect 169398 315922 186970 315978
rect 187026 315922 187094 315978
rect 187150 315922 187218 315978
rect 187274 315922 187342 315978
rect 187398 315922 219878 315978
rect 219934 315922 220002 315978
rect 220058 315922 250598 315978
rect 250654 315922 250722 315978
rect 250778 315922 281318 315978
rect 281374 315922 281442 315978
rect 281498 315922 312038 315978
rect 312094 315922 312162 315978
rect 312218 315922 342758 315978
rect 342814 315922 342882 315978
rect 342938 315922 373478 315978
rect 373534 315922 373602 315978
rect 373658 315922 404198 315978
rect 404254 315922 404322 315978
rect 404378 315922 434918 315978
rect 434974 315922 435042 315978
rect 435098 315922 465638 315978
rect 465694 315922 465762 315978
rect 465818 315922 496358 315978
rect 496414 315922 496482 315978
rect 496538 315922 510970 315978
rect 511026 315922 511094 315978
rect 511150 315922 511218 315978
rect 511274 315922 511342 315978
rect 511398 315922 528970 315978
rect 529026 315922 529094 315978
rect 529150 315922 529218 315978
rect 529274 315922 529342 315978
rect 529398 315922 546970 315978
rect 547026 315922 547094 315978
rect 547150 315922 547218 315978
rect 547274 315922 547342 315978
rect 547398 315922 564970 315978
rect 565026 315922 565094 315978
rect 565150 315922 565218 315978
rect 565274 315922 565342 315978
rect 565398 315922 582970 315978
rect 583026 315922 583094 315978
rect 583150 315922 583218 315978
rect 583274 315922 583342 315978
rect 583398 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 3250 310350
rect 3306 310294 3374 310350
rect 3430 310294 3498 310350
rect 3554 310294 3622 310350
rect 3678 310294 21250 310350
rect 21306 310294 21374 310350
rect 21430 310294 21498 310350
rect 21554 310294 21622 310350
rect 21678 310294 39250 310350
rect 39306 310294 39374 310350
rect 39430 310294 39498 310350
rect 39554 310294 39622 310350
rect 39678 310294 57250 310350
rect 57306 310294 57374 310350
rect 57430 310294 57498 310350
rect 57554 310294 57622 310350
rect 57678 310294 75250 310350
rect 75306 310294 75374 310350
rect 75430 310294 75498 310350
rect 75554 310294 75622 310350
rect 75678 310294 93250 310350
rect 93306 310294 93374 310350
rect 93430 310294 93498 310350
rect 93554 310294 93622 310350
rect 93678 310294 111250 310350
rect 111306 310294 111374 310350
rect 111430 310294 111498 310350
rect 111554 310294 111622 310350
rect 111678 310294 129250 310350
rect 129306 310294 129374 310350
rect 129430 310294 129498 310350
rect 129554 310294 129622 310350
rect 129678 310294 147250 310350
rect 147306 310294 147374 310350
rect 147430 310294 147498 310350
rect 147554 310294 147622 310350
rect 147678 310294 165250 310350
rect 165306 310294 165374 310350
rect 165430 310294 165498 310350
rect 165554 310294 165622 310350
rect 165678 310294 183250 310350
rect 183306 310294 183374 310350
rect 183430 310294 183498 310350
rect 183554 310294 183622 310350
rect 183678 310294 201250 310350
rect 201306 310294 201374 310350
rect 201430 310294 201498 310350
rect 201554 310294 201622 310350
rect 201678 310294 204518 310350
rect 204574 310294 204642 310350
rect 204698 310294 235238 310350
rect 235294 310294 235362 310350
rect 235418 310294 265958 310350
rect 266014 310294 266082 310350
rect 266138 310294 296678 310350
rect 296734 310294 296802 310350
rect 296858 310294 327398 310350
rect 327454 310294 327522 310350
rect 327578 310294 358118 310350
rect 358174 310294 358242 310350
rect 358298 310294 388838 310350
rect 388894 310294 388962 310350
rect 389018 310294 419558 310350
rect 419614 310294 419682 310350
rect 419738 310294 450278 310350
rect 450334 310294 450402 310350
rect 450458 310294 480998 310350
rect 481054 310294 481122 310350
rect 481178 310294 507250 310350
rect 507306 310294 507374 310350
rect 507430 310294 507498 310350
rect 507554 310294 507622 310350
rect 507678 310294 525250 310350
rect 525306 310294 525374 310350
rect 525430 310294 525498 310350
rect 525554 310294 525622 310350
rect 525678 310294 543250 310350
rect 543306 310294 543374 310350
rect 543430 310294 543498 310350
rect 543554 310294 543622 310350
rect 543678 310294 561250 310350
rect 561306 310294 561374 310350
rect 561430 310294 561498 310350
rect 561554 310294 561622 310350
rect 561678 310294 579250 310350
rect 579306 310294 579374 310350
rect 579430 310294 579498 310350
rect 579554 310294 579622 310350
rect 579678 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 3250 310226
rect 3306 310170 3374 310226
rect 3430 310170 3498 310226
rect 3554 310170 3622 310226
rect 3678 310170 21250 310226
rect 21306 310170 21374 310226
rect 21430 310170 21498 310226
rect 21554 310170 21622 310226
rect 21678 310170 39250 310226
rect 39306 310170 39374 310226
rect 39430 310170 39498 310226
rect 39554 310170 39622 310226
rect 39678 310170 57250 310226
rect 57306 310170 57374 310226
rect 57430 310170 57498 310226
rect 57554 310170 57622 310226
rect 57678 310170 75250 310226
rect 75306 310170 75374 310226
rect 75430 310170 75498 310226
rect 75554 310170 75622 310226
rect 75678 310170 93250 310226
rect 93306 310170 93374 310226
rect 93430 310170 93498 310226
rect 93554 310170 93622 310226
rect 93678 310170 111250 310226
rect 111306 310170 111374 310226
rect 111430 310170 111498 310226
rect 111554 310170 111622 310226
rect 111678 310170 129250 310226
rect 129306 310170 129374 310226
rect 129430 310170 129498 310226
rect 129554 310170 129622 310226
rect 129678 310170 147250 310226
rect 147306 310170 147374 310226
rect 147430 310170 147498 310226
rect 147554 310170 147622 310226
rect 147678 310170 165250 310226
rect 165306 310170 165374 310226
rect 165430 310170 165498 310226
rect 165554 310170 165622 310226
rect 165678 310170 183250 310226
rect 183306 310170 183374 310226
rect 183430 310170 183498 310226
rect 183554 310170 183622 310226
rect 183678 310170 201250 310226
rect 201306 310170 201374 310226
rect 201430 310170 201498 310226
rect 201554 310170 201622 310226
rect 201678 310170 204518 310226
rect 204574 310170 204642 310226
rect 204698 310170 235238 310226
rect 235294 310170 235362 310226
rect 235418 310170 265958 310226
rect 266014 310170 266082 310226
rect 266138 310170 296678 310226
rect 296734 310170 296802 310226
rect 296858 310170 327398 310226
rect 327454 310170 327522 310226
rect 327578 310170 358118 310226
rect 358174 310170 358242 310226
rect 358298 310170 388838 310226
rect 388894 310170 388962 310226
rect 389018 310170 419558 310226
rect 419614 310170 419682 310226
rect 419738 310170 450278 310226
rect 450334 310170 450402 310226
rect 450458 310170 480998 310226
rect 481054 310170 481122 310226
rect 481178 310170 507250 310226
rect 507306 310170 507374 310226
rect 507430 310170 507498 310226
rect 507554 310170 507622 310226
rect 507678 310170 525250 310226
rect 525306 310170 525374 310226
rect 525430 310170 525498 310226
rect 525554 310170 525622 310226
rect 525678 310170 543250 310226
rect 543306 310170 543374 310226
rect 543430 310170 543498 310226
rect 543554 310170 543622 310226
rect 543678 310170 561250 310226
rect 561306 310170 561374 310226
rect 561430 310170 561498 310226
rect 561554 310170 561622 310226
rect 561678 310170 579250 310226
rect 579306 310170 579374 310226
rect 579430 310170 579498 310226
rect 579554 310170 579622 310226
rect 579678 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 3250 310102
rect 3306 310046 3374 310102
rect 3430 310046 3498 310102
rect 3554 310046 3622 310102
rect 3678 310046 21250 310102
rect 21306 310046 21374 310102
rect 21430 310046 21498 310102
rect 21554 310046 21622 310102
rect 21678 310046 39250 310102
rect 39306 310046 39374 310102
rect 39430 310046 39498 310102
rect 39554 310046 39622 310102
rect 39678 310046 57250 310102
rect 57306 310046 57374 310102
rect 57430 310046 57498 310102
rect 57554 310046 57622 310102
rect 57678 310046 75250 310102
rect 75306 310046 75374 310102
rect 75430 310046 75498 310102
rect 75554 310046 75622 310102
rect 75678 310046 93250 310102
rect 93306 310046 93374 310102
rect 93430 310046 93498 310102
rect 93554 310046 93622 310102
rect 93678 310046 111250 310102
rect 111306 310046 111374 310102
rect 111430 310046 111498 310102
rect 111554 310046 111622 310102
rect 111678 310046 129250 310102
rect 129306 310046 129374 310102
rect 129430 310046 129498 310102
rect 129554 310046 129622 310102
rect 129678 310046 147250 310102
rect 147306 310046 147374 310102
rect 147430 310046 147498 310102
rect 147554 310046 147622 310102
rect 147678 310046 165250 310102
rect 165306 310046 165374 310102
rect 165430 310046 165498 310102
rect 165554 310046 165622 310102
rect 165678 310046 183250 310102
rect 183306 310046 183374 310102
rect 183430 310046 183498 310102
rect 183554 310046 183622 310102
rect 183678 310046 201250 310102
rect 201306 310046 201374 310102
rect 201430 310046 201498 310102
rect 201554 310046 201622 310102
rect 201678 310046 204518 310102
rect 204574 310046 204642 310102
rect 204698 310046 235238 310102
rect 235294 310046 235362 310102
rect 235418 310046 265958 310102
rect 266014 310046 266082 310102
rect 266138 310046 296678 310102
rect 296734 310046 296802 310102
rect 296858 310046 327398 310102
rect 327454 310046 327522 310102
rect 327578 310046 358118 310102
rect 358174 310046 358242 310102
rect 358298 310046 388838 310102
rect 388894 310046 388962 310102
rect 389018 310046 419558 310102
rect 419614 310046 419682 310102
rect 419738 310046 450278 310102
rect 450334 310046 450402 310102
rect 450458 310046 480998 310102
rect 481054 310046 481122 310102
rect 481178 310046 507250 310102
rect 507306 310046 507374 310102
rect 507430 310046 507498 310102
rect 507554 310046 507622 310102
rect 507678 310046 525250 310102
rect 525306 310046 525374 310102
rect 525430 310046 525498 310102
rect 525554 310046 525622 310102
rect 525678 310046 543250 310102
rect 543306 310046 543374 310102
rect 543430 310046 543498 310102
rect 543554 310046 543622 310102
rect 543678 310046 561250 310102
rect 561306 310046 561374 310102
rect 561430 310046 561498 310102
rect 561554 310046 561622 310102
rect 561678 310046 579250 310102
rect 579306 310046 579374 310102
rect 579430 310046 579498 310102
rect 579554 310046 579622 310102
rect 579678 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 3250 309978
rect 3306 309922 3374 309978
rect 3430 309922 3498 309978
rect 3554 309922 3622 309978
rect 3678 309922 21250 309978
rect 21306 309922 21374 309978
rect 21430 309922 21498 309978
rect 21554 309922 21622 309978
rect 21678 309922 39250 309978
rect 39306 309922 39374 309978
rect 39430 309922 39498 309978
rect 39554 309922 39622 309978
rect 39678 309922 57250 309978
rect 57306 309922 57374 309978
rect 57430 309922 57498 309978
rect 57554 309922 57622 309978
rect 57678 309922 75250 309978
rect 75306 309922 75374 309978
rect 75430 309922 75498 309978
rect 75554 309922 75622 309978
rect 75678 309922 93250 309978
rect 93306 309922 93374 309978
rect 93430 309922 93498 309978
rect 93554 309922 93622 309978
rect 93678 309922 111250 309978
rect 111306 309922 111374 309978
rect 111430 309922 111498 309978
rect 111554 309922 111622 309978
rect 111678 309922 129250 309978
rect 129306 309922 129374 309978
rect 129430 309922 129498 309978
rect 129554 309922 129622 309978
rect 129678 309922 147250 309978
rect 147306 309922 147374 309978
rect 147430 309922 147498 309978
rect 147554 309922 147622 309978
rect 147678 309922 165250 309978
rect 165306 309922 165374 309978
rect 165430 309922 165498 309978
rect 165554 309922 165622 309978
rect 165678 309922 183250 309978
rect 183306 309922 183374 309978
rect 183430 309922 183498 309978
rect 183554 309922 183622 309978
rect 183678 309922 201250 309978
rect 201306 309922 201374 309978
rect 201430 309922 201498 309978
rect 201554 309922 201622 309978
rect 201678 309922 204518 309978
rect 204574 309922 204642 309978
rect 204698 309922 235238 309978
rect 235294 309922 235362 309978
rect 235418 309922 265958 309978
rect 266014 309922 266082 309978
rect 266138 309922 296678 309978
rect 296734 309922 296802 309978
rect 296858 309922 327398 309978
rect 327454 309922 327522 309978
rect 327578 309922 358118 309978
rect 358174 309922 358242 309978
rect 358298 309922 388838 309978
rect 388894 309922 388962 309978
rect 389018 309922 419558 309978
rect 419614 309922 419682 309978
rect 419738 309922 450278 309978
rect 450334 309922 450402 309978
rect 450458 309922 480998 309978
rect 481054 309922 481122 309978
rect 481178 309922 507250 309978
rect 507306 309922 507374 309978
rect 507430 309922 507498 309978
rect 507554 309922 507622 309978
rect 507678 309922 525250 309978
rect 525306 309922 525374 309978
rect 525430 309922 525498 309978
rect 525554 309922 525622 309978
rect 525678 309922 543250 309978
rect 543306 309922 543374 309978
rect 543430 309922 543498 309978
rect 543554 309922 543622 309978
rect 543678 309922 561250 309978
rect 561306 309922 561374 309978
rect 561430 309922 561498 309978
rect 561554 309922 561622 309978
rect 561678 309922 579250 309978
rect 579306 309922 579374 309978
rect 579430 309922 579498 309978
rect 579554 309922 579622 309978
rect 579678 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 6970 298350
rect 7026 298294 7094 298350
rect 7150 298294 7218 298350
rect 7274 298294 7342 298350
rect 7398 298294 24970 298350
rect 25026 298294 25094 298350
rect 25150 298294 25218 298350
rect 25274 298294 25342 298350
rect 25398 298294 42970 298350
rect 43026 298294 43094 298350
rect 43150 298294 43218 298350
rect 43274 298294 43342 298350
rect 43398 298294 60970 298350
rect 61026 298294 61094 298350
rect 61150 298294 61218 298350
rect 61274 298294 61342 298350
rect 61398 298294 78970 298350
rect 79026 298294 79094 298350
rect 79150 298294 79218 298350
rect 79274 298294 79342 298350
rect 79398 298294 96970 298350
rect 97026 298294 97094 298350
rect 97150 298294 97218 298350
rect 97274 298294 97342 298350
rect 97398 298294 114970 298350
rect 115026 298294 115094 298350
rect 115150 298294 115218 298350
rect 115274 298294 115342 298350
rect 115398 298294 132970 298350
rect 133026 298294 133094 298350
rect 133150 298294 133218 298350
rect 133274 298294 133342 298350
rect 133398 298294 150970 298350
rect 151026 298294 151094 298350
rect 151150 298294 151218 298350
rect 151274 298294 151342 298350
rect 151398 298294 168970 298350
rect 169026 298294 169094 298350
rect 169150 298294 169218 298350
rect 169274 298294 169342 298350
rect 169398 298294 186970 298350
rect 187026 298294 187094 298350
rect 187150 298294 187218 298350
rect 187274 298294 187342 298350
rect 187398 298294 219878 298350
rect 219934 298294 220002 298350
rect 220058 298294 250598 298350
rect 250654 298294 250722 298350
rect 250778 298294 281318 298350
rect 281374 298294 281442 298350
rect 281498 298294 312038 298350
rect 312094 298294 312162 298350
rect 312218 298294 342758 298350
rect 342814 298294 342882 298350
rect 342938 298294 373478 298350
rect 373534 298294 373602 298350
rect 373658 298294 404198 298350
rect 404254 298294 404322 298350
rect 404378 298294 434918 298350
rect 434974 298294 435042 298350
rect 435098 298294 465638 298350
rect 465694 298294 465762 298350
rect 465818 298294 496358 298350
rect 496414 298294 496482 298350
rect 496538 298294 510970 298350
rect 511026 298294 511094 298350
rect 511150 298294 511218 298350
rect 511274 298294 511342 298350
rect 511398 298294 528970 298350
rect 529026 298294 529094 298350
rect 529150 298294 529218 298350
rect 529274 298294 529342 298350
rect 529398 298294 546970 298350
rect 547026 298294 547094 298350
rect 547150 298294 547218 298350
rect 547274 298294 547342 298350
rect 547398 298294 564970 298350
rect 565026 298294 565094 298350
rect 565150 298294 565218 298350
rect 565274 298294 565342 298350
rect 565398 298294 582970 298350
rect 583026 298294 583094 298350
rect 583150 298294 583218 298350
rect 583274 298294 583342 298350
rect 583398 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 6970 298226
rect 7026 298170 7094 298226
rect 7150 298170 7218 298226
rect 7274 298170 7342 298226
rect 7398 298170 24970 298226
rect 25026 298170 25094 298226
rect 25150 298170 25218 298226
rect 25274 298170 25342 298226
rect 25398 298170 42970 298226
rect 43026 298170 43094 298226
rect 43150 298170 43218 298226
rect 43274 298170 43342 298226
rect 43398 298170 60970 298226
rect 61026 298170 61094 298226
rect 61150 298170 61218 298226
rect 61274 298170 61342 298226
rect 61398 298170 78970 298226
rect 79026 298170 79094 298226
rect 79150 298170 79218 298226
rect 79274 298170 79342 298226
rect 79398 298170 96970 298226
rect 97026 298170 97094 298226
rect 97150 298170 97218 298226
rect 97274 298170 97342 298226
rect 97398 298170 114970 298226
rect 115026 298170 115094 298226
rect 115150 298170 115218 298226
rect 115274 298170 115342 298226
rect 115398 298170 132970 298226
rect 133026 298170 133094 298226
rect 133150 298170 133218 298226
rect 133274 298170 133342 298226
rect 133398 298170 150970 298226
rect 151026 298170 151094 298226
rect 151150 298170 151218 298226
rect 151274 298170 151342 298226
rect 151398 298170 168970 298226
rect 169026 298170 169094 298226
rect 169150 298170 169218 298226
rect 169274 298170 169342 298226
rect 169398 298170 186970 298226
rect 187026 298170 187094 298226
rect 187150 298170 187218 298226
rect 187274 298170 187342 298226
rect 187398 298170 219878 298226
rect 219934 298170 220002 298226
rect 220058 298170 250598 298226
rect 250654 298170 250722 298226
rect 250778 298170 281318 298226
rect 281374 298170 281442 298226
rect 281498 298170 312038 298226
rect 312094 298170 312162 298226
rect 312218 298170 342758 298226
rect 342814 298170 342882 298226
rect 342938 298170 373478 298226
rect 373534 298170 373602 298226
rect 373658 298170 404198 298226
rect 404254 298170 404322 298226
rect 404378 298170 434918 298226
rect 434974 298170 435042 298226
rect 435098 298170 465638 298226
rect 465694 298170 465762 298226
rect 465818 298170 496358 298226
rect 496414 298170 496482 298226
rect 496538 298170 510970 298226
rect 511026 298170 511094 298226
rect 511150 298170 511218 298226
rect 511274 298170 511342 298226
rect 511398 298170 528970 298226
rect 529026 298170 529094 298226
rect 529150 298170 529218 298226
rect 529274 298170 529342 298226
rect 529398 298170 546970 298226
rect 547026 298170 547094 298226
rect 547150 298170 547218 298226
rect 547274 298170 547342 298226
rect 547398 298170 564970 298226
rect 565026 298170 565094 298226
rect 565150 298170 565218 298226
rect 565274 298170 565342 298226
rect 565398 298170 582970 298226
rect 583026 298170 583094 298226
rect 583150 298170 583218 298226
rect 583274 298170 583342 298226
rect 583398 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 6970 298102
rect 7026 298046 7094 298102
rect 7150 298046 7218 298102
rect 7274 298046 7342 298102
rect 7398 298046 24970 298102
rect 25026 298046 25094 298102
rect 25150 298046 25218 298102
rect 25274 298046 25342 298102
rect 25398 298046 42970 298102
rect 43026 298046 43094 298102
rect 43150 298046 43218 298102
rect 43274 298046 43342 298102
rect 43398 298046 60970 298102
rect 61026 298046 61094 298102
rect 61150 298046 61218 298102
rect 61274 298046 61342 298102
rect 61398 298046 78970 298102
rect 79026 298046 79094 298102
rect 79150 298046 79218 298102
rect 79274 298046 79342 298102
rect 79398 298046 96970 298102
rect 97026 298046 97094 298102
rect 97150 298046 97218 298102
rect 97274 298046 97342 298102
rect 97398 298046 114970 298102
rect 115026 298046 115094 298102
rect 115150 298046 115218 298102
rect 115274 298046 115342 298102
rect 115398 298046 132970 298102
rect 133026 298046 133094 298102
rect 133150 298046 133218 298102
rect 133274 298046 133342 298102
rect 133398 298046 150970 298102
rect 151026 298046 151094 298102
rect 151150 298046 151218 298102
rect 151274 298046 151342 298102
rect 151398 298046 168970 298102
rect 169026 298046 169094 298102
rect 169150 298046 169218 298102
rect 169274 298046 169342 298102
rect 169398 298046 186970 298102
rect 187026 298046 187094 298102
rect 187150 298046 187218 298102
rect 187274 298046 187342 298102
rect 187398 298046 219878 298102
rect 219934 298046 220002 298102
rect 220058 298046 250598 298102
rect 250654 298046 250722 298102
rect 250778 298046 281318 298102
rect 281374 298046 281442 298102
rect 281498 298046 312038 298102
rect 312094 298046 312162 298102
rect 312218 298046 342758 298102
rect 342814 298046 342882 298102
rect 342938 298046 373478 298102
rect 373534 298046 373602 298102
rect 373658 298046 404198 298102
rect 404254 298046 404322 298102
rect 404378 298046 434918 298102
rect 434974 298046 435042 298102
rect 435098 298046 465638 298102
rect 465694 298046 465762 298102
rect 465818 298046 496358 298102
rect 496414 298046 496482 298102
rect 496538 298046 510970 298102
rect 511026 298046 511094 298102
rect 511150 298046 511218 298102
rect 511274 298046 511342 298102
rect 511398 298046 528970 298102
rect 529026 298046 529094 298102
rect 529150 298046 529218 298102
rect 529274 298046 529342 298102
rect 529398 298046 546970 298102
rect 547026 298046 547094 298102
rect 547150 298046 547218 298102
rect 547274 298046 547342 298102
rect 547398 298046 564970 298102
rect 565026 298046 565094 298102
rect 565150 298046 565218 298102
rect 565274 298046 565342 298102
rect 565398 298046 582970 298102
rect 583026 298046 583094 298102
rect 583150 298046 583218 298102
rect 583274 298046 583342 298102
rect 583398 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 6970 297978
rect 7026 297922 7094 297978
rect 7150 297922 7218 297978
rect 7274 297922 7342 297978
rect 7398 297922 24970 297978
rect 25026 297922 25094 297978
rect 25150 297922 25218 297978
rect 25274 297922 25342 297978
rect 25398 297922 42970 297978
rect 43026 297922 43094 297978
rect 43150 297922 43218 297978
rect 43274 297922 43342 297978
rect 43398 297922 60970 297978
rect 61026 297922 61094 297978
rect 61150 297922 61218 297978
rect 61274 297922 61342 297978
rect 61398 297922 78970 297978
rect 79026 297922 79094 297978
rect 79150 297922 79218 297978
rect 79274 297922 79342 297978
rect 79398 297922 96970 297978
rect 97026 297922 97094 297978
rect 97150 297922 97218 297978
rect 97274 297922 97342 297978
rect 97398 297922 114970 297978
rect 115026 297922 115094 297978
rect 115150 297922 115218 297978
rect 115274 297922 115342 297978
rect 115398 297922 132970 297978
rect 133026 297922 133094 297978
rect 133150 297922 133218 297978
rect 133274 297922 133342 297978
rect 133398 297922 150970 297978
rect 151026 297922 151094 297978
rect 151150 297922 151218 297978
rect 151274 297922 151342 297978
rect 151398 297922 168970 297978
rect 169026 297922 169094 297978
rect 169150 297922 169218 297978
rect 169274 297922 169342 297978
rect 169398 297922 186970 297978
rect 187026 297922 187094 297978
rect 187150 297922 187218 297978
rect 187274 297922 187342 297978
rect 187398 297922 219878 297978
rect 219934 297922 220002 297978
rect 220058 297922 250598 297978
rect 250654 297922 250722 297978
rect 250778 297922 281318 297978
rect 281374 297922 281442 297978
rect 281498 297922 312038 297978
rect 312094 297922 312162 297978
rect 312218 297922 342758 297978
rect 342814 297922 342882 297978
rect 342938 297922 373478 297978
rect 373534 297922 373602 297978
rect 373658 297922 404198 297978
rect 404254 297922 404322 297978
rect 404378 297922 434918 297978
rect 434974 297922 435042 297978
rect 435098 297922 465638 297978
rect 465694 297922 465762 297978
rect 465818 297922 496358 297978
rect 496414 297922 496482 297978
rect 496538 297922 510970 297978
rect 511026 297922 511094 297978
rect 511150 297922 511218 297978
rect 511274 297922 511342 297978
rect 511398 297922 528970 297978
rect 529026 297922 529094 297978
rect 529150 297922 529218 297978
rect 529274 297922 529342 297978
rect 529398 297922 546970 297978
rect 547026 297922 547094 297978
rect 547150 297922 547218 297978
rect 547274 297922 547342 297978
rect 547398 297922 564970 297978
rect 565026 297922 565094 297978
rect 565150 297922 565218 297978
rect 565274 297922 565342 297978
rect 565398 297922 582970 297978
rect 583026 297922 583094 297978
rect 583150 297922 583218 297978
rect 583274 297922 583342 297978
rect 583398 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 3250 292350
rect 3306 292294 3374 292350
rect 3430 292294 3498 292350
rect 3554 292294 3622 292350
rect 3678 292294 21250 292350
rect 21306 292294 21374 292350
rect 21430 292294 21498 292350
rect 21554 292294 21622 292350
rect 21678 292294 39250 292350
rect 39306 292294 39374 292350
rect 39430 292294 39498 292350
rect 39554 292294 39622 292350
rect 39678 292294 57250 292350
rect 57306 292294 57374 292350
rect 57430 292294 57498 292350
rect 57554 292294 57622 292350
rect 57678 292294 75250 292350
rect 75306 292294 75374 292350
rect 75430 292294 75498 292350
rect 75554 292294 75622 292350
rect 75678 292294 93250 292350
rect 93306 292294 93374 292350
rect 93430 292294 93498 292350
rect 93554 292294 93622 292350
rect 93678 292294 111250 292350
rect 111306 292294 111374 292350
rect 111430 292294 111498 292350
rect 111554 292294 111622 292350
rect 111678 292294 129250 292350
rect 129306 292294 129374 292350
rect 129430 292294 129498 292350
rect 129554 292294 129622 292350
rect 129678 292294 147250 292350
rect 147306 292294 147374 292350
rect 147430 292294 147498 292350
rect 147554 292294 147622 292350
rect 147678 292294 165250 292350
rect 165306 292294 165374 292350
rect 165430 292294 165498 292350
rect 165554 292294 165622 292350
rect 165678 292294 183250 292350
rect 183306 292294 183374 292350
rect 183430 292294 183498 292350
rect 183554 292294 183622 292350
rect 183678 292294 201250 292350
rect 201306 292294 201374 292350
rect 201430 292294 201498 292350
rect 201554 292294 201622 292350
rect 201678 292294 204518 292350
rect 204574 292294 204642 292350
rect 204698 292294 235238 292350
rect 235294 292294 235362 292350
rect 235418 292294 265958 292350
rect 266014 292294 266082 292350
rect 266138 292294 296678 292350
rect 296734 292294 296802 292350
rect 296858 292294 327398 292350
rect 327454 292294 327522 292350
rect 327578 292294 358118 292350
rect 358174 292294 358242 292350
rect 358298 292294 388838 292350
rect 388894 292294 388962 292350
rect 389018 292294 419558 292350
rect 419614 292294 419682 292350
rect 419738 292294 450278 292350
rect 450334 292294 450402 292350
rect 450458 292294 480998 292350
rect 481054 292294 481122 292350
rect 481178 292294 507250 292350
rect 507306 292294 507374 292350
rect 507430 292294 507498 292350
rect 507554 292294 507622 292350
rect 507678 292294 525250 292350
rect 525306 292294 525374 292350
rect 525430 292294 525498 292350
rect 525554 292294 525622 292350
rect 525678 292294 543250 292350
rect 543306 292294 543374 292350
rect 543430 292294 543498 292350
rect 543554 292294 543622 292350
rect 543678 292294 561250 292350
rect 561306 292294 561374 292350
rect 561430 292294 561498 292350
rect 561554 292294 561622 292350
rect 561678 292294 579250 292350
rect 579306 292294 579374 292350
rect 579430 292294 579498 292350
rect 579554 292294 579622 292350
rect 579678 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 3250 292226
rect 3306 292170 3374 292226
rect 3430 292170 3498 292226
rect 3554 292170 3622 292226
rect 3678 292170 21250 292226
rect 21306 292170 21374 292226
rect 21430 292170 21498 292226
rect 21554 292170 21622 292226
rect 21678 292170 39250 292226
rect 39306 292170 39374 292226
rect 39430 292170 39498 292226
rect 39554 292170 39622 292226
rect 39678 292170 57250 292226
rect 57306 292170 57374 292226
rect 57430 292170 57498 292226
rect 57554 292170 57622 292226
rect 57678 292170 75250 292226
rect 75306 292170 75374 292226
rect 75430 292170 75498 292226
rect 75554 292170 75622 292226
rect 75678 292170 93250 292226
rect 93306 292170 93374 292226
rect 93430 292170 93498 292226
rect 93554 292170 93622 292226
rect 93678 292170 111250 292226
rect 111306 292170 111374 292226
rect 111430 292170 111498 292226
rect 111554 292170 111622 292226
rect 111678 292170 129250 292226
rect 129306 292170 129374 292226
rect 129430 292170 129498 292226
rect 129554 292170 129622 292226
rect 129678 292170 147250 292226
rect 147306 292170 147374 292226
rect 147430 292170 147498 292226
rect 147554 292170 147622 292226
rect 147678 292170 165250 292226
rect 165306 292170 165374 292226
rect 165430 292170 165498 292226
rect 165554 292170 165622 292226
rect 165678 292170 183250 292226
rect 183306 292170 183374 292226
rect 183430 292170 183498 292226
rect 183554 292170 183622 292226
rect 183678 292170 201250 292226
rect 201306 292170 201374 292226
rect 201430 292170 201498 292226
rect 201554 292170 201622 292226
rect 201678 292170 204518 292226
rect 204574 292170 204642 292226
rect 204698 292170 235238 292226
rect 235294 292170 235362 292226
rect 235418 292170 265958 292226
rect 266014 292170 266082 292226
rect 266138 292170 296678 292226
rect 296734 292170 296802 292226
rect 296858 292170 327398 292226
rect 327454 292170 327522 292226
rect 327578 292170 358118 292226
rect 358174 292170 358242 292226
rect 358298 292170 388838 292226
rect 388894 292170 388962 292226
rect 389018 292170 419558 292226
rect 419614 292170 419682 292226
rect 419738 292170 450278 292226
rect 450334 292170 450402 292226
rect 450458 292170 480998 292226
rect 481054 292170 481122 292226
rect 481178 292170 507250 292226
rect 507306 292170 507374 292226
rect 507430 292170 507498 292226
rect 507554 292170 507622 292226
rect 507678 292170 525250 292226
rect 525306 292170 525374 292226
rect 525430 292170 525498 292226
rect 525554 292170 525622 292226
rect 525678 292170 543250 292226
rect 543306 292170 543374 292226
rect 543430 292170 543498 292226
rect 543554 292170 543622 292226
rect 543678 292170 561250 292226
rect 561306 292170 561374 292226
rect 561430 292170 561498 292226
rect 561554 292170 561622 292226
rect 561678 292170 579250 292226
rect 579306 292170 579374 292226
rect 579430 292170 579498 292226
rect 579554 292170 579622 292226
rect 579678 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 3250 292102
rect 3306 292046 3374 292102
rect 3430 292046 3498 292102
rect 3554 292046 3622 292102
rect 3678 292046 21250 292102
rect 21306 292046 21374 292102
rect 21430 292046 21498 292102
rect 21554 292046 21622 292102
rect 21678 292046 39250 292102
rect 39306 292046 39374 292102
rect 39430 292046 39498 292102
rect 39554 292046 39622 292102
rect 39678 292046 57250 292102
rect 57306 292046 57374 292102
rect 57430 292046 57498 292102
rect 57554 292046 57622 292102
rect 57678 292046 75250 292102
rect 75306 292046 75374 292102
rect 75430 292046 75498 292102
rect 75554 292046 75622 292102
rect 75678 292046 93250 292102
rect 93306 292046 93374 292102
rect 93430 292046 93498 292102
rect 93554 292046 93622 292102
rect 93678 292046 111250 292102
rect 111306 292046 111374 292102
rect 111430 292046 111498 292102
rect 111554 292046 111622 292102
rect 111678 292046 129250 292102
rect 129306 292046 129374 292102
rect 129430 292046 129498 292102
rect 129554 292046 129622 292102
rect 129678 292046 147250 292102
rect 147306 292046 147374 292102
rect 147430 292046 147498 292102
rect 147554 292046 147622 292102
rect 147678 292046 165250 292102
rect 165306 292046 165374 292102
rect 165430 292046 165498 292102
rect 165554 292046 165622 292102
rect 165678 292046 183250 292102
rect 183306 292046 183374 292102
rect 183430 292046 183498 292102
rect 183554 292046 183622 292102
rect 183678 292046 201250 292102
rect 201306 292046 201374 292102
rect 201430 292046 201498 292102
rect 201554 292046 201622 292102
rect 201678 292046 204518 292102
rect 204574 292046 204642 292102
rect 204698 292046 235238 292102
rect 235294 292046 235362 292102
rect 235418 292046 265958 292102
rect 266014 292046 266082 292102
rect 266138 292046 296678 292102
rect 296734 292046 296802 292102
rect 296858 292046 327398 292102
rect 327454 292046 327522 292102
rect 327578 292046 358118 292102
rect 358174 292046 358242 292102
rect 358298 292046 388838 292102
rect 388894 292046 388962 292102
rect 389018 292046 419558 292102
rect 419614 292046 419682 292102
rect 419738 292046 450278 292102
rect 450334 292046 450402 292102
rect 450458 292046 480998 292102
rect 481054 292046 481122 292102
rect 481178 292046 507250 292102
rect 507306 292046 507374 292102
rect 507430 292046 507498 292102
rect 507554 292046 507622 292102
rect 507678 292046 525250 292102
rect 525306 292046 525374 292102
rect 525430 292046 525498 292102
rect 525554 292046 525622 292102
rect 525678 292046 543250 292102
rect 543306 292046 543374 292102
rect 543430 292046 543498 292102
rect 543554 292046 543622 292102
rect 543678 292046 561250 292102
rect 561306 292046 561374 292102
rect 561430 292046 561498 292102
rect 561554 292046 561622 292102
rect 561678 292046 579250 292102
rect 579306 292046 579374 292102
rect 579430 292046 579498 292102
rect 579554 292046 579622 292102
rect 579678 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 3250 291978
rect 3306 291922 3374 291978
rect 3430 291922 3498 291978
rect 3554 291922 3622 291978
rect 3678 291922 21250 291978
rect 21306 291922 21374 291978
rect 21430 291922 21498 291978
rect 21554 291922 21622 291978
rect 21678 291922 39250 291978
rect 39306 291922 39374 291978
rect 39430 291922 39498 291978
rect 39554 291922 39622 291978
rect 39678 291922 57250 291978
rect 57306 291922 57374 291978
rect 57430 291922 57498 291978
rect 57554 291922 57622 291978
rect 57678 291922 75250 291978
rect 75306 291922 75374 291978
rect 75430 291922 75498 291978
rect 75554 291922 75622 291978
rect 75678 291922 93250 291978
rect 93306 291922 93374 291978
rect 93430 291922 93498 291978
rect 93554 291922 93622 291978
rect 93678 291922 111250 291978
rect 111306 291922 111374 291978
rect 111430 291922 111498 291978
rect 111554 291922 111622 291978
rect 111678 291922 129250 291978
rect 129306 291922 129374 291978
rect 129430 291922 129498 291978
rect 129554 291922 129622 291978
rect 129678 291922 147250 291978
rect 147306 291922 147374 291978
rect 147430 291922 147498 291978
rect 147554 291922 147622 291978
rect 147678 291922 165250 291978
rect 165306 291922 165374 291978
rect 165430 291922 165498 291978
rect 165554 291922 165622 291978
rect 165678 291922 183250 291978
rect 183306 291922 183374 291978
rect 183430 291922 183498 291978
rect 183554 291922 183622 291978
rect 183678 291922 201250 291978
rect 201306 291922 201374 291978
rect 201430 291922 201498 291978
rect 201554 291922 201622 291978
rect 201678 291922 204518 291978
rect 204574 291922 204642 291978
rect 204698 291922 235238 291978
rect 235294 291922 235362 291978
rect 235418 291922 265958 291978
rect 266014 291922 266082 291978
rect 266138 291922 296678 291978
rect 296734 291922 296802 291978
rect 296858 291922 327398 291978
rect 327454 291922 327522 291978
rect 327578 291922 358118 291978
rect 358174 291922 358242 291978
rect 358298 291922 388838 291978
rect 388894 291922 388962 291978
rect 389018 291922 419558 291978
rect 419614 291922 419682 291978
rect 419738 291922 450278 291978
rect 450334 291922 450402 291978
rect 450458 291922 480998 291978
rect 481054 291922 481122 291978
rect 481178 291922 507250 291978
rect 507306 291922 507374 291978
rect 507430 291922 507498 291978
rect 507554 291922 507622 291978
rect 507678 291922 525250 291978
rect 525306 291922 525374 291978
rect 525430 291922 525498 291978
rect 525554 291922 525622 291978
rect 525678 291922 543250 291978
rect 543306 291922 543374 291978
rect 543430 291922 543498 291978
rect 543554 291922 543622 291978
rect 543678 291922 561250 291978
rect 561306 291922 561374 291978
rect 561430 291922 561498 291978
rect 561554 291922 561622 291978
rect 561678 291922 579250 291978
rect 579306 291922 579374 291978
rect 579430 291922 579498 291978
rect 579554 291922 579622 291978
rect 579678 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 6970 280350
rect 7026 280294 7094 280350
rect 7150 280294 7218 280350
rect 7274 280294 7342 280350
rect 7398 280294 24970 280350
rect 25026 280294 25094 280350
rect 25150 280294 25218 280350
rect 25274 280294 25342 280350
rect 25398 280294 42970 280350
rect 43026 280294 43094 280350
rect 43150 280294 43218 280350
rect 43274 280294 43342 280350
rect 43398 280294 60970 280350
rect 61026 280294 61094 280350
rect 61150 280294 61218 280350
rect 61274 280294 61342 280350
rect 61398 280294 78970 280350
rect 79026 280294 79094 280350
rect 79150 280294 79218 280350
rect 79274 280294 79342 280350
rect 79398 280294 96970 280350
rect 97026 280294 97094 280350
rect 97150 280294 97218 280350
rect 97274 280294 97342 280350
rect 97398 280294 114970 280350
rect 115026 280294 115094 280350
rect 115150 280294 115218 280350
rect 115274 280294 115342 280350
rect 115398 280294 132970 280350
rect 133026 280294 133094 280350
rect 133150 280294 133218 280350
rect 133274 280294 133342 280350
rect 133398 280294 150970 280350
rect 151026 280294 151094 280350
rect 151150 280294 151218 280350
rect 151274 280294 151342 280350
rect 151398 280294 168970 280350
rect 169026 280294 169094 280350
rect 169150 280294 169218 280350
rect 169274 280294 169342 280350
rect 169398 280294 186970 280350
rect 187026 280294 187094 280350
rect 187150 280294 187218 280350
rect 187274 280294 187342 280350
rect 187398 280294 219878 280350
rect 219934 280294 220002 280350
rect 220058 280294 250598 280350
rect 250654 280294 250722 280350
rect 250778 280294 281318 280350
rect 281374 280294 281442 280350
rect 281498 280294 312038 280350
rect 312094 280294 312162 280350
rect 312218 280294 342758 280350
rect 342814 280294 342882 280350
rect 342938 280294 373478 280350
rect 373534 280294 373602 280350
rect 373658 280294 404198 280350
rect 404254 280294 404322 280350
rect 404378 280294 434918 280350
rect 434974 280294 435042 280350
rect 435098 280294 465638 280350
rect 465694 280294 465762 280350
rect 465818 280294 496358 280350
rect 496414 280294 496482 280350
rect 496538 280294 510970 280350
rect 511026 280294 511094 280350
rect 511150 280294 511218 280350
rect 511274 280294 511342 280350
rect 511398 280294 528970 280350
rect 529026 280294 529094 280350
rect 529150 280294 529218 280350
rect 529274 280294 529342 280350
rect 529398 280294 546970 280350
rect 547026 280294 547094 280350
rect 547150 280294 547218 280350
rect 547274 280294 547342 280350
rect 547398 280294 564970 280350
rect 565026 280294 565094 280350
rect 565150 280294 565218 280350
rect 565274 280294 565342 280350
rect 565398 280294 582970 280350
rect 583026 280294 583094 280350
rect 583150 280294 583218 280350
rect 583274 280294 583342 280350
rect 583398 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 6970 280226
rect 7026 280170 7094 280226
rect 7150 280170 7218 280226
rect 7274 280170 7342 280226
rect 7398 280170 24970 280226
rect 25026 280170 25094 280226
rect 25150 280170 25218 280226
rect 25274 280170 25342 280226
rect 25398 280170 42970 280226
rect 43026 280170 43094 280226
rect 43150 280170 43218 280226
rect 43274 280170 43342 280226
rect 43398 280170 60970 280226
rect 61026 280170 61094 280226
rect 61150 280170 61218 280226
rect 61274 280170 61342 280226
rect 61398 280170 78970 280226
rect 79026 280170 79094 280226
rect 79150 280170 79218 280226
rect 79274 280170 79342 280226
rect 79398 280170 96970 280226
rect 97026 280170 97094 280226
rect 97150 280170 97218 280226
rect 97274 280170 97342 280226
rect 97398 280170 114970 280226
rect 115026 280170 115094 280226
rect 115150 280170 115218 280226
rect 115274 280170 115342 280226
rect 115398 280170 132970 280226
rect 133026 280170 133094 280226
rect 133150 280170 133218 280226
rect 133274 280170 133342 280226
rect 133398 280170 150970 280226
rect 151026 280170 151094 280226
rect 151150 280170 151218 280226
rect 151274 280170 151342 280226
rect 151398 280170 168970 280226
rect 169026 280170 169094 280226
rect 169150 280170 169218 280226
rect 169274 280170 169342 280226
rect 169398 280170 186970 280226
rect 187026 280170 187094 280226
rect 187150 280170 187218 280226
rect 187274 280170 187342 280226
rect 187398 280170 219878 280226
rect 219934 280170 220002 280226
rect 220058 280170 250598 280226
rect 250654 280170 250722 280226
rect 250778 280170 281318 280226
rect 281374 280170 281442 280226
rect 281498 280170 312038 280226
rect 312094 280170 312162 280226
rect 312218 280170 342758 280226
rect 342814 280170 342882 280226
rect 342938 280170 373478 280226
rect 373534 280170 373602 280226
rect 373658 280170 404198 280226
rect 404254 280170 404322 280226
rect 404378 280170 434918 280226
rect 434974 280170 435042 280226
rect 435098 280170 465638 280226
rect 465694 280170 465762 280226
rect 465818 280170 496358 280226
rect 496414 280170 496482 280226
rect 496538 280170 510970 280226
rect 511026 280170 511094 280226
rect 511150 280170 511218 280226
rect 511274 280170 511342 280226
rect 511398 280170 528970 280226
rect 529026 280170 529094 280226
rect 529150 280170 529218 280226
rect 529274 280170 529342 280226
rect 529398 280170 546970 280226
rect 547026 280170 547094 280226
rect 547150 280170 547218 280226
rect 547274 280170 547342 280226
rect 547398 280170 564970 280226
rect 565026 280170 565094 280226
rect 565150 280170 565218 280226
rect 565274 280170 565342 280226
rect 565398 280170 582970 280226
rect 583026 280170 583094 280226
rect 583150 280170 583218 280226
rect 583274 280170 583342 280226
rect 583398 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 6970 280102
rect 7026 280046 7094 280102
rect 7150 280046 7218 280102
rect 7274 280046 7342 280102
rect 7398 280046 24970 280102
rect 25026 280046 25094 280102
rect 25150 280046 25218 280102
rect 25274 280046 25342 280102
rect 25398 280046 42970 280102
rect 43026 280046 43094 280102
rect 43150 280046 43218 280102
rect 43274 280046 43342 280102
rect 43398 280046 60970 280102
rect 61026 280046 61094 280102
rect 61150 280046 61218 280102
rect 61274 280046 61342 280102
rect 61398 280046 78970 280102
rect 79026 280046 79094 280102
rect 79150 280046 79218 280102
rect 79274 280046 79342 280102
rect 79398 280046 96970 280102
rect 97026 280046 97094 280102
rect 97150 280046 97218 280102
rect 97274 280046 97342 280102
rect 97398 280046 114970 280102
rect 115026 280046 115094 280102
rect 115150 280046 115218 280102
rect 115274 280046 115342 280102
rect 115398 280046 132970 280102
rect 133026 280046 133094 280102
rect 133150 280046 133218 280102
rect 133274 280046 133342 280102
rect 133398 280046 150970 280102
rect 151026 280046 151094 280102
rect 151150 280046 151218 280102
rect 151274 280046 151342 280102
rect 151398 280046 168970 280102
rect 169026 280046 169094 280102
rect 169150 280046 169218 280102
rect 169274 280046 169342 280102
rect 169398 280046 186970 280102
rect 187026 280046 187094 280102
rect 187150 280046 187218 280102
rect 187274 280046 187342 280102
rect 187398 280046 219878 280102
rect 219934 280046 220002 280102
rect 220058 280046 250598 280102
rect 250654 280046 250722 280102
rect 250778 280046 281318 280102
rect 281374 280046 281442 280102
rect 281498 280046 312038 280102
rect 312094 280046 312162 280102
rect 312218 280046 342758 280102
rect 342814 280046 342882 280102
rect 342938 280046 373478 280102
rect 373534 280046 373602 280102
rect 373658 280046 404198 280102
rect 404254 280046 404322 280102
rect 404378 280046 434918 280102
rect 434974 280046 435042 280102
rect 435098 280046 465638 280102
rect 465694 280046 465762 280102
rect 465818 280046 496358 280102
rect 496414 280046 496482 280102
rect 496538 280046 510970 280102
rect 511026 280046 511094 280102
rect 511150 280046 511218 280102
rect 511274 280046 511342 280102
rect 511398 280046 528970 280102
rect 529026 280046 529094 280102
rect 529150 280046 529218 280102
rect 529274 280046 529342 280102
rect 529398 280046 546970 280102
rect 547026 280046 547094 280102
rect 547150 280046 547218 280102
rect 547274 280046 547342 280102
rect 547398 280046 564970 280102
rect 565026 280046 565094 280102
rect 565150 280046 565218 280102
rect 565274 280046 565342 280102
rect 565398 280046 582970 280102
rect 583026 280046 583094 280102
rect 583150 280046 583218 280102
rect 583274 280046 583342 280102
rect 583398 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 6970 279978
rect 7026 279922 7094 279978
rect 7150 279922 7218 279978
rect 7274 279922 7342 279978
rect 7398 279922 24970 279978
rect 25026 279922 25094 279978
rect 25150 279922 25218 279978
rect 25274 279922 25342 279978
rect 25398 279922 42970 279978
rect 43026 279922 43094 279978
rect 43150 279922 43218 279978
rect 43274 279922 43342 279978
rect 43398 279922 60970 279978
rect 61026 279922 61094 279978
rect 61150 279922 61218 279978
rect 61274 279922 61342 279978
rect 61398 279922 78970 279978
rect 79026 279922 79094 279978
rect 79150 279922 79218 279978
rect 79274 279922 79342 279978
rect 79398 279922 96970 279978
rect 97026 279922 97094 279978
rect 97150 279922 97218 279978
rect 97274 279922 97342 279978
rect 97398 279922 114970 279978
rect 115026 279922 115094 279978
rect 115150 279922 115218 279978
rect 115274 279922 115342 279978
rect 115398 279922 132970 279978
rect 133026 279922 133094 279978
rect 133150 279922 133218 279978
rect 133274 279922 133342 279978
rect 133398 279922 150970 279978
rect 151026 279922 151094 279978
rect 151150 279922 151218 279978
rect 151274 279922 151342 279978
rect 151398 279922 168970 279978
rect 169026 279922 169094 279978
rect 169150 279922 169218 279978
rect 169274 279922 169342 279978
rect 169398 279922 186970 279978
rect 187026 279922 187094 279978
rect 187150 279922 187218 279978
rect 187274 279922 187342 279978
rect 187398 279922 219878 279978
rect 219934 279922 220002 279978
rect 220058 279922 250598 279978
rect 250654 279922 250722 279978
rect 250778 279922 281318 279978
rect 281374 279922 281442 279978
rect 281498 279922 312038 279978
rect 312094 279922 312162 279978
rect 312218 279922 342758 279978
rect 342814 279922 342882 279978
rect 342938 279922 373478 279978
rect 373534 279922 373602 279978
rect 373658 279922 404198 279978
rect 404254 279922 404322 279978
rect 404378 279922 434918 279978
rect 434974 279922 435042 279978
rect 435098 279922 465638 279978
rect 465694 279922 465762 279978
rect 465818 279922 496358 279978
rect 496414 279922 496482 279978
rect 496538 279922 510970 279978
rect 511026 279922 511094 279978
rect 511150 279922 511218 279978
rect 511274 279922 511342 279978
rect 511398 279922 528970 279978
rect 529026 279922 529094 279978
rect 529150 279922 529218 279978
rect 529274 279922 529342 279978
rect 529398 279922 546970 279978
rect 547026 279922 547094 279978
rect 547150 279922 547218 279978
rect 547274 279922 547342 279978
rect 547398 279922 564970 279978
rect 565026 279922 565094 279978
rect 565150 279922 565218 279978
rect 565274 279922 565342 279978
rect 565398 279922 582970 279978
rect 583026 279922 583094 279978
rect 583150 279922 583218 279978
rect 583274 279922 583342 279978
rect 583398 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 3250 274350
rect 3306 274294 3374 274350
rect 3430 274294 3498 274350
rect 3554 274294 3622 274350
rect 3678 274294 21250 274350
rect 21306 274294 21374 274350
rect 21430 274294 21498 274350
rect 21554 274294 21622 274350
rect 21678 274294 39250 274350
rect 39306 274294 39374 274350
rect 39430 274294 39498 274350
rect 39554 274294 39622 274350
rect 39678 274294 57250 274350
rect 57306 274294 57374 274350
rect 57430 274294 57498 274350
rect 57554 274294 57622 274350
rect 57678 274294 75250 274350
rect 75306 274294 75374 274350
rect 75430 274294 75498 274350
rect 75554 274294 75622 274350
rect 75678 274294 93250 274350
rect 93306 274294 93374 274350
rect 93430 274294 93498 274350
rect 93554 274294 93622 274350
rect 93678 274294 111250 274350
rect 111306 274294 111374 274350
rect 111430 274294 111498 274350
rect 111554 274294 111622 274350
rect 111678 274294 129250 274350
rect 129306 274294 129374 274350
rect 129430 274294 129498 274350
rect 129554 274294 129622 274350
rect 129678 274294 147250 274350
rect 147306 274294 147374 274350
rect 147430 274294 147498 274350
rect 147554 274294 147622 274350
rect 147678 274294 165250 274350
rect 165306 274294 165374 274350
rect 165430 274294 165498 274350
rect 165554 274294 165622 274350
rect 165678 274294 183250 274350
rect 183306 274294 183374 274350
rect 183430 274294 183498 274350
rect 183554 274294 183622 274350
rect 183678 274294 201250 274350
rect 201306 274294 201374 274350
rect 201430 274294 201498 274350
rect 201554 274294 201622 274350
rect 201678 274294 204518 274350
rect 204574 274294 204642 274350
rect 204698 274294 235238 274350
rect 235294 274294 235362 274350
rect 235418 274294 265958 274350
rect 266014 274294 266082 274350
rect 266138 274294 296678 274350
rect 296734 274294 296802 274350
rect 296858 274294 327398 274350
rect 327454 274294 327522 274350
rect 327578 274294 358118 274350
rect 358174 274294 358242 274350
rect 358298 274294 388838 274350
rect 388894 274294 388962 274350
rect 389018 274294 419558 274350
rect 419614 274294 419682 274350
rect 419738 274294 450278 274350
rect 450334 274294 450402 274350
rect 450458 274294 480998 274350
rect 481054 274294 481122 274350
rect 481178 274294 507250 274350
rect 507306 274294 507374 274350
rect 507430 274294 507498 274350
rect 507554 274294 507622 274350
rect 507678 274294 525250 274350
rect 525306 274294 525374 274350
rect 525430 274294 525498 274350
rect 525554 274294 525622 274350
rect 525678 274294 543250 274350
rect 543306 274294 543374 274350
rect 543430 274294 543498 274350
rect 543554 274294 543622 274350
rect 543678 274294 561250 274350
rect 561306 274294 561374 274350
rect 561430 274294 561498 274350
rect 561554 274294 561622 274350
rect 561678 274294 579250 274350
rect 579306 274294 579374 274350
rect 579430 274294 579498 274350
rect 579554 274294 579622 274350
rect 579678 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 3250 274226
rect 3306 274170 3374 274226
rect 3430 274170 3498 274226
rect 3554 274170 3622 274226
rect 3678 274170 21250 274226
rect 21306 274170 21374 274226
rect 21430 274170 21498 274226
rect 21554 274170 21622 274226
rect 21678 274170 39250 274226
rect 39306 274170 39374 274226
rect 39430 274170 39498 274226
rect 39554 274170 39622 274226
rect 39678 274170 57250 274226
rect 57306 274170 57374 274226
rect 57430 274170 57498 274226
rect 57554 274170 57622 274226
rect 57678 274170 75250 274226
rect 75306 274170 75374 274226
rect 75430 274170 75498 274226
rect 75554 274170 75622 274226
rect 75678 274170 93250 274226
rect 93306 274170 93374 274226
rect 93430 274170 93498 274226
rect 93554 274170 93622 274226
rect 93678 274170 111250 274226
rect 111306 274170 111374 274226
rect 111430 274170 111498 274226
rect 111554 274170 111622 274226
rect 111678 274170 129250 274226
rect 129306 274170 129374 274226
rect 129430 274170 129498 274226
rect 129554 274170 129622 274226
rect 129678 274170 147250 274226
rect 147306 274170 147374 274226
rect 147430 274170 147498 274226
rect 147554 274170 147622 274226
rect 147678 274170 165250 274226
rect 165306 274170 165374 274226
rect 165430 274170 165498 274226
rect 165554 274170 165622 274226
rect 165678 274170 183250 274226
rect 183306 274170 183374 274226
rect 183430 274170 183498 274226
rect 183554 274170 183622 274226
rect 183678 274170 201250 274226
rect 201306 274170 201374 274226
rect 201430 274170 201498 274226
rect 201554 274170 201622 274226
rect 201678 274170 204518 274226
rect 204574 274170 204642 274226
rect 204698 274170 235238 274226
rect 235294 274170 235362 274226
rect 235418 274170 265958 274226
rect 266014 274170 266082 274226
rect 266138 274170 296678 274226
rect 296734 274170 296802 274226
rect 296858 274170 327398 274226
rect 327454 274170 327522 274226
rect 327578 274170 358118 274226
rect 358174 274170 358242 274226
rect 358298 274170 388838 274226
rect 388894 274170 388962 274226
rect 389018 274170 419558 274226
rect 419614 274170 419682 274226
rect 419738 274170 450278 274226
rect 450334 274170 450402 274226
rect 450458 274170 480998 274226
rect 481054 274170 481122 274226
rect 481178 274170 507250 274226
rect 507306 274170 507374 274226
rect 507430 274170 507498 274226
rect 507554 274170 507622 274226
rect 507678 274170 525250 274226
rect 525306 274170 525374 274226
rect 525430 274170 525498 274226
rect 525554 274170 525622 274226
rect 525678 274170 543250 274226
rect 543306 274170 543374 274226
rect 543430 274170 543498 274226
rect 543554 274170 543622 274226
rect 543678 274170 561250 274226
rect 561306 274170 561374 274226
rect 561430 274170 561498 274226
rect 561554 274170 561622 274226
rect 561678 274170 579250 274226
rect 579306 274170 579374 274226
rect 579430 274170 579498 274226
rect 579554 274170 579622 274226
rect 579678 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 3250 274102
rect 3306 274046 3374 274102
rect 3430 274046 3498 274102
rect 3554 274046 3622 274102
rect 3678 274046 21250 274102
rect 21306 274046 21374 274102
rect 21430 274046 21498 274102
rect 21554 274046 21622 274102
rect 21678 274046 39250 274102
rect 39306 274046 39374 274102
rect 39430 274046 39498 274102
rect 39554 274046 39622 274102
rect 39678 274046 57250 274102
rect 57306 274046 57374 274102
rect 57430 274046 57498 274102
rect 57554 274046 57622 274102
rect 57678 274046 75250 274102
rect 75306 274046 75374 274102
rect 75430 274046 75498 274102
rect 75554 274046 75622 274102
rect 75678 274046 93250 274102
rect 93306 274046 93374 274102
rect 93430 274046 93498 274102
rect 93554 274046 93622 274102
rect 93678 274046 111250 274102
rect 111306 274046 111374 274102
rect 111430 274046 111498 274102
rect 111554 274046 111622 274102
rect 111678 274046 129250 274102
rect 129306 274046 129374 274102
rect 129430 274046 129498 274102
rect 129554 274046 129622 274102
rect 129678 274046 147250 274102
rect 147306 274046 147374 274102
rect 147430 274046 147498 274102
rect 147554 274046 147622 274102
rect 147678 274046 165250 274102
rect 165306 274046 165374 274102
rect 165430 274046 165498 274102
rect 165554 274046 165622 274102
rect 165678 274046 183250 274102
rect 183306 274046 183374 274102
rect 183430 274046 183498 274102
rect 183554 274046 183622 274102
rect 183678 274046 201250 274102
rect 201306 274046 201374 274102
rect 201430 274046 201498 274102
rect 201554 274046 201622 274102
rect 201678 274046 204518 274102
rect 204574 274046 204642 274102
rect 204698 274046 235238 274102
rect 235294 274046 235362 274102
rect 235418 274046 265958 274102
rect 266014 274046 266082 274102
rect 266138 274046 296678 274102
rect 296734 274046 296802 274102
rect 296858 274046 327398 274102
rect 327454 274046 327522 274102
rect 327578 274046 358118 274102
rect 358174 274046 358242 274102
rect 358298 274046 388838 274102
rect 388894 274046 388962 274102
rect 389018 274046 419558 274102
rect 419614 274046 419682 274102
rect 419738 274046 450278 274102
rect 450334 274046 450402 274102
rect 450458 274046 480998 274102
rect 481054 274046 481122 274102
rect 481178 274046 507250 274102
rect 507306 274046 507374 274102
rect 507430 274046 507498 274102
rect 507554 274046 507622 274102
rect 507678 274046 525250 274102
rect 525306 274046 525374 274102
rect 525430 274046 525498 274102
rect 525554 274046 525622 274102
rect 525678 274046 543250 274102
rect 543306 274046 543374 274102
rect 543430 274046 543498 274102
rect 543554 274046 543622 274102
rect 543678 274046 561250 274102
rect 561306 274046 561374 274102
rect 561430 274046 561498 274102
rect 561554 274046 561622 274102
rect 561678 274046 579250 274102
rect 579306 274046 579374 274102
rect 579430 274046 579498 274102
rect 579554 274046 579622 274102
rect 579678 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 3250 273978
rect 3306 273922 3374 273978
rect 3430 273922 3498 273978
rect 3554 273922 3622 273978
rect 3678 273922 21250 273978
rect 21306 273922 21374 273978
rect 21430 273922 21498 273978
rect 21554 273922 21622 273978
rect 21678 273922 39250 273978
rect 39306 273922 39374 273978
rect 39430 273922 39498 273978
rect 39554 273922 39622 273978
rect 39678 273922 57250 273978
rect 57306 273922 57374 273978
rect 57430 273922 57498 273978
rect 57554 273922 57622 273978
rect 57678 273922 75250 273978
rect 75306 273922 75374 273978
rect 75430 273922 75498 273978
rect 75554 273922 75622 273978
rect 75678 273922 93250 273978
rect 93306 273922 93374 273978
rect 93430 273922 93498 273978
rect 93554 273922 93622 273978
rect 93678 273922 111250 273978
rect 111306 273922 111374 273978
rect 111430 273922 111498 273978
rect 111554 273922 111622 273978
rect 111678 273922 129250 273978
rect 129306 273922 129374 273978
rect 129430 273922 129498 273978
rect 129554 273922 129622 273978
rect 129678 273922 147250 273978
rect 147306 273922 147374 273978
rect 147430 273922 147498 273978
rect 147554 273922 147622 273978
rect 147678 273922 165250 273978
rect 165306 273922 165374 273978
rect 165430 273922 165498 273978
rect 165554 273922 165622 273978
rect 165678 273922 183250 273978
rect 183306 273922 183374 273978
rect 183430 273922 183498 273978
rect 183554 273922 183622 273978
rect 183678 273922 201250 273978
rect 201306 273922 201374 273978
rect 201430 273922 201498 273978
rect 201554 273922 201622 273978
rect 201678 273922 204518 273978
rect 204574 273922 204642 273978
rect 204698 273922 235238 273978
rect 235294 273922 235362 273978
rect 235418 273922 265958 273978
rect 266014 273922 266082 273978
rect 266138 273922 296678 273978
rect 296734 273922 296802 273978
rect 296858 273922 327398 273978
rect 327454 273922 327522 273978
rect 327578 273922 358118 273978
rect 358174 273922 358242 273978
rect 358298 273922 388838 273978
rect 388894 273922 388962 273978
rect 389018 273922 419558 273978
rect 419614 273922 419682 273978
rect 419738 273922 450278 273978
rect 450334 273922 450402 273978
rect 450458 273922 480998 273978
rect 481054 273922 481122 273978
rect 481178 273922 507250 273978
rect 507306 273922 507374 273978
rect 507430 273922 507498 273978
rect 507554 273922 507622 273978
rect 507678 273922 525250 273978
rect 525306 273922 525374 273978
rect 525430 273922 525498 273978
rect 525554 273922 525622 273978
rect 525678 273922 543250 273978
rect 543306 273922 543374 273978
rect 543430 273922 543498 273978
rect 543554 273922 543622 273978
rect 543678 273922 561250 273978
rect 561306 273922 561374 273978
rect 561430 273922 561498 273978
rect 561554 273922 561622 273978
rect 561678 273922 579250 273978
rect 579306 273922 579374 273978
rect 579430 273922 579498 273978
rect 579554 273922 579622 273978
rect 579678 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 6970 262350
rect 7026 262294 7094 262350
rect 7150 262294 7218 262350
rect 7274 262294 7342 262350
rect 7398 262294 24970 262350
rect 25026 262294 25094 262350
rect 25150 262294 25218 262350
rect 25274 262294 25342 262350
rect 25398 262294 42970 262350
rect 43026 262294 43094 262350
rect 43150 262294 43218 262350
rect 43274 262294 43342 262350
rect 43398 262294 60970 262350
rect 61026 262294 61094 262350
rect 61150 262294 61218 262350
rect 61274 262294 61342 262350
rect 61398 262294 78970 262350
rect 79026 262294 79094 262350
rect 79150 262294 79218 262350
rect 79274 262294 79342 262350
rect 79398 262294 96970 262350
rect 97026 262294 97094 262350
rect 97150 262294 97218 262350
rect 97274 262294 97342 262350
rect 97398 262294 114970 262350
rect 115026 262294 115094 262350
rect 115150 262294 115218 262350
rect 115274 262294 115342 262350
rect 115398 262294 132970 262350
rect 133026 262294 133094 262350
rect 133150 262294 133218 262350
rect 133274 262294 133342 262350
rect 133398 262294 150970 262350
rect 151026 262294 151094 262350
rect 151150 262294 151218 262350
rect 151274 262294 151342 262350
rect 151398 262294 168970 262350
rect 169026 262294 169094 262350
rect 169150 262294 169218 262350
rect 169274 262294 169342 262350
rect 169398 262294 186970 262350
rect 187026 262294 187094 262350
rect 187150 262294 187218 262350
rect 187274 262294 187342 262350
rect 187398 262294 219878 262350
rect 219934 262294 220002 262350
rect 220058 262294 250598 262350
rect 250654 262294 250722 262350
rect 250778 262294 281318 262350
rect 281374 262294 281442 262350
rect 281498 262294 312038 262350
rect 312094 262294 312162 262350
rect 312218 262294 342758 262350
rect 342814 262294 342882 262350
rect 342938 262294 373478 262350
rect 373534 262294 373602 262350
rect 373658 262294 404198 262350
rect 404254 262294 404322 262350
rect 404378 262294 434918 262350
rect 434974 262294 435042 262350
rect 435098 262294 465638 262350
rect 465694 262294 465762 262350
rect 465818 262294 496358 262350
rect 496414 262294 496482 262350
rect 496538 262294 510970 262350
rect 511026 262294 511094 262350
rect 511150 262294 511218 262350
rect 511274 262294 511342 262350
rect 511398 262294 528970 262350
rect 529026 262294 529094 262350
rect 529150 262294 529218 262350
rect 529274 262294 529342 262350
rect 529398 262294 546970 262350
rect 547026 262294 547094 262350
rect 547150 262294 547218 262350
rect 547274 262294 547342 262350
rect 547398 262294 564970 262350
rect 565026 262294 565094 262350
rect 565150 262294 565218 262350
rect 565274 262294 565342 262350
rect 565398 262294 582970 262350
rect 583026 262294 583094 262350
rect 583150 262294 583218 262350
rect 583274 262294 583342 262350
rect 583398 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 6970 262226
rect 7026 262170 7094 262226
rect 7150 262170 7218 262226
rect 7274 262170 7342 262226
rect 7398 262170 24970 262226
rect 25026 262170 25094 262226
rect 25150 262170 25218 262226
rect 25274 262170 25342 262226
rect 25398 262170 42970 262226
rect 43026 262170 43094 262226
rect 43150 262170 43218 262226
rect 43274 262170 43342 262226
rect 43398 262170 60970 262226
rect 61026 262170 61094 262226
rect 61150 262170 61218 262226
rect 61274 262170 61342 262226
rect 61398 262170 78970 262226
rect 79026 262170 79094 262226
rect 79150 262170 79218 262226
rect 79274 262170 79342 262226
rect 79398 262170 96970 262226
rect 97026 262170 97094 262226
rect 97150 262170 97218 262226
rect 97274 262170 97342 262226
rect 97398 262170 114970 262226
rect 115026 262170 115094 262226
rect 115150 262170 115218 262226
rect 115274 262170 115342 262226
rect 115398 262170 132970 262226
rect 133026 262170 133094 262226
rect 133150 262170 133218 262226
rect 133274 262170 133342 262226
rect 133398 262170 150970 262226
rect 151026 262170 151094 262226
rect 151150 262170 151218 262226
rect 151274 262170 151342 262226
rect 151398 262170 168970 262226
rect 169026 262170 169094 262226
rect 169150 262170 169218 262226
rect 169274 262170 169342 262226
rect 169398 262170 186970 262226
rect 187026 262170 187094 262226
rect 187150 262170 187218 262226
rect 187274 262170 187342 262226
rect 187398 262170 219878 262226
rect 219934 262170 220002 262226
rect 220058 262170 250598 262226
rect 250654 262170 250722 262226
rect 250778 262170 281318 262226
rect 281374 262170 281442 262226
rect 281498 262170 312038 262226
rect 312094 262170 312162 262226
rect 312218 262170 342758 262226
rect 342814 262170 342882 262226
rect 342938 262170 373478 262226
rect 373534 262170 373602 262226
rect 373658 262170 404198 262226
rect 404254 262170 404322 262226
rect 404378 262170 434918 262226
rect 434974 262170 435042 262226
rect 435098 262170 465638 262226
rect 465694 262170 465762 262226
rect 465818 262170 496358 262226
rect 496414 262170 496482 262226
rect 496538 262170 510970 262226
rect 511026 262170 511094 262226
rect 511150 262170 511218 262226
rect 511274 262170 511342 262226
rect 511398 262170 528970 262226
rect 529026 262170 529094 262226
rect 529150 262170 529218 262226
rect 529274 262170 529342 262226
rect 529398 262170 546970 262226
rect 547026 262170 547094 262226
rect 547150 262170 547218 262226
rect 547274 262170 547342 262226
rect 547398 262170 564970 262226
rect 565026 262170 565094 262226
rect 565150 262170 565218 262226
rect 565274 262170 565342 262226
rect 565398 262170 582970 262226
rect 583026 262170 583094 262226
rect 583150 262170 583218 262226
rect 583274 262170 583342 262226
rect 583398 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 6970 262102
rect 7026 262046 7094 262102
rect 7150 262046 7218 262102
rect 7274 262046 7342 262102
rect 7398 262046 24970 262102
rect 25026 262046 25094 262102
rect 25150 262046 25218 262102
rect 25274 262046 25342 262102
rect 25398 262046 42970 262102
rect 43026 262046 43094 262102
rect 43150 262046 43218 262102
rect 43274 262046 43342 262102
rect 43398 262046 60970 262102
rect 61026 262046 61094 262102
rect 61150 262046 61218 262102
rect 61274 262046 61342 262102
rect 61398 262046 78970 262102
rect 79026 262046 79094 262102
rect 79150 262046 79218 262102
rect 79274 262046 79342 262102
rect 79398 262046 96970 262102
rect 97026 262046 97094 262102
rect 97150 262046 97218 262102
rect 97274 262046 97342 262102
rect 97398 262046 114970 262102
rect 115026 262046 115094 262102
rect 115150 262046 115218 262102
rect 115274 262046 115342 262102
rect 115398 262046 132970 262102
rect 133026 262046 133094 262102
rect 133150 262046 133218 262102
rect 133274 262046 133342 262102
rect 133398 262046 150970 262102
rect 151026 262046 151094 262102
rect 151150 262046 151218 262102
rect 151274 262046 151342 262102
rect 151398 262046 168970 262102
rect 169026 262046 169094 262102
rect 169150 262046 169218 262102
rect 169274 262046 169342 262102
rect 169398 262046 186970 262102
rect 187026 262046 187094 262102
rect 187150 262046 187218 262102
rect 187274 262046 187342 262102
rect 187398 262046 219878 262102
rect 219934 262046 220002 262102
rect 220058 262046 250598 262102
rect 250654 262046 250722 262102
rect 250778 262046 281318 262102
rect 281374 262046 281442 262102
rect 281498 262046 312038 262102
rect 312094 262046 312162 262102
rect 312218 262046 342758 262102
rect 342814 262046 342882 262102
rect 342938 262046 373478 262102
rect 373534 262046 373602 262102
rect 373658 262046 404198 262102
rect 404254 262046 404322 262102
rect 404378 262046 434918 262102
rect 434974 262046 435042 262102
rect 435098 262046 465638 262102
rect 465694 262046 465762 262102
rect 465818 262046 496358 262102
rect 496414 262046 496482 262102
rect 496538 262046 510970 262102
rect 511026 262046 511094 262102
rect 511150 262046 511218 262102
rect 511274 262046 511342 262102
rect 511398 262046 528970 262102
rect 529026 262046 529094 262102
rect 529150 262046 529218 262102
rect 529274 262046 529342 262102
rect 529398 262046 546970 262102
rect 547026 262046 547094 262102
rect 547150 262046 547218 262102
rect 547274 262046 547342 262102
rect 547398 262046 564970 262102
rect 565026 262046 565094 262102
rect 565150 262046 565218 262102
rect 565274 262046 565342 262102
rect 565398 262046 582970 262102
rect 583026 262046 583094 262102
rect 583150 262046 583218 262102
rect 583274 262046 583342 262102
rect 583398 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 6970 261978
rect 7026 261922 7094 261978
rect 7150 261922 7218 261978
rect 7274 261922 7342 261978
rect 7398 261922 24970 261978
rect 25026 261922 25094 261978
rect 25150 261922 25218 261978
rect 25274 261922 25342 261978
rect 25398 261922 42970 261978
rect 43026 261922 43094 261978
rect 43150 261922 43218 261978
rect 43274 261922 43342 261978
rect 43398 261922 60970 261978
rect 61026 261922 61094 261978
rect 61150 261922 61218 261978
rect 61274 261922 61342 261978
rect 61398 261922 78970 261978
rect 79026 261922 79094 261978
rect 79150 261922 79218 261978
rect 79274 261922 79342 261978
rect 79398 261922 96970 261978
rect 97026 261922 97094 261978
rect 97150 261922 97218 261978
rect 97274 261922 97342 261978
rect 97398 261922 114970 261978
rect 115026 261922 115094 261978
rect 115150 261922 115218 261978
rect 115274 261922 115342 261978
rect 115398 261922 132970 261978
rect 133026 261922 133094 261978
rect 133150 261922 133218 261978
rect 133274 261922 133342 261978
rect 133398 261922 150970 261978
rect 151026 261922 151094 261978
rect 151150 261922 151218 261978
rect 151274 261922 151342 261978
rect 151398 261922 168970 261978
rect 169026 261922 169094 261978
rect 169150 261922 169218 261978
rect 169274 261922 169342 261978
rect 169398 261922 186970 261978
rect 187026 261922 187094 261978
rect 187150 261922 187218 261978
rect 187274 261922 187342 261978
rect 187398 261922 219878 261978
rect 219934 261922 220002 261978
rect 220058 261922 250598 261978
rect 250654 261922 250722 261978
rect 250778 261922 281318 261978
rect 281374 261922 281442 261978
rect 281498 261922 312038 261978
rect 312094 261922 312162 261978
rect 312218 261922 342758 261978
rect 342814 261922 342882 261978
rect 342938 261922 373478 261978
rect 373534 261922 373602 261978
rect 373658 261922 404198 261978
rect 404254 261922 404322 261978
rect 404378 261922 434918 261978
rect 434974 261922 435042 261978
rect 435098 261922 465638 261978
rect 465694 261922 465762 261978
rect 465818 261922 496358 261978
rect 496414 261922 496482 261978
rect 496538 261922 510970 261978
rect 511026 261922 511094 261978
rect 511150 261922 511218 261978
rect 511274 261922 511342 261978
rect 511398 261922 528970 261978
rect 529026 261922 529094 261978
rect 529150 261922 529218 261978
rect 529274 261922 529342 261978
rect 529398 261922 546970 261978
rect 547026 261922 547094 261978
rect 547150 261922 547218 261978
rect 547274 261922 547342 261978
rect 547398 261922 564970 261978
rect 565026 261922 565094 261978
rect 565150 261922 565218 261978
rect 565274 261922 565342 261978
rect 565398 261922 582970 261978
rect 583026 261922 583094 261978
rect 583150 261922 583218 261978
rect 583274 261922 583342 261978
rect 583398 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 3250 256350
rect 3306 256294 3374 256350
rect 3430 256294 3498 256350
rect 3554 256294 3622 256350
rect 3678 256294 21250 256350
rect 21306 256294 21374 256350
rect 21430 256294 21498 256350
rect 21554 256294 21622 256350
rect 21678 256294 39250 256350
rect 39306 256294 39374 256350
rect 39430 256294 39498 256350
rect 39554 256294 39622 256350
rect 39678 256294 57250 256350
rect 57306 256294 57374 256350
rect 57430 256294 57498 256350
rect 57554 256294 57622 256350
rect 57678 256294 75250 256350
rect 75306 256294 75374 256350
rect 75430 256294 75498 256350
rect 75554 256294 75622 256350
rect 75678 256294 93250 256350
rect 93306 256294 93374 256350
rect 93430 256294 93498 256350
rect 93554 256294 93622 256350
rect 93678 256294 111250 256350
rect 111306 256294 111374 256350
rect 111430 256294 111498 256350
rect 111554 256294 111622 256350
rect 111678 256294 129250 256350
rect 129306 256294 129374 256350
rect 129430 256294 129498 256350
rect 129554 256294 129622 256350
rect 129678 256294 147250 256350
rect 147306 256294 147374 256350
rect 147430 256294 147498 256350
rect 147554 256294 147622 256350
rect 147678 256294 165250 256350
rect 165306 256294 165374 256350
rect 165430 256294 165498 256350
rect 165554 256294 165622 256350
rect 165678 256294 183250 256350
rect 183306 256294 183374 256350
rect 183430 256294 183498 256350
rect 183554 256294 183622 256350
rect 183678 256294 201250 256350
rect 201306 256294 201374 256350
rect 201430 256294 201498 256350
rect 201554 256294 201622 256350
rect 201678 256294 204518 256350
rect 204574 256294 204642 256350
rect 204698 256294 235238 256350
rect 235294 256294 235362 256350
rect 235418 256294 265958 256350
rect 266014 256294 266082 256350
rect 266138 256294 296678 256350
rect 296734 256294 296802 256350
rect 296858 256294 327398 256350
rect 327454 256294 327522 256350
rect 327578 256294 358118 256350
rect 358174 256294 358242 256350
rect 358298 256294 388838 256350
rect 388894 256294 388962 256350
rect 389018 256294 419558 256350
rect 419614 256294 419682 256350
rect 419738 256294 450278 256350
rect 450334 256294 450402 256350
rect 450458 256294 480998 256350
rect 481054 256294 481122 256350
rect 481178 256294 507250 256350
rect 507306 256294 507374 256350
rect 507430 256294 507498 256350
rect 507554 256294 507622 256350
rect 507678 256294 525250 256350
rect 525306 256294 525374 256350
rect 525430 256294 525498 256350
rect 525554 256294 525622 256350
rect 525678 256294 543250 256350
rect 543306 256294 543374 256350
rect 543430 256294 543498 256350
rect 543554 256294 543622 256350
rect 543678 256294 561250 256350
rect 561306 256294 561374 256350
rect 561430 256294 561498 256350
rect 561554 256294 561622 256350
rect 561678 256294 579250 256350
rect 579306 256294 579374 256350
rect 579430 256294 579498 256350
rect 579554 256294 579622 256350
rect 579678 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 3250 256226
rect 3306 256170 3374 256226
rect 3430 256170 3498 256226
rect 3554 256170 3622 256226
rect 3678 256170 21250 256226
rect 21306 256170 21374 256226
rect 21430 256170 21498 256226
rect 21554 256170 21622 256226
rect 21678 256170 39250 256226
rect 39306 256170 39374 256226
rect 39430 256170 39498 256226
rect 39554 256170 39622 256226
rect 39678 256170 57250 256226
rect 57306 256170 57374 256226
rect 57430 256170 57498 256226
rect 57554 256170 57622 256226
rect 57678 256170 75250 256226
rect 75306 256170 75374 256226
rect 75430 256170 75498 256226
rect 75554 256170 75622 256226
rect 75678 256170 93250 256226
rect 93306 256170 93374 256226
rect 93430 256170 93498 256226
rect 93554 256170 93622 256226
rect 93678 256170 111250 256226
rect 111306 256170 111374 256226
rect 111430 256170 111498 256226
rect 111554 256170 111622 256226
rect 111678 256170 129250 256226
rect 129306 256170 129374 256226
rect 129430 256170 129498 256226
rect 129554 256170 129622 256226
rect 129678 256170 147250 256226
rect 147306 256170 147374 256226
rect 147430 256170 147498 256226
rect 147554 256170 147622 256226
rect 147678 256170 165250 256226
rect 165306 256170 165374 256226
rect 165430 256170 165498 256226
rect 165554 256170 165622 256226
rect 165678 256170 183250 256226
rect 183306 256170 183374 256226
rect 183430 256170 183498 256226
rect 183554 256170 183622 256226
rect 183678 256170 201250 256226
rect 201306 256170 201374 256226
rect 201430 256170 201498 256226
rect 201554 256170 201622 256226
rect 201678 256170 204518 256226
rect 204574 256170 204642 256226
rect 204698 256170 235238 256226
rect 235294 256170 235362 256226
rect 235418 256170 265958 256226
rect 266014 256170 266082 256226
rect 266138 256170 296678 256226
rect 296734 256170 296802 256226
rect 296858 256170 327398 256226
rect 327454 256170 327522 256226
rect 327578 256170 358118 256226
rect 358174 256170 358242 256226
rect 358298 256170 388838 256226
rect 388894 256170 388962 256226
rect 389018 256170 419558 256226
rect 419614 256170 419682 256226
rect 419738 256170 450278 256226
rect 450334 256170 450402 256226
rect 450458 256170 480998 256226
rect 481054 256170 481122 256226
rect 481178 256170 507250 256226
rect 507306 256170 507374 256226
rect 507430 256170 507498 256226
rect 507554 256170 507622 256226
rect 507678 256170 525250 256226
rect 525306 256170 525374 256226
rect 525430 256170 525498 256226
rect 525554 256170 525622 256226
rect 525678 256170 543250 256226
rect 543306 256170 543374 256226
rect 543430 256170 543498 256226
rect 543554 256170 543622 256226
rect 543678 256170 561250 256226
rect 561306 256170 561374 256226
rect 561430 256170 561498 256226
rect 561554 256170 561622 256226
rect 561678 256170 579250 256226
rect 579306 256170 579374 256226
rect 579430 256170 579498 256226
rect 579554 256170 579622 256226
rect 579678 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 3250 256102
rect 3306 256046 3374 256102
rect 3430 256046 3498 256102
rect 3554 256046 3622 256102
rect 3678 256046 21250 256102
rect 21306 256046 21374 256102
rect 21430 256046 21498 256102
rect 21554 256046 21622 256102
rect 21678 256046 39250 256102
rect 39306 256046 39374 256102
rect 39430 256046 39498 256102
rect 39554 256046 39622 256102
rect 39678 256046 57250 256102
rect 57306 256046 57374 256102
rect 57430 256046 57498 256102
rect 57554 256046 57622 256102
rect 57678 256046 75250 256102
rect 75306 256046 75374 256102
rect 75430 256046 75498 256102
rect 75554 256046 75622 256102
rect 75678 256046 93250 256102
rect 93306 256046 93374 256102
rect 93430 256046 93498 256102
rect 93554 256046 93622 256102
rect 93678 256046 111250 256102
rect 111306 256046 111374 256102
rect 111430 256046 111498 256102
rect 111554 256046 111622 256102
rect 111678 256046 129250 256102
rect 129306 256046 129374 256102
rect 129430 256046 129498 256102
rect 129554 256046 129622 256102
rect 129678 256046 147250 256102
rect 147306 256046 147374 256102
rect 147430 256046 147498 256102
rect 147554 256046 147622 256102
rect 147678 256046 165250 256102
rect 165306 256046 165374 256102
rect 165430 256046 165498 256102
rect 165554 256046 165622 256102
rect 165678 256046 183250 256102
rect 183306 256046 183374 256102
rect 183430 256046 183498 256102
rect 183554 256046 183622 256102
rect 183678 256046 201250 256102
rect 201306 256046 201374 256102
rect 201430 256046 201498 256102
rect 201554 256046 201622 256102
rect 201678 256046 204518 256102
rect 204574 256046 204642 256102
rect 204698 256046 235238 256102
rect 235294 256046 235362 256102
rect 235418 256046 265958 256102
rect 266014 256046 266082 256102
rect 266138 256046 296678 256102
rect 296734 256046 296802 256102
rect 296858 256046 327398 256102
rect 327454 256046 327522 256102
rect 327578 256046 358118 256102
rect 358174 256046 358242 256102
rect 358298 256046 388838 256102
rect 388894 256046 388962 256102
rect 389018 256046 419558 256102
rect 419614 256046 419682 256102
rect 419738 256046 450278 256102
rect 450334 256046 450402 256102
rect 450458 256046 480998 256102
rect 481054 256046 481122 256102
rect 481178 256046 507250 256102
rect 507306 256046 507374 256102
rect 507430 256046 507498 256102
rect 507554 256046 507622 256102
rect 507678 256046 525250 256102
rect 525306 256046 525374 256102
rect 525430 256046 525498 256102
rect 525554 256046 525622 256102
rect 525678 256046 543250 256102
rect 543306 256046 543374 256102
rect 543430 256046 543498 256102
rect 543554 256046 543622 256102
rect 543678 256046 561250 256102
rect 561306 256046 561374 256102
rect 561430 256046 561498 256102
rect 561554 256046 561622 256102
rect 561678 256046 579250 256102
rect 579306 256046 579374 256102
rect 579430 256046 579498 256102
rect 579554 256046 579622 256102
rect 579678 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 3250 255978
rect 3306 255922 3374 255978
rect 3430 255922 3498 255978
rect 3554 255922 3622 255978
rect 3678 255922 21250 255978
rect 21306 255922 21374 255978
rect 21430 255922 21498 255978
rect 21554 255922 21622 255978
rect 21678 255922 39250 255978
rect 39306 255922 39374 255978
rect 39430 255922 39498 255978
rect 39554 255922 39622 255978
rect 39678 255922 57250 255978
rect 57306 255922 57374 255978
rect 57430 255922 57498 255978
rect 57554 255922 57622 255978
rect 57678 255922 75250 255978
rect 75306 255922 75374 255978
rect 75430 255922 75498 255978
rect 75554 255922 75622 255978
rect 75678 255922 93250 255978
rect 93306 255922 93374 255978
rect 93430 255922 93498 255978
rect 93554 255922 93622 255978
rect 93678 255922 111250 255978
rect 111306 255922 111374 255978
rect 111430 255922 111498 255978
rect 111554 255922 111622 255978
rect 111678 255922 129250 255978
rect 129306 255922 129374 255978
rect 129430 255922 129498 255978
rect 129554 255922 129622 255978
rect 129678 255922 147250 255978
rect 147306 255922 147374 255978
rect 147430 255922 147498 255978
rect 147554 255922 147622 255978
rect 147678 255922 165250 255978
rect 165306 255922 165374 255978
rect 165430 255922 165498 255978
rect 165554 255922 165622 255978
rect 165678 255922 183250 255978
rect 183306 255922 183374 255978
rect 183430 255922 183498 255978
rect 183554 255922 183622 255978
rect 183678 255922 201250 255978
rect 201306 255922 201374 255978
rect 201430 255922 201498 255978
rect 201554 255922 201622 255978
rect 201678 255922 204518 255978
rect 204574 255922 204642 255978
rect 204698 255922 235238 255978
rect 235294 255922 235362 255978
rect 235418 255922 265958 255978
rect 266014 255922 266082 255978
rect 266138 255922 296678 255978
rect 296734 255922 296802 255978
rect 296858 255922 327398 255978
rect 327454 255922 327522 255978
rect 327578 255922 358118 255978
rect 358174 255922 358242 255978
rect 358298 255922 388838 255978
rect 388894 255922 388962 255978
rect 389018 255922 419558 255978
rect 419614 255922 419682 255978
rect 419738 255922 450278 255978
rect 450334 255922 450402 255978
rect 450458 255922 480998 255978
rect 481054 255922 481122 255978
rect 481178 255922 507250 255978
rect 507306 255922 507374 255978
rect 507430 255922 507498 255978
rect 507554 255922 507622 255978
rect 507678 255922 525250 255978
rect 525306 255922 525374 255978
rect 525430 255922 525498 255978
rect 525554 255922 525622 255978
rect 525678 255922 543250 255978
rect 543306 255922 543374 255978
rect 543430 255922 543498 255978
rect 543554 255922 543622 255978
rect 543678 255922 561250 255978
rect 561306 255922 561374 255978
rect 561430 255922 561498 255978
rect 561554 255922 561622 255978
rect 561678 255922 579250 255978
rect 579306 255922 579374 255978
rect 579430 255922 579498 255978
rect 579554 255922 579622 255978
rect 579678 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 6970 244350
rect 7026 244294 7094 244350
rect 7150 244294 7218 244350
rect 7274 244294 7342 244350
rect 7398 244294 24970 244350
rect 25026 244294 25094 244350
rect 25150 244294 25218 244350
rect 25274 244294 25342 244350
rect 25398 244294 42970 244350
rect 43026 244294 43094 244350
rect 43150 244294 43218 244350
rect 43274 244294 43342 244350
rect 43398 244294 60970 244350
rect 61026 244294 61094 244350
rect 61150 244294 61218 244350
rect 61274 244294 61342 244350
rect 61398 244294 78970 244350
rect 79026 244294 79094 244350
rect 79150 244294 79218 244350
rect 79274 244294 79342 244350
rect 79398 244294 96970 244350
rect 97026 244294 97094 244350
rect 97150 244294 97218 244350
rect 97274 244294 97342 244350
rect 97398 244294 114970 244350
rect 115026 244294 115094 244350
rect 115150 244294 115218 244350
rect 115274 244294 115342 244350
rect 115398 244294 132970 244350
rect 133026 244294 133094 244350
rect 133150 244294 133218 244350
rect 133274 244294 133342 244350
rect 133398 244294 150970 244350
rect 151026 244294 151094 244350
rect 151150 244294 151218 244350
rect 151274 244294 151342 244350
rect 151398 244294 168970 244350
rect 169026 244294 169094 244350
rect 169150 244294 169218 244350
rect 169274 244294 169342 244350
rect 169398 244294 186970 244350
rect 187026 244294 187094 244350
rect 187150 244294 187218 244350
rect 187274 244294 187342 244350
rect 187398 244294 219878 244350
rect 219934 244294 220002 244350
rect 220058 244294 250598 244350
rect 250654 244294 250722 244350
rect 250778 244294 281318 244350
rect 281374 244294 281442 244350
rect 281498 244294 312038 244350
rect 312094 244294 312162 244350
rect 312218 244294 342758 244350
rect 342814 244294 342882 244350
rect 342938 244294 373478 244350
rect 373534 244294 373602 244350
rect 373658 244294 404198 244350
rect 404254 244294 404322 244350
rect 404378 244294 434918 244350
rect 434974 244294 435042 244350
rect 435098 244294 465638 244350
rect 465694 244294 465762 244350
rect 465818 244294 496358 244350
rect 496414 244294 496482 244350
rect 496538 244294 510970 244350
rect 511026 244294 511094 244350
rect 511150 244294 511218 244350
rect 511274 244294 511342 244350
rect 511398 244294 528970 244350
rect 529026 244294 529094 244350
rect 529150 244294 529218 244350
rect 529274 244294 529342 244350
rect 529398 244294 546970 244350
rect 547026 244294 547094 244350
rect 547150 244294 547218 244350
rect 547274 244294 547342 244350
rect 547398 244294 564970 244350
rect 565026 244294 565094 244350
rect 565150 244294 565218 244350
rect 565274 244294 565342 244350
rect 565398 244294 582970 244350
rect 583026 244294 583094 244350
rect 583150 244294 583218 244350
rect 583274 244294 583342 244350
rect 583398 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 6970 244226
rect 7026 244170 7094 244226
rect 7150 244170 7218 244226
rect 7274 244170 7342 244226
rect 7398 244170 24970 244226
rect 25026 244170 25094 244226
rect 25150 244170 25218 244226
rect 25274 244170 25342 244226
rect 25398 244170 42970 244226
rect 43026 244170 43094 244226
rect 43150 244170 43218 244226
rect 43274 244170 43342 244226
rect 43398 244170 60970 244226
rect 61026 244170 61094 244226
rect 61150 244170 61218 244226
rect 61274 244170 61342 244226
rect 61398 244170 78970 244226
rect 79026 244170 79094 244226
rect 79150 244170 79218 244226
rect 79274 244170 79342 244226
rect 79398 244170 96970 244226
rect 97026 244170 97094 244226
rect 97150 244170 97218 244226
rect 97274 244170 97342 244226
rect 97398 244170 114970 244226
rect 115026 244170 115094 244226
rect 115150 244170 115218 244226
rect 115274 244170 115342 244226
rect 115398 244170 132970 244226
rect 133026 244170 133094 244226
rect 133150 244170 133218 244226
rect 133274 244170 133342 244226
rect 133398 244170 150970 244226
rect 151026 244170 151094 244226
rect 151150 244170 151218 244226
rect 151274 244170 151342 244226
rect 151398 244170 168970 244226
rect 169026 244170 169094 244226
rect 169150 244170 169218 244226
rect 169274 244170 169342 244226
rect 169398 244170 186970 244226
rect 187026 244170 187094 244226
rect 187150 244170 187218 244226
rect 187274 244170 187342 244226
rect 187398 244170 219878 244226
rect 219934 244170 220002 244226
rect 220058 244170 250598 244226
rect 250654 244170 250722 244226
rect 250778 244170 281318 244226
rect 281374 244170 281442 244226
rect 281498 244170 312038 244226
rect 312094 244170 312162 244226
rect 312218 244170 342758 244226
rect 342814 244170 342882 244226
rect 342938 244170 373478 244226
rect 373534 244170 373602 244226
rect 373658 244170 404198 244226
rect 404254 244170 404322 244226
rect 404378 244170 434918 244226
rect 434974 244170 435042 244226
rect 435098 244170 465638 244226
rect 465694 244170 465762 244226
rect 465818 244170 496358 244226
rect 496414 244170 496482 244226
rect 496538 244170 510970 244226
rect 511026 244170 511094 244226
rect 511150 244170 511218 244226
rect 511274 244170 511342 244226
rect 511398 244170 528970 244226
rect 529026 244170 529094 244226
rect 529150 244170 529218 244226
rect 529274 244170 529342 244226
rect 529398 244170 546970 244226
rect 547026 244170 547094 244226
rect 547150 244170 547218 244226
rect 547274 244170 547342 244226
rect 547398 244170 564970 244226
rect 565026 244170 565094 244226
rect 565150 244170 565218 244226
rect 565274 244170 565342 244226
rect 565398 244170 582970 244226
rect 583026 244170 583094 244226
rect 583150 244170 583218 244226
rect 583274 244170 583342 244226
rect 583398 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 6970 244102
rect 7026 244046 7094 244102
rect 7150 244046 7218 244102
rect 7274 244046 7342 244102
rect 7398 244046 24970 244102
rect 25026 244046 25094 244102
rect 25150 244046 25218 244102
rect 25274 244046 25342 244102
rect 25398 244046 42970 244102
rect 43026 244046 43094 244102
rect 43150 244046 43218 244102
rect 43274 244046 43342 244102
rect 43398 244046 60970 244102
rect 61026 244046 61094 244102
rect 61150 244046 61218 244102
rect 61274 244046 61342 244102
rect 61398 244046 78970 244102
rect 79026 244046 79094 244102
rect 79150 244046 79218 244102
rect 79274 244046 79342 244102
rect 79398 244046 96970 244102
rect 97026 244046 97094 244102
rect 97150 244046 97218 244102
rect 97274 244046 97342 244102
rect 97398 244046 114970 244102
rect 115026 244046 115094 244102
rect 115150 244046 115218 244102
rect 115274 244046 115342 244102
rect 115398 244046 132970 244102
rect 133026 244046 133094 244102
rect 133150 244046 133218 244102
rect 133274 244046 133342 244102
rect 133398 244046 150970 244102
rect 151026 244046 151094 244102
rect 151150 244046 151218 244102
rect 151274 244046 151342 244102
rect 151398 244046 168970 244102
rect 169026 244046 169094 244102
rect 169150 244046 169218 244102
rect 169274 244046 169342 244102
rect 169398 244046 186970 244102
rect 187026 244046 187094 244102
rect 187150 244046 187218 244102
rect 187274 244046 187342 244102
rect 187398 244046 219878 244102
rect 219934 244046 220002 244102
rect 220058 244046 250598 244102
rect 250654 244046 250722 244102
rect 250778 244046 281318 244102
rect 281374 244046 281442 244102
rect 281498 244046 312038 244102
rect 312094 244046 312162 244102
rect 312218 244046 342758 244102
rect 342814 244046 342882 244102
rect 342938 244046 373478 244102
rect 373534 244046 373602 244102
rect 373658 244046 404198 244102
rect 404254 244046 404322 244102
rect 404378 244046 434918 244102
rect 434974 244046 435042 244102
rect 435098 244046 465638 244102
rect 465694 244046 465762 244102
rect 465818 244046 496358 244102
rect 496414 244046 496482 244102
rect 496538 244046 510970 244102
rect 511026 244046 511094 244102
rect 511150 244046 511218 244102
rect 511274 244046 511342 244102
rect 511398 244046 528970 244102
rect 529026 244046 529094 244102
rect 529150 244046 529218 244102
rect 529274 244046 529342 244102
rect 529398 244046 546970 244102
rect 547026 244046 547094 244102
rect 547150 244046 547218 244102
rect 547274 244046 547342 244102
rect 547398 244046 564970 244102
rect 565026 244046 565094 244102
rect 565150 244046 565218 244102
rect 565274 244046 565342 244102
rect 565398 244046 582970 244102
rect 583026 244046 583094 244102
rect 583150 244046 583218 244102
rect 583274 244046 583342 244102
rect 583398 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 6970 243978
rect 7026 243922 7094 243978
rect 7150 243922 7218 243978
rect 7274 243922 7342 243978
rect 7398 243922 24970 243978
rect 25026 243922 25094 243978
rect 25150 243922 25218 243978
rect 25274 243922 25342 243978
rect 25398 243922 42970 243978
rect 43026 243922 43094 243978
rect 43150 243922 43218 243978
rect 43274 243922 43342 243978
rect 43398 243922 60970 243978
rect 61026 243922 61094 243978
rect 61150 243922 61218 243978
rect 61274 243922 61342 243978
rect 61398 243922 78970 243978
rect 79026 243922 79094 243978
rect 79150 243922 79218 243978
rect 79274 243922 79342 243978
rect 79398 243922 96970 243978
rect 97026 243922 97094 243978
rect 97150 243922 97218 243978
rect 97274 243922 97342 243978
rect 97398 243922 114970 243978
rect 115026 243922 115094 243978
rect 115150 243922 115218 243978
rect 115274 243922 115342 243978
rect 115398 243922 132970 243978
rect 133026 243922 133094 243978
rect 133150 243922 133218 243978
rect 133274 243922 133342 243978
rect 133398 243922 150970 243978
rect 151026 243922 151094 243978
rect 151150 243922 151218 243978
rect 151274 243922 151342 243978
rect 151398 243922 168970 243978
rect 169026 243922 169094 243978
rect 169150 243922 169218 243978
rect 169274 243922 169342 243978
rect 169398 243922 186970 243978
rect 187026 243922 187094 243978
rect 187150 243922 187218 243978
rect 187274 243922 187342 243978
rect 187398 243922 219878 243978
rect 219934 243922 220002 243978
rect 220058 243922 250598 243978
rect 250654 243922 250722 243978
rect 250778 243922 281318 243978
rect 281374 243922 281442 243978
rect 281498 243922 312038 243978
rect 312094 243922 312162 243978
rect 312218 243922 342758 243978
rect 342814 243922 342882 243978
rect 342938 243922 373478 243978
rect 373534 243922 373602 243978
rect 373658 243922 404198 243978
rect 404254 243922 404322 243978
rect 404378 243922 434918 243978
rect 434974 243922 435042 243978
rect 435098 243922 465638 243978
rect 465694 243922 465762 243978
rect 465818 243922 496358 243978
rect 496414 243922 496482 243978
rect 496538 243922 510970 243978
rect 511026 243922 511094 243978
rect 511150 243922 511218 243978
rect 511274 243922 511342 243978
rect 511398 243922 528970 243978
rect 529026 243922 529094 243978
rect 529150 243922 529218 243978
rect 529274 243922 529342 243978
rect 529398 243922 546970 243978
rect 547026 243922 547094 243978
rect 547150 243922 547218 243978
rect 547274 243922 547342 243978
rect 547398 243922 564970 243978
rect 565026 243922 565094 243978
rect 565150 243922 565218 243978
rect 565274 243922 565342 243978
rect 565398 243922 582970 243978
rect 583026 243922 583094 243978
rect 583150 243922 583218 243978
rect 583274 243922 583342 243978
rect 583398 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 3250 238350
rect 3306 238294 3374 238350
rect 3430 238294 3498 238350
rect 3554 238294 3622 238350
rect 3678 238294 21250 238350
rect 21306 238294 21374 238350
rect 21430 238294 21498 238350
rect 21554 238294 21622 238350
rect 21678 238294 39250 238350
rect 39306 238294 39374 238350
rect 39430 238294 39498 238350
rect 39554 238294 39622 238350
rect 39678 238294 57250 238350
rect 57306 238294 57374 238350
rect 57430 238294 57498 238350
rect 57554 238294 57622 238350
rect 57678 238294 75250 238350
rect 75306 238294 75374 238350
rect 75430 238294 75498 238350
rect 75554 238294 75622 238350
rect 75678 238294 93250 238350
rect 93306 238294 93374 238350
rect 93430 238294 93498 238350
rect 93554 238294 93622 238350
rect 93678 238294 111250 238350
rect 111306 238294 111374 238350
rect 111430 238294 111498 238350
rect 111554 238294 111622 238350
rect 111678 238294 129250 238350
rect 129306 238294 129374 238350
rect 129430 238294 129498 238350
rect 129554 238294 129622 238350
rect 129678 238294 147250 238350
rect 147306 238294 147374 238350
rect 147430 238294 147498 238350
rect 147554 238294 147622 238350
rect 147678 238294 165250 238350
rect 165306 238294 165374 238350
rect 165430 238294 165498 238350
rect 165554 238294 165622 238350
rect 165678 238294 183250 238350
rect 183306 238294 183374 238350
rect 183430 238294 183498 238350
rect 183554 238294 183622 238350
rect 183678 238294 201250 238350
rect 201306 238294 201374 238350
rect 201430 238294 201498 238350
rect 201554 238294 201622 238350
rect 201678 238294 204518 238350
rect 204574 238294 204642 238350
rect 204698 238294 235238 238350
rect 235294 238294 235362 238350
rect 235418 238294 265958 238350
rect 266014 238294 266082 238350
rect 266138 238294 296678 238350
rect 296734 238294 296802 238350
rect 296858 238294 327398 238350
rect 327454 238294 327522 238350
rect 327578 238294 358118 238350
rect 358174 238294 358242 238350
rect 358298 238294 388838 238350
rect 388894 238294 388962 238350
rect 389018 238294 419558 238350
rect 419614 238294 419682 238350
rect 419738 238294 450278 238350
rect 450334 238294 450402 238350
rect 450458 238294 480998 238350
rect 481054 238294 481122 238350
rect 481178 238294 507250 238350
rect 507306 238294 507374 238350
rect 507430 238294 507498 238350
rect 507554 238294 507622 238350
rect 507678 238294 525250 238350
rect 525306 238294 525374 238350
rect 525430 238294 525498 238350
rect 525554 238294 525622 238350
rect 525678 238294 543250 238350
rect 543306 238294 543374 238350
rect 543430 238294 543498 238350
rect 543554 238294 543622 238350
rect 543678 238294 561250 238350
rect 561306 238294 561374 238350
rect 561430 238294 561498 238350
rect 561554 238294 561622 238350
rect 561678 238294 579250 238350
rect 579306 238294 579374 238350
rect 579430 238294 579498 238350
rect 579554 238294 579622 238350
rect 579678 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 3250 238226
rect 3306 238170 3374 238226
rect 3430 238170 3498 238226
rect 3554 238170 3622 238226
rect 3678 238170 21250 238226
rect 21306 238170 21374 238226
rect 21430 238170 21498 238226
rect 21554 238170 21622 238226
rect 21678 238170 39250 238226
rect 39306 238170 39374 238226
rect 39430 238170 39498 238226
rect 39554 238170 39622 238226
rect 39678 238170 57250 238226
rect 57306 238170 57374 238226
rect 57430 238170 57498 238226
rect 57554 238170 57622 238226
rect 57678 238170 75250 238226
rect 75306 238170 75374 238226
rect 75430 238170 75498 238226
rect 75554 238170 75622 238226
rect 75678 238170 93250 238226
rect 93306 238170 93374 238226
rect 93430 238170 93498 238226
rect 93554 238170 93622 238226
rect 93678 238170 111250 238226
rect 111306 238170 111374 238226
rect 111430 238170 111498 238226
rect 111554 238170 111622 238226
rect 111678 238170 129250 238226
rect 129306 238170 129374 238226
rect 129430 238170 129498 238226
rect 129554 238170 129622 238226
rect 129678 238170 147250 238226
rect 147306 238170 147374 238226
rect 147430 238170 147498 238226
rect 147554 238170 147622 238226
rect 147678 238170 165250 238226
rect 165306 238170 165374 238226
rect 165430 238170 165498 238226
rect 165554 238170 165622 238226
rect 165678 238170 183250 238226
rect 183306 238170 183374 238226
rect 183430 238170 183498 238226
rect 183554 238170 183622 238226
rect 183678 238170 201250 238226
rect 201306 238170 201374 238226
rect 201430 238170 201498 238226
rect 201554 238170 201622 238226
rect 201678 238170 204518 238226
rect 204574 238170 204642 238226
rect 204698 238170 235238 238226
rect 235294 238170 235362 238226
rect 235418 238170 265958 238226
rect 266014 238170 266082 238226
rect 266138 238170 296678 238226
rect 296734 238170 296802 238226
rect 296858 238170 327398 238226
rect 327454 238170 327522 238226
rect 327578 238170 358118 238226
rect 358174 238170 358242 238226
rect 358298 238170 388838 238226
rect 388894 238170 388962 238226
rect 389018 238170 419558 238226
rect 419614 238170 419682 238226
rect 419738 238170 450278 238226
rect 450334 238170 450402 238226
rect 450458 238170 480998 238226
rect 481054 238170 481122 238226
rect 481178 238170 507250 238226
rect 507306 238170 507374 238226
rect 507430 238170 507498 238226
rect 507554 238170 507622 238226
rect 507678 238170 525250 238226
rect 525306 238170 525374 238226
rect 525430 238170 525498 238226
rect 525554 238170 525622 238226
rect 525678 238170 543250 238226
rect 543306 238170 543374 238226
rect 543430 238170 543498 238226
rect 543554 238170 543622 238226
rect 543678 238170 561250 238226
rect 561306 238170 561374 238226
rect 561430 238170 561498 238226
rect 561554 238170 561622 238226
rect 561678 238170 579250 238226
rect 579306 238170 579374 238226
rect 579430 238170 579498 238226
rect 579554 238170 579622 238226
rect 579678 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 3250 238102
rect 3306 238046 3374 238102
rect 3430 238046 3498 238102
rect 3554 238046 3622 238102
rect 3678 238046 21250 238102
rect 21306 238046 21374 238102
rect 21430 238046 21498 238102
rect 21554 238046 21622 238102
rect 21678 238046 39250 238102
rect 39306 238046 39374 238102
rect 39430 238046 39498 238102
rect 39554 238046 39622 238102
rect 39678 238046 57250 238102
rect 57306 238046 57374 238102
rect 57430 238046 57498 238102
rect 57554 238046 57622 238102
rect 57678 238046 75250 238102
rect 75306 238046 75374 238102
rect 75430 238046 75498 238102
rect 75554 238046 75622 238102
rect 75678 238046 93250 238102
rect 93306 238046 93374 238102
rect 93430 238046 93498 238102
rect 93554 238046 93622 238102
rect 93678 238046 111250 238102
rect 111306 238046 111374 238102
rect 111430 238046 111498 238102
rect 111554 238046 111622 238102
rect 111678 238046 129250 238102
rect 129306 238046 129374 238102
rect 129430 238046 129498 238102
rect 129554 238046 129622 238102
rect 129678 238046 147250 238102
rect 147306 238046 147374 238102
rect 147430 238046 147498 238102
rect 147554 238046 147622 238102
rect 147678 238046 165250 238102
rect 165306 238046 165374 238102
rect 165430 238046 165498 238102
rect 165554 238046 165622 238102
rect 165678 238046 183250 238102
rect 183306 238046 183374 238102
rect 183430 238046 183498 238102
rect 183554 238046 183622 238102
rect 183678 238046 201250 238102
rect 201306 238046 201374 238102
rect 201430 238046 201498 238102
rect 201554 238046 201622 238102
rect 201678 238046 204518 238102
rect 204574 238046 204642 238102
rect 204698 238046 235238 238102
rect 235294 238046 235362 238102
rect 235418 238046 265958 238102
rect 266014 238046 266082 238102
rect 266138 238046 296678 238102
rect 296734 238046 296802 238102
rect 296858 238046 327398 238102
rect 327454 238046 327522 238102
rect 327578 238046 358118 238102
rect 358174 238046 358242 238102
rect 358298 238046 388838 238102
rect 388894 238046 388962 238102
rect 389018 238046 419558 238102
rect 419614 238046 419682 238102
rect 419738 238046 450278 238102
rect 450334 238046 450402 238102
rect 450458 238046 480998 238102
rect 481054 238046 481122 238102
rect 481178 238046 507250 238102
rect 507306 238046 507374 238102
rect 507430 238046 507498 238102
rect 507554 238046 507622 238102
rect 507678 238046 525250 238102
rect 525306 238046 525374 238102
rect 525430 238046 525498 238102
rect 525554 238046 525622 238102
rect 525678 238046 543250 238102
rect 543306 238046 543374 238102
rect 543430 238046 543498 238102
rect 543554 238046 543622 238102
rect 543678 238046 561250 238102
rect 561306 238046 561374 238102
rect 561430 238046 561498 238102
rect 561554 238046 561622 238102
rect 561678 238046 579250 238102
rect 579306 238046 579374 238102
rect 579430 238046 579498 238102
rect 579554 238046 579622 238102
rect 579678 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 3250 237978
rect 3306 237922 3374 237978
rect 3430 237922 3498 237978
rect 3554 237922 3622 237978
rect 3678 237922 21250 237978
rect 21306 237922 21374 237978
rect 21430 237922 21498 237978
rect 21554 237922 21622 237978
rect 21678 237922 39250 237978
rect 39306 237922 39374 237978
rect 39430 237922 39498 237978
rect 39554 237922 39622 237978
rect 39678 237922 57250 237978
rect 57306 237922 57374 237978
rect 57430 237922 57498 237978
rect 57554 237922 57622 237978
rect 57678 237922 75250 237978
rect 75306 237922 75374 237978
rect 75430 237922 75498 237978
rect 75554 237922 75622 237978
rect 75678 237922 93250 237978
rect 93306 237922 93374 237978
rect 93430 237922 93498 237978
rect 93554 237922 93622 237978
rect 93678 237922 111250 237978
rect 111306 237922 111374 237978
rect 111430 237922 111498 237978
rect 111554 237922 111622 237978
rect 111678 237922 129250 237978
rect 129306 237922 129374 237978
rect 129430 237922 129498 237978
rect 129554 237922 129622 237978
rect 129678 237922 147250 237978
rect 147306 237922 147374 237978
rect 147430 237922 147498 237978
rect 147554 237922 147622 237978
rect 147678 237922 165250 237978
rect 165306 237922 165374 237978
rect 165430 237922 165498 237978
rect 165554 237922 165622 237978
rect 165678 237922 183250 237978
rect 183306 237922 183374 237978
rect 183430 237922 183498 237978
rect 183554 237922 183622 237978
rect 183678 237922 201250 237978
rect 201306 237922 201374 237978
rect 201430 237922 201498 237978
rect 201554 237922 201622 237978
rect 201678 237922 204518 237978
rect 204574 237922 204642 237978
rect 204698 237922 235238 237978
rect 235294 237922 235362 237978
rect 235418 237922 265958 237978
rect 266014 237922 266082 237978
rect 266138 237922 296678 237978
rect 296734 237922 296802 237978
rect 296858 237922 327398 237978
rect 327454 237922 327522 237978
rect 327578 237922 358118 237978
rect 358174 237922 358242 237978
rect 358298 237922 388838 237978
rect 388894 237922 388962 237978
rect 389018 237922 419558 237978
rect 419614 237922 419682 237978
rect 419738 237922 450278 237978
rect 450334 237922 450402 237978
rect 450458 237922 480998 237978
rect 481054 237922 481122 237978
rect 481178 237922 507250 237978
rect 507306 237922 507374 237978
rect 507430 237922 507498 237978
rect 507554 237922 507622 237978
rect 507678 237922 525250 237978
rect 525306 237922 525374 237978
rect 525430 237922 525498 237978
rect 525554 237922 525622 237978
rect 525678 237922 543250 237978
rect 543306 237922 543374 237978
rect 543430 237922 543498 237978
rect 543554 237922 543622 237978
rect 543678 237922 561250 237978
rect 561306 237922 561374 237978
rect 561430 237922 561498 237978
rect 561554 237922 561622 237978
rect 561678 237922 579250 237978
rect 579306 237922 579374 237978
rect 579430 237922 579498 237978
rect 579554 237922 579622 237978
rect 579678 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 6970 226350
rect 7026 226294 7094 226350
rect 7150 226294 7218 226350
rect 7274 226294 7342 226350
rect 7398 226294 24970 226350
rect 25026 226294 25094 226350
rect 25150 226294 25218 226350
rect 25274 226294 25342 226350
rect 25398 226294 42970 226350
rect 43026 226294 43094 226350
rect 43150 226294 43218 226350
rect 43274 226294 43342 226350
rect 43398 226294 60970 226350
rect 61026 226294 61094 226350
rect 61150 226294 61218 226350
rect 61274 226294 61342 226350
rect 61398 226294 78970 226350
rect 79026 226294 79094 226350
rect 79150 226294 79218 226350
rect 79274 226294 79342 226350
rect 79398 226294 96970 226350
rect 97026 226294 97094 226350
rect 97150 226294 97218 226350
rect 97274 226294 97342 226350
rect 97398 226294 114970 226350
rect 115026 226294 115094 226350
rect 115150 226294 115218 226350
rect 115274 226294 115342 226350
rect 115398 226294 132970 226350
rect 133026 226294 133094 226350
rect 133150 226294 133218 226350
rect 133274 226294 133342 226350
rect 133398 226294 150970 226350
rect 151026 226294 151094 226350
rect 151150 226294 151218 226350
rect 151274 226294 151342 226350
rect 151398 226294 168970 226350
rect 169026 226294 169094 226350
rect 169150 226294 169218 226350
rect 169274 226294 169342 226350
rect 169398 226294 186970 226350
rect 187026 226294 187094 226350
rect 187150 226294 187218 226350
rect 187274 226294 187342 226350
rect 187398 226294 219878 226350
rect 219934 226294 220002 226350
rect 220058 226294 250598 226350
rect 250654 226294 250722 226350
rect 250778 226294 281318 226350
rect 281374 226294 281442 226350
rect 281498 226294 312038 226350
rect 312094 226294 312162 226350
rect 312218 226294 342758 226350
rect 342814 226294 342882 226350
rect 342938 226294 373478 226350
rect 373534 226294 373602 226350
rect 373658 226294 404198 226350
rect 404254 226294 404322 226350
rect 404378 226294 434918 226350
rect 434974 226294 435042 226350
rect 435098 226294 465638 226350
rect 465694 226294 465762 226350
rect 465818 226294 496358 226350
rect 496414 226294 496482 226350
rect 496538 226294 510970 226350
rect 511026 226294 511094 226350
rect 511150 226294 511218 226350
rect 511274 226294 511342 226350
rect 511398 226294 528970 226350
rect 529026 226294 529094 226350
rect 529150 226294 529218 226350
rect 529274 226294 529342 226350
rect 529398 226294 546970 226350
rect 547026 226294 547094 226350
rect 547150 226294 547218 226350
rect 547274 226294 547342 226350
rect 547398 226294 564970 226350
rect 565026 226294 565094 226350
rect 565150 226294 565218 226350
rect 565274 226294 565342 226350
rect 565398 226294 582970 226350
rect 583026 226294 583094 226350
rect 583150 226294 583218 226350
rect 583274 226294 583342 226350
rect 583398 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 6970 226226
rect 7026 226170 7094 226226
rect 7150 226170 7218 226226
rect 7274 226170 7342 226226
rect 7398 226170 24970 226226
rect 25026 226170 25094 226226
rect 25150 226170 25218 226226
rect 25274 226170 25342 226226
rect 25398 226170 42970 226226
rect 43026 226170 43094 226226
rect 43150 226170 43218 226226
rect 43274 226170 43342 226226
rect 43398 226170 60970 226226
rect 61026 226170 61094 226226
rect 61150 226170 61218 226226
rect 61274 226170 61342 226226
rect 61398 226170 78970 226226
rect 79026 226170 79094 226226
rect 79150 226170 79218 226226
rect 79274 226170 79342 226226
rect 79398 226170 96970 226226
rect 97026 226170 97094 226226
rect 97150 226170 97218 226226
rect 97274 226170 97342 226226
rect 97398 226170 114970 226226
rect 115026 226170 115094 226226
rect 115150 226170 115218 226226
rect 115274 226170 115342 226226
rect 115398 226170 132970 226226
rect 133026 226170 133094 226226
rect 133150 226170 133218 226226
rect 133274 226170 133342 226226
rect 133398 226170 150970 226226
rect 151026 226170 151094 226226
rect 151150 226170 151218 226226
rect 151274 226170 151342 226226
rect 151398 226170 168970 226226
rect 169026 226170 169094 226226
rect 169150 226170 169218 226226
rect 169274 226170 169342 226226
rect 169398 226170 186970 226226
rect 187026 226170 187094 226226
rect 187150 226170 187218 226226
rect 187274 226170 187342 226226
rect 187398 226170 219878 226226
rect 219934 226170 220002 226226
rect 220058 226170 250598 226226
rect 250654 226170 250722 226226
rect 250778 226170 281318 226226
rect 281374 226170 281442 226226
rect 281498 226170 312038 226226
rect 312094 226170 312162 226226
rect 312218 226170 342758 226226
rect 342814 226170 342882 226226
rect 342938 226170 373478 226226
rect 373534 226170 373602 226226
rect 373658 226170 404198 226226
rect 404254 226170 404322 226226
rect 404378 226170 434918 226226
rect 434974 226170 435042 226226
rect 435098 226170 465638 226226
rect 465694 226170 465762 226226
rect 465818 226170 496358 226226
rect 496414 226170 496482 226226
rect 496538 226170 510970 226226
rect 511026 226170 511094 226226
rect 511150 226170 511218 226226
rect 511274 226170 511342 226226
rect 511398 226170 528970 226226
rect 529026 226170 529094 226226
rect 529150 226170 529218 226226
rect 529274 226170 529342 226226
rect 529398 226170 546970 226226
rect 547026 226170 547094 226226
rect 547150 226170 547218 226226
rect 547274 226170 547342 226226
rect 547398 226170 564970 226226
rect 565026 226170 565094 226226
rect 565150 226170 565218 226226
rect 565274 226170 565342 226226
rect 565398 226170 582970 226226
rect 583026 226170 583094 226226
rect 583150 226170 583218 226226
rect 583274 226170 583342 226226
rect 583398 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 6970 226102
rect 7026 226046 7094 226102
rect 7150 226046 7218 226102
rect 7274 226046 7342 226102
rect 7398 226046 24970 226102
rect 25026 226046 25094 226102
rect 25150 226046 25218 226102
rect 25274 226046 25342 226102
rect 25398 226046 42970 226102
rect 43026 226046 43094 226102
rect 43150 226046 43218 226102
rect 43274 226046 43342 226102
rect 43398 226046 60970 226102
rect 61026 226046 61094 226102
rect 61150 226046 61218 226102
rect 61274 226046 61342 226102
rect 61398 226046 78970 226102
rect 79026 226046 79094 226102
rect 79150 226046 79218 226102
rect 79274 226046 79342 226102
rect 79398 226046 96970 226102
rect 97026 226046 97094 226102
rect 97150 226046 97218 226102
rect 97274 226046 97342 226102
rect 97398 226046 114970 226102
rect 115026 226046 115094 226102
rect 115150 226046 115218 226102
rect 115274 226046 115342 226102
rect 115398 226046 132970 226102
rect 133026 226046 133094 226102
rect 133150 226046 133218 226102
rect 133274 226046 133342 226102
rect 133398 226046 150970 226102
rect 151026 226046 151094 226102
rect 151150 226046 151218 226102
rect 151274 226046 151342 226102
rect 151398 226046 168970 226102
rect 169026 226046 169094 226102
rect 169150 226046 169218 226102
rect 169274 226046 169342 226102
rect 169398 226046 186970 226102
rect 187026 226046 187094 226102
rect 187150 226046 187218 226102
rect 187274 226046 187342 226102
rect 187398 226046 219878 226102
rect 219934 226046 220002 226102
rect 220058 226046 250598 226102
rect 250654 226046 250722 226102
rect 250778 226046 281318 226102
rect 281374 226046 281442 226102
rect 281498 226046 312038 226102
rect 312094 226046 312162 226102
rect 312218 226046 342758 226102
rect 342814 226046 342882 226102
rect 342938 226046 373478 226102
rect 373534 226046 373602 226102
rect 373658 226046 404198 226102
rect 404254 226046 404322 226102
rect 404378 226046 434918 226102
rect 434974 226046 435042 226102
rect 435098 226046 465638 226102
rect 465694 226046 465762 226102
rect 465818 226046 496358 226102
rect 496414 226046 496482 226102
rect 496538 226046 510970 226102
rect 511026 226046 511094 226102
rect 511150 226046 511218 226102
rect 511274 226046 511342 226102
rect 511398 226046 528970 226102
rect 529026 226046 529094 226102
rect 529150 226046 529218 226102
rect 529274 226046 529342 226102
rect 529398 226046 546970 226102
rect 547026 226046 547094 226102
rect 547150 226046 547218 226102
rect 547274 226046 547342 226102
rect 547398 226046 564970 226102
rect 565026 226046 565094 226102
rect 565150 226046 565218 226102
rect 565274 226046 565342 226102
rect 565398 226046 582970 226102
rect 583026 226046 583094 226102
rect 583150 226046 583218 226102
rect 583274 226046 583342 226102
rect 583398 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 6970 225978
rect 7026 225922 7094 225978
rect 7150 225922 7218 225978
rect 7274 225922 7342 225978
rect 7398 225922 24970 225978
rect 25026 225922 25094 225978
rect 25150 225922 25218 225978
rect 25274 225922 25342 225978
rect 25398 225922 42970 225978
rect 43026 225922 43094 225978
rect 43150 225922 43218 225978
rect 43274 225922 43342 225978
rect 43398 225922 60970 225978
rect 61026 225922 61094 225978
rect 61150 225922 61218 225978
rect 61274 225922 61342 225978
rect 61398 225922 78970 225978
rect 79026 225922 79094 225978
rect 79150 225922 79218 225978
rect 79274 225922 79342 225978
rect 79398 225922 96970 225978
rect 97026 225922 97094 225978
rect 97150 225922 97218 225978
rect 97274 225922 97342 225978
rect 97398 225922 114970 225978
rect 115026 225922 115094 225978
rect 115150 225922 115218 225978
rect 115274 225922 115342 225978
rect 115398 225922 132970 225978
rect 133026 225922 133094 225978
rect 133150 225922 133218 225978
rect 133274 225922 133342 225978
rect 133398 225922 150970 225978
rect 151026 225922 151094 225978
rect 151150 225922 151218 225978
rect 151274 225922 151342 225978
rect 151398 225922 168970 225978
rect 169026 225922 169094 225978
rect 169150 225922 169218 225978
rect 169274 225922 169342 225978
rect 169398 225922 186970 225978
rect 187026 225922 187094 225978
rect 187150 225922 187218 225978
rect 187274 225922 187342 225978
rect 187398 225922 219878 225978
rect 219934 225922 220002 225978
rect 220058 225922 250598 225978
rect 250654 225922 250722 225978
rect 250778 225922 281318 225978
rect 281374 225922 281442 225978
rect 281498 225922 312038 225978
rect 312094 225922 312162 225978
rect 312218 225922 342758 225978
rect 342814 225922 342882 225978
rect 342938 225922 373478 225978
rect 373534 225922 373602 225978
rect 373658 225922 404198 225978
rect 404254 225922 404322 225978
rect 404378 225922 434918 225978
rect 434974 225922 435042 225978
rect 435098 225922 465638 225978
rect 465694 225922 465762 225978
rect 465818 225922 496358 225978
rect 496414 225922 496482 225978
rect 496538 225922 510970 225978
rect 511026 225922 511094 225978
rect 511150 225922 511218 225978
rect 511274 225922 511342 225978
rect 511398 225922 528970 225978
rect 529026 225922 529094 225978
rect 529150 225922 529218 225978
rect 529274 225922 529342 225978
rect 529398 225922 546970 225978
rect 547026 225922 547094 225978
rect 547150 225922 547218 225978
rect 547274 225922 547342 225978
rect 547398 225922 564970 225978
rect 565026 225922 565094 225978
rect 565150 225922 565218 225978
rect 565274 225922 565342 225978
rect 565398 225922 582970 225978
rect 583026 225922 583094 225978
rect 583150 225922 583218 225978
rect 583274 225922 583342 225978
rect 583398 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 3250 220350
rect 3306 220294 3374 220350
rect 3430 220294 3498 220350
rect 3554 220294 3622 220350
rect 3678 220294 21250 220350
rect 21306 220294 21374 220350
rect 21430 220294 21498 220350
rect 21554 220294 21622 220350
rect 21678 220294 39250 220350
rect 39306 220294 39374 220350
rect 39430 220294 39498 220350
rect 39554 220294 39622 220350
rect 39678 220294 57250 220350
rect 57306 220294 57374 220350
rect 57430 220294 57498 220350
rect 57554 220294 57622 220350
rect 57678 220294 75250 220350
rect 75306 220294 75374 220350
rect 75430 220294 75498 220350
rect 75554 220294 75622 220350
rect 75678 220294 93250 220350
rect 93306 220294 93374 220350
rect 93430 220294 93498 220350
rect 93554 220294 93622 220350
rect 93678 220294 111250 220350
rect 111306 220294 111374 220350
rect 111430 220294 111498 220350
rect 111554 220294 111622 220350
rect 111678 220294 129250 220350
rect 129306 220294 129374 220350
rect 129430 220294 129498 220350
rect 129554 220294 129622 220350
rect 129678 220294 147250 220350
rect 147306 220294 147374 220350
rect 147430 220294 147498 220350
rect 147554 220294 147622 220350
rect 147678 220294 165250 220350
rect 165306 220294 165374 220350
rect 165430 220294 165498 220350
rect 165554 220294 165622 220350
rect 165678 220294 183250 220350
rect 183306 220294 183374 220350
rect 183430 220294 183498 220350
rect 183554 220294 183622 220350
rect 183678 220294 201250 220350
rect 201306 220294 201374 220350
rect 201430 220294 201498 220350
rect 201554 220294 201622 220350
rect 201678 220294 204518 220350
rect 204574 220294 204642 220350
rect 204698 220294 235238 220350
rect 235294 220294 235362 220350
rect 235418 220294 265958 220350
rect 266014 220294 266082 220350
rect 266138 220294 296678 220350
rect 296734 220294 296802 220350
rect 296858 220294 327398 220350
rect 327454 220294 327522 220350
rect 327578 220294 358118 220350
rect 358174 220294 358242 220350
rect 358298 220294 388838 220350
rect 388894 220294 388962 220350
rect 389018 220294 419558 220350
rect 419614 220294 419682 220350
rect 419738 220294 450278 220350
rect 450334 220294 450402 220350
rect 450458 220294 480998 220350
rect 481054 220294 481122 220350
rect 481178 220294 507250 220350
rect 507306 220294 507374 220350
rect 507430 220294 507498 220350
rect 507554 220294 507622 220350
rect 507678 220294 525250 220350
rect 525306 220294 525374 220350
rect 525430 220294 525498 220350
rect 525554 220294 525622 220350
rect 525678 220294 543250 220350
rect 543306 220294 543374 220350
rect 543430 220294 543498 220350
rect 543554 220294 543622 220350
rect 543678 220294 561250 220350
rect 561306 220294 561374 220350
rect 561430 220294 561498 220350
rect 561554 220294 561622 220350
rect 561678 220294 579250 220350
rect 579306 220294 579374 220350
rect 579430 220294 579498 220350
rect 579554 220294 579622 220350
rect 579678 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 3250 220226
rect 3306 220170 3374 220226
rect 3430 220170 3498 220226
rect 3554 220170 3622 220226
rect 3678 220170 21250 220226
rect 21306 220170 21374 220226
rect 21430 220170 21498 220226
rect 21554 220170 21622 220226
rect 21678 220170 39250 220226
rect 39306 220170 39374 220226
rect 39430 220170 39498 220226
rect 39554 220170 39622 220226
rect 39678 220170 57250 220226
rect 57306 220170 57374 220226
rect 57430 220170 57498 220226
rect 57554 220170 57622 220226
rect 57678 220170 75250 220226
rect 75306 220170 75374 220226
rect 75430 220170 75498 220226
rect 75554 220170 75622 220226
rect 75678 220170 93250 220226
rect 93306 220170 93374 220226
rect 93430 220170 93498 220226
rect 93554 220170 93622 220226
rect 93678 220170 111250 220226
rect 111306 220170 111374 220226
rect 111430 220170 111498 220226
rect 111554 220170 111622 220226
rect 111678 220170 129250 220226
rect 129306 220170 129374 220226
rect 129430 220170 129498 220226
rect 129554 220170 129622 220226
rect 129678 220170 147250 220226
rect 147306 220170 147374 220226
rect 147430 220170 147498 220226
rect 147554 220170 147622 220226
rect 147678 220170 165250 220226
rect 165306 220170 165374 220226
rect 165430 220170 165498 220226
rect 165554 220170 165622 220226
rect 165678 220170 183250 220226
rect 183306 220170 183374 220226
rect 183430 220170 183498 220226
rect 183554 220170 183622 220226
rect 183678 220170 201250 220226
rect 201306 220170 201374 220226
rect 201430 220170 201498 220226
rect 201554 220170 201622 220226
rect 201678 220170 204518 220226
rect 204574 220170 204642 220226
rect 204698 220170 235238 220226
rect 235294 220170 235362 220226
rect 235418 220170 265958 220226
rect 266014 220170 266082 220226
rect 266138 220170 296678 220226
rect 296734 220170 296802 220226
rect 296858 220170 327398 220226
rect 327454 220170 327522 220226
rect 327578 220170 358118 220226
rect 358174 220170 358242 220226
rect 358298 220170 388838 220226
rect 388894 220170 388962 220226
rect 389018 220170 419558 220226
rect 419614 220170 419682 220226
rect 419738 220170 450278 220226
rect 450334 220170 450402 220226
rect 450458 220170 480998 220226
rect 481054 220170 481122 220226
rect 481178 220170 507250 220226
rect 507306 220170 507374 220226
rect 507430 220170 507498 220226
rect 507554 220170 507622 220226
rect 507678 220170 525250 220226
rect 525306 220170 525374 220226
rect 525430 220170 525498 220226
rect 525554 220170 525622 220226
rect 525678 220170 543250 220226
rect 543306 220170 543374 220226
rect 543430 220170 543498 220226
rect 543554 220170 543622 220226
rect 543678 220170 561250 220226
rect 561306 220170 561374 220226
rect 561430 220170 561498 220226
rect 561554 220170 561622 220226
rect 561678 220170 579250 220226
rect 579306 220170 579374 220226
rect 579430 220170 579498 220226
rect 579554 220170 579622 220226
rect 579678 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 3250 220102
rect 3306 220046 3374 220102
rect 3430 220046 3498 220102
rect 3554 220046 3622 220102
rect 3678 220046 21250 220102
rect 21306 220046 21374 220102
rect 21430 220046 21498 220102
rect 21554 220046 21622 220102
rect 21678 220046 39250 220102
rect 39306 220046 39374 220102
rect 39430 220046 39498 220102
rect 39554 220046 39622 220102
rect 39678 220046 57250 220102
rect 57306 220046 57374 220102
rect 57430 220046 57498 220102
rect 57554 220046 57622 220102
rect 57678 220046 75250 220102
rect 75306 220046 75374 220102
rect 75430 220046 75498 220102
rect 75554 220046 75622 220102
rect 75678 220046 93250 220102
rect 93306 220046 93374 220102
rect 93430 220046 93498 220102
rect 93554 220046 93622 220102
rect 93678 220046 111250 220102
rect 111306 220046 111374 220102
rect 111430 220046 111498 220102
rect 111554 220046 111622 220102
rect 111678 220046 129250 220102
rect 129306 220046 129374 220102
rect 129430 220046 129498 220102
rect 129554 220046 129622 220102
rect 129678 220046 147250 220102
rect 147306 220046 147374 220102
rect 147430 220046 147498 220102
rect 147554 220046 147622 220102
rect 147678 220046 165250 220102
rect 165306 220046 165374 220102
rect 165430 220046 165498 220102
rect 165554 220046 165622 220102
rect 165678 220046 183250 220102
rect 183306 220046 183374 220102
rect 183430 220046 183498 220102
rect 183554 220046 183622 220102
rect 183678 220046 201250 220102
rect 201306 220046 201374 220102
rect 201430 220046 201498 220102
rect 201554 220046 201622 220102
rect 201678 220046 204518 220102
rect 204574 220046 204642 220102
rect 204698 220046 235238 220102
rect 235294 220046 235362 220102
rect 235418 220046 265958 220102
rect 266014 220046 266082 220102
rect 266138 220046 296678 220102
rect 296734 220046 296802 220102
rect 296858 220046 327398 220102
rect 327454 220046 327522 220102
rect 327578 220046 358118 220102
rect 358174 220046 358242 220102
rect 358298 220046 388838 220102
rect 388894 220046 388962 220102
rect 389018 220046 419558 220102
rect 419614 220046 419682 220102
rect 419738 220046 450278 220102
rect 450334 220046 450402 220102
rect 450458 220046 480998 220102
rect 481054 220046 481122 220102
rect 481178 220046 507250 220102
rect 507306 220046 507374 220102
rect 507430 220046 507498 220102
rect 507554 220046 507622 220102
rect 507678 220046 525250 220102
rect 525306 220046 525374 220102
rect 525430 220046 525498 220102
rect 525554 220046 525622 220102
rect 525678 220046 543250 220102
rect 543306 220046 543374 220102
rect 543430 220046 543498 220102
rect 543554 220046 543622 220102
rect 543678 220046 561250 220102
rect 561306 220046 561374 220102
rect 561430 220046 561498 220102
rect 561554 220046 561622 220102
rect 561678 220046 579250 220102
rect 579306 220046 579374 220102
rect 579430 220046 579498 220102
rect 579554 220046 579622 220102
rect 579678 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 3250 219978
rect 3306 219922 3374 219978
rect 3430 219922 3498 219978
rect 3554 219922 3622 219978
rect 3678 219922 21250 219978
rect 21306 219922 21374 219978
rect 21430 219922 21498 219978
rect 21554 219922 21622 219978
rect 21678 219922 39250 219978
rect 39306 219922 39374 219978
rect 39430 219922 39498 219978
rect 39554 219922 39622 219978
rect 39678 219922 57250 219978
rect 57306 219922 57374 219978
rect 57430 219922 57498 219978
rect 57554 219922 57622 219978
rect 57678 219922 75250 219978
rect 75306 219922 75374 219978
rect 75430 219922 75498 219978
rect 75554 219922 75622 219978
rect 75678 219922 93250 219978
rect 93306 219922 93374 219978
rect 93430 219922 93498 219978
rect 93554 219922 93622 219978
rect 93678 219922 111250 219978
rect 111306 219922 111374 219978
rect 111430 219922 111498 219978
rect 111554 219922 111622 219978
rect 111678 219922 129250 219978
rect 129306 219922 129374 219978
rect 129430 219922 129498 219978
rect 129554 219922 129622 219978
rect 129678 219922 147250 219978
rect 147306 219922 147374 219978
rect 147430 219922 147498 219978
rect 147554 219922 147622 219978
rect 147678 219922 165250 219978
rect 165306 219922 165374 219978
rect 165430 219922 165498 219978
rect 165554 219922 165622 219978
rect 165678 219922 183250 219978
rect 183306 219922 183374 219978
rect 183430 219922 183498 219978
rect 183554 219922 183622 219978
rect 183678 219922 201250 219978
rect 201306 219922 201374 219978
rect 201430 219922 201498 219978
rect 201554 219922 201622 219978
rect 201678 219922 204518 219978
rect 204574 219922 204642 219978
rect 204698 219922 235238 219978
rect 235294 219922 235362 219978
rect 235418 219922 265958 219978
rect 266014 219922 266082 219978
rect 266138 219922 296678 219978
rect 296734 219922 296802 219978
rect 296858 219922 327398 219978
rect 327454 219922 327522 219978
rect 327578 219922 358118 219978
rect 358174 219922 358242 219978
rect 358298 219922 388838 219978
rect 388894 219922 388962 219978
rect 389018 219922 419558 219978
rect 419614 219922 419682 219978
rect 419738 219922 450278 219978
rect 450334 219922 450402 219978
rect 450458 219922 480998 219978
rect 481054 219922 481122 219978
rect 481178 219922 507250 219978
rect 507306 219922 507374 219978
rect 507430 219922 507498 219978
rect 507554 219922 507622 219978
rect 507678 219922 525250 219978
rect 525306 219922 525374 219978
rect 525430 219922 525498 219978
rect 525554 219922 525622 219978
rect 525678 219922 543250 219978
rect 543306 219922 543374 219978
rect 543430 219922 543498 219978
rect 543554 219922 543622 219978
rect 543678 219922 561250 219978
rect 561306 219922 561374 219978
rect 561430 219922 561498 219978
rect 561554 219922 561622 219978
rect 561678 219922 579250 219978
rect 579306 219922 579374 219978
rect 579430 219922 579498 219978
rect 579554 219922 579622 219978
rect 579678 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 6970 208350
rect 7026 208294 7094 208350
rect 7150 208294 7218 208350
rect 7274 208294 7342 208350
rect 7398 208294 24970 208350
rect 25026 208294 25094 208350
rect 25150 208294 25218 208350
rect 25274 208294 25342 208350
rect 25398 208294 42970 208350
rect 43026 208294 43094 208350
rect 43150 208294 43218 208350
rect 43274 208294 43342 208350
rect 43398 208294 60970 208350
rect 61026 208294 61094 208350
rect 61150 208294 61218 208350
rect 61274 208294 61342 208350
rect 61398 208294 78970 208350
rect 79026 208294 79094 208350
rect 79150 208294 79218 208350
rect 79274 208294 79342 208350
rect 79398 208294 96970 208350
rect 97026 208294 97094 208350
rect 97150 208294 97218 208350
rect 97274 208294 97342 208350
rect 97398 208294 114970 208350
rect 115026 208294 115094 208350
rect 115150 208294 115218 208350
rect 115274 208294 115342 208350
rect 115398 208294 132970 208350
rect 133026 208294 133094 208350
rect 133150 208294 133218 208350
rect 133274 208294 133342 208350
rect 133398 208294 150970 208350
rect 151026 208294 151094 208350
rect 151150 208294 151218 208350
rect 151274 208294 151342 208350
rect 151398 208294 168970 208350
rect 169026 208294 169094 208350
rect 169150 208294 169218 208350
rect 169274 208294 169342 208350
rect 169398 208294 186970 208350
rect 187026 208294 187094 208350
rect 187150 208294 187218 208350
rect 187274 208294 187342 208350
rect 187398 208294 204970 208350
rect 205026 208294 205094 208350
rect 205150 208294 205218 208350
rect 205274 208294 205342 208350
rect 205398 208294 219878 208350
rect 219934 208294 220002 208350
rect 220058 208294 222970 208350
rect 223026 208294 223094 208350
rect 223150 208294 223218 208350
rect 223274 208294 223342 208350
rect 223398 208294 240970 208350
rect 241026 208294 241094 208350
rect 241150 208294 241218 208350
rect 241274 208294 241342 208350
rect 241398 208294 250598 208350
rect 250654 208294 250722 208350
rect 250778 208294 258970 208350
rect 259026 208294 259094 208350
rect 259150 208294 259218 208350
rect 259274 208294 259342 208350
rect 259398 208294 276970 208350
rect 277026 208294 277094 208350
rect 277150 208294 277218 208350
rect 277274 208294 277342 208350
rect 277398 208294 281318 208350
rect 281374 208294 281442 208350
rect 281498 208294 294970 208350
rect 295026 208294 295094 208350
rect 295150 208294 295218 208350
rect 295274 208294 295342 208350
rect 295398 208294 312038 208350
rect 312094 208294 312162 208350
rect 312218 208294 312970 208350
rect 313026 208294 313094 208350
rect 313150 208294 313218 208350
rect 313274 208294 313342 208350
rect 313398 208294 330970 208350
rect 331026 208294 331094 208350
rect 331150 208294 331218 208350
rect 331274 208294 331342 208350
rect 331398 208294 342758 208350
rect 342814 208294 342882 208350
rect 342938 208294 348970 208350
rect 349026 208294 349094 208350
rect 349150 208294 349218 208350
rect 349274 208294 349342 208350
rect 349398 208294 366970 208350
rect 367026 208294 367094 208350
rect 367150 208294 367218 208350
rect 367274 208294 367342 208350
rect 367398 208294 373478 208350
rect 373534 208294 373602 208350
rect 373658 208294 384970 208350
rect 385026 208294 385094 208350
rect 385150 208294 385218 208350
rect 385274 208294 385342 208350
rect 385398 208294 402970 208350
rect 403026 208294 403094 208350
rect 403150 208294 403218 208350
rect 403274 208294 403342 208350
rect 403398 208294 404198 208350
rect 404254 208294 404322 208350
rect 404378 208294 420970 208350
rect 421026 208294 421094 208350
rect 421150 208294 421218 208350
rect 421274 208294 421342 208350
rect 421398 208294 434918 208350
rect 434974 208294 435042 208350
rect 435098 208294 438970 208350
rect 439026 208294 439094 208350
rect 439150 208294 439218 208350
rect 439274 208294 439342 208350
rect 439398 208294 456970 208350
rect 457026 208294 457094 208350
rect 457150 208294 457218 208350
rect 457274 208294 457342 208350
rect 457398 208294 465638 208350
rect 465694 208294 465762 208350
rect 465818 208294 474970 208350
rect 475026 208294 475094 208350
rect 475150 208294 475218 208350
rect 475274 208294 475342 208350
rect 475398 208294 492970 208350
rect 493026 208294 493094 208350
rect 493150 208294 493218 208350
rect 493274 208294 493342 208350
rect 493398 208294 496358 208350
rect 496414 208294 496482 208350
rect 496538 208294 510970 208350
rect 511026 208294 511094 208350
rect 511150 208294 511218 208350
rect 511274 208294 511342 208350
rect 511398 208294 528970 208350
rect 529026 208294 529094 208350
rect 529150 208294 529218 208350
rect 529274 208294 529342 208350
rect 529398 208294 546970 208350
rect 547026 208294 547094 208350
rect 547150 208294 547218 208350
rect 547274 208294 547342 208350
rect 547398 208294 564970 208350
rect 565026 208294 565094 208350
rect 565150 208294 565218 208350
rect 565274 208294 565342 208350
rect 565398 208294 582970 208350
rect 583026 208294 583094 208350
rect 583150 208294 583218 208350
rect 583274 208294 583342 208350
rect 583398 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 6970 208226
rect 7026 208170 7094 208226
rect 7150 208170 7218 208226
rect 7274 208170 7342 208226
rect 7398 208170 24970 208226
rect 25026 208170 25094 208226
rect 25150 208170 25218 208226
rect 25274 208170 25342 208226
rect 25398 208170 42970 208226
rect 43026 208170 43094 208226
rect 43150 208170 43218 208226
rect 43274 208170 43342 208226
rect 43398 208170 60970 208226
rect 61026 208170 61094 208226
rect 61150 208170 61218 208226
rect 61274 208170 61342 208226
rect 61398 208170 78970 208226
rect 79026 208170 79094 208226
rect 79150 208170 79218 208226
rect 79274 208170 79342 208226
rect 79398 208170 96970 208226
rect 97026 208170 97094 208226
rect 97150 208170 97218 208226
rect 97274 208170 97342 208226
rect 97398 208170 114970 208226
rect 115026 208170 115094 208226
rect 115150 208170 115218 208226
rect 115274 208170 115342 208226
rect 115398 208170 132970 208226
rect 133026 208170 133094 208226
rect 133150 208170 133218 208226
rect 133274 208170 133342 208226
rect 133398 208170 150970 208226
rect 151026 208170 151094 208226
rect 151150 208170 151218 208226
rect 151274 208170 151342 208226
rect 151398 208170 168970 208226
rect 169026 208170 169094 208226
rect 169150 208170 169218 208226
rect 169274 208170 169342 208226
rect 169398 208170 186970 208226
rect 187026 208170 187094 208226
rect 187150 208170 187218 208226
rect 187274 208170 187342 208226
rect 187398 208170 204970 208226
rect 205026 208170 205094 208226
rect 205150 208170 205218 208226
rect 205274 208170 205342 208226
rect 205398 208170 219878 208226
rect 219934 208170 220002 208226
rect 220058 208170 222970 208226
rect 223026 208170 223094 208226
rect 223150 208170 223218 208226
rect 223274 208170 223342 208226
rect 223398 208170 240970 208226
rect 241026 208170 241094 208226
rect 241150 208170 241218 208226
rect 241274 208170 241342 208226
rect 241398 208170 250598 208226
rect 250654 208170 250722 208226
rect 250778 208170 258970 208226
rect 259026 208170 259094 208226
rect 259150 208170 259218 208226
rect 259274 208170 259342 208226
rect 259398 208170 276970 208226
rect 277026 208170 277094 208226
rect 277150 208170 277218 208226
rect 277274 208170 277342 208226
rect 277398 208170 281318 208226
rect 281374 208170 281442 208226
rect 281498 208170 294970 208226
rect 295026 208170 295094 208226
rect 295150 208170 295218 208226
rect 295274 208170 295342 208226
rect 295398 208170 312038 208226
rect 312094 208170 312162 208226
rect 312218 208170 312970 208226
rect 313026 208170 313094 208226
rect 313150 208170 313218 208226
rect 313274 208170 313342 208226
rect 313398 208170 330970 208226
rect 331026 208170 331094 208226
rect 331150 208170 331218 208226
rect 331274 208170 331342 208226
rect 331398 208170 342758 208226
rect 342814 208170 342882 208226
rect 342938 208170 348970 208226
rect 349026 208170 349094 208226
rect 349150 208170 349218 208226
rect 349274 208170 349342 208226
rect 349398 208170 366970 208226
rect 367026 208170 367094 208226
rect 367150 208170 367218 208226
rect 367274 208170 367342 208226
rect 367398 208170 373478 208226
rect 373534 208170 373602 208226
rect 373658 208170 384970 208226
rect 385026 208170 385094 208226
rect 385150 208170 385218 208226
rect 385274 208170 385342 208226
rect 385398 208170 402970 208226
rect 403026 208170 403094 208226
rect 403150 208170 403218 208226
rect 403274 208170 403342 208226
rect 403398 208170 404198 208226
rect 404254 208170 404322 208226
rect 404378 208170 420970 208226
rect 421026 208170 421094 208226
rect 421150 208170 421218 208226
rect 421274 208170 421342 208226
rect 421398 208170 434918 208226
rect 434974 208170 435042 208226
rect 435098 208170 438970 208226
rect 439026 208170 439094 208226
rect 439150 208170 439218 208226
rect 439274 208170 439342 208226
rect 439398 208170 456970 208226
rect 457026 208170 457094 208226
rect 457150 208170 457218 208226
rect 457274 208170 457342 208226
rect 457398 208170 465638 208226
rect 465694 208170 465762 208226
rect 465818 208170 474970 208226
rect 475026 208170 475094 208226
rect 475150 208170 475218 208226
rect 475274 208170 475342 208226
rect 475398 208170 492970 208226
rect 493026 208170 493094 208226
rect 493150 208170 493218 208226
rect 493274 208170 493342 208226
rect 493398 208170 496358 208226
rect 496414 208170 496482 208226
rect 496538 208170 510970 208226
rect 511026 208170 511094 208226
rect 511150 208170 511218 208226
rect 511274 208170 511342 208226
rect 511398 208170 528970 208226
rect 529026 208170 529094 208226
rect 529150 208170 529218 208226
rect 529274 208170 529342 208226
rect 529398 208170 546970 208226
rect 547026 208170 547094 208226
rect 547150 208170 547218 208226
rect 547274 208170 547342 208226
rect 547398 208170 564970 208226
rect 565026 208170 565094 208226
rect 565150 208170 565218 208226
rect 565274 208170 565342 208226
rect 565398 208170 582970 208226
rect 583026 208170 583094 208226
rect 583150 208170 583218 208226
rect 583274 208170 583342 208226
rect 583398 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 6970 208102
rect 7026 208046 7094 208102
rect 7150 208046 7218 208102
rect 7274 208046 7342 208102
rect 7398 208046 24970 208102
rect 25026 208046 25094 208102
rect 25150 208046 25218 208102
rect 25274 208046 25342 208102
rect 25398 208046 42970 208102
rect 43026 208046 43094 208102
rect 43150 208046 43218 208102
rect 43274 208046 43342 208102
rect 43398 208046 60970 208102
rect 61026 208046 61094 208102
rect 61150 208046 61218 208102
rect 61274 208046 61342 208102
rect 61398 208046 78970 208102
rect 79026 208046 79094 208102
rect 79150 208046 79218 208102
rect 79274 208046 79342 208102
rect 79398 208046 96970 208102
rect 97026 208046 97094 208102
rect 97150 208046 97218 208102
rect 97274 208046 97342 208102
rect 97398 208046 114970 208102
rect 115026 208046 115094 208102
rect 115150 208046 115218 208102
rect 115274 208046 115342 208102
rect 115398 208046 132970 208102
rect 133026 208046 133094 208102
rect 133150 208046 133218 208102
rect 133274 208046 133342 208102
rect 133398 208046 150970 208102
rect 151026 208046 151094 208102
rect 151150 208046 151218 208102
rect 151274 208046 151342 208102
rect 151398 208046 168970 208102
rect 169026 208046 169094 208102
rect 169150 208046 169218 208102
rect 169274 208046 169342 208102
rect 169398 208046 186970 208102
rect 187026 208046 187094 208102
rect 187150 208046 187218 208102
rect 187274 208046 187342 208102
rect 187398 208046 204970 208102
rect 205026 208046 205094 208102
rect 205150 208046 205218 208102
rect 205274 208046 205342 208102
rect 205398 208046 219878 208102
rect 219934 208046 220002 208102
rect 220058 208046 222970 208102
rect 223026 208046 223094 208102
rect 223150 208046 223218 208102
rect 223274 208046 223342 208102
rect 223398 208046 240970 208102
rect 241026 208046 241094 208102
rect 241150 208046 241218 208102
rect 241274 208046 241342 208102
rect 241398 208046 250598 208102
rect 250654 208046 250722 208102
rect 250778 208046 258970 208102
rect 259026 208046 259094 208102
rect 259150 208046 259218 208102
rect 259274 208046 259342 208102
rect 259398 208046 276970 208102
rect 277026 208046 277094 208102
rect 277150 208046 277218 208102
rect 277274 208046 277342 208102
rect 277398 208046 281318 208102
rect 281374 208046 281442 208102
rect 281498 208046 294970 208102
rect 295026 208046 295094 208102
rect 295150 208046 295218 208102
rect 295274 208046 295342 208102
rect 295398 208046 312038 208102
rect 312094 208046 312162 208102
rect 312218 208046 312970 208102
rect 313026 208046 313094 208102
rect 313150 208046 313218 208102
rect 313274 208046 313342 208102
rect 313398 208046 330970 208102
rect 331026 208046 331094 208102
rect 331150 208046 331218 208102
rect 331274 208046 331342 208102
rect 331398 208046 342758 208102
rect 342814 208046 342882 208102
rect 342938 208046 348970 208102
rect 349026 208046 349094 208102
rect 349150 208046 349218 208102
rect 349274 208046 349342 208102
rect 349398 208046 366970 208102
rect 367026 208046 367094 208102
rect 367150 208046 367218 208102
rect 367274 208046 367342 208102
rect 367398 208046 373478 208102
rect 373534 208046 373602 208102
rect 373658 208046 384970 208102
rect 385026 208046 385094 208102
rect 385150 208046 385218 208102
rect 385274 208046 385342 208102
rect 385398 208046 402970 208102
rect 403026 208046 403094 208102
rect 403150 208046 403218 208102
rect 403274 208046 403342 208102
rect 403398 208046 404198 208102
rect 404254 208046 404322 208102
rect 404378 208046 420970 208102
rect 421026 208046 421094 208102
rect 421150 208046 421218 208102
rect 421274 208046 421342 208102
rect 421398 208046 434918 208102
rect 434974 208046 435042 208102
rect 435098 208046 438970 208102
rect 439026 208046 439094 208102
rect 439150 208046 439218 208102
rect 439274 208046 439342 208102
rect 439398 208046 456970 208102
rect 457026 208046 457094 208102
rect 457150 208046 457218 208102
rect 457274 208046 457342 208102
rect 457398 208046 465638 208102
rect 465694 208046 465762 208102
rect 465818 208046 474970 208102
rect 475026 208046 475094 208102
rect 475150 208046 475218 208102
rect 475274 208046 475342 208102
rect 475398 208046 492970 208102
rect 493026 208046 493094 208102
rect 493150 208046 493218 208102
rect 493274 208046 493342 208102
rect 493398 208046 496358 208102
rect 496414 208046 496482 208102
rect 496538 208046 510970 208102
rect 511026 208046 511094 208102
rect 511150 208046 511218 208102
rect 511274 208046 511342 208102
rect 511398 208046 528970 208102
rect 529026 208046 529094 208102
rect 529150 208046 529218 208102
rect 529274 208046 529342 208102
rect 529398 208046 546970 208102
rect 547026 208046 547094 208102
rect 547150 208046 547218 208102
rect 547274 208046 547342 208102
rect 547398 208046 564970 208102
rect 565026 208046 565094 208102
rect 565150 208046 565218 208102
rect 565274 208046 565342 208102
rect 565398 208046 582970 208102
rect 583026 208046 583094 208102
rect 583150 208046 583218 208102
rect 583274 208046 583342 208102
rect 583398 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 6970 207978
rect 7026 207922 7094 207978
rect 7150 207922 7218 207978
rect 7274 207922 7342 207978
rect 7398 207922 24970 207978
rect 25026 207922 25094 207978
rect 25150 207922 25218 207978
rect 25274 207922 25342 207978
rect 25398 207922 42970 207978
rect 43026 207922 43094 207978
rect 43150 207922 43218 207978
rect 43274 207922 43342 207978
rect 43398 207922 60970 207978
rect 61026 207922 61094 207978
rect 61150 207922 61218 207978
rect 61274 207922 61342 207978
rect 61398 207922 78970 207978
rect 79026 207922 79094 207978
rect 79150 207922 79218 207978
rect 79274 207922 79342 207978
rect 79398 207922 96970 207978
rect 97026 207922 97094 207978
rect 97150 207922 97218 207978
rect 97274 207922 97342 207978
rect 97398 207922 114970 207978
rect 115026 207922 115094 207978
rect 115150 207922 115218 207978
rect 115274 207922 115342 207978
rect 115398 207922 132970 207978
rect 133026 207922 133094 207978
rect 133150 207922 133218 207978
rect 133274 207922 133342 207978
rect 133398 207922 150970 207978
rect 151026 207922 151094 207978
rect 151150 207922 151218 207978
rect 151274 207922 151342 207978
rect 151398 207922 168970 207978
rect 169026 207922 169094 207978
rect 169150 207922 169218 207978
rect 169274 207922 169342 207978
rect 169398 207922 186970 207978
rect 187026 207922 187094 207978
rect 187150 207922 187218 207978
rect 187274 207922 187342 207978
rect 187398 207922 204970 207978
rect 205026 207922 205094 207978
rect 205150 207922 205218 207978
rect 205274 207922 205342 207978
rect 205398 207922 219878 207978
rect 219934 207922 220002 207978
rect 220058 207922 222970 207978
rect 223026 207922 223094 207978
rect 223150 207922 223218 207978
rect 223274 207922 223342 207978
rect 223398 207922 240970 207978
rect 241026 207922 241094 207978
rect 241150 207922 241218 207978
rect 241274 207922 241342 207978
rect 241398 207922 250598 207978
rect 250654 207922 250722 207978
rect 250778 207922 258970 207978
rect 259026 207922 259094 207978
rect 259150 207922 259218 207978
rect 259274 207922 259342 207978
rect 259398 207922 276970 207978
rect 277026 207922 277094 207978
rect 277150 207922 277218 207978
rect 277274 207922 277342 207978
rect 277398 207922 281318 207978
rect 281374 207922 281442 207978
rect 281498 207922 294970 207978
rect 295026 207922 295094 207978
rect 295150 207922 295218 207978
rect 295274 207922 295342 207978
rect 295398 207922 312038 207978
rect 312094 207922 312162 207978
rect 312218 207922 312970 207978
rect 313026 207922 313094 207978
rect 313150 207922 313218 207978
rect 313274 207922 313342 207978
rect 313398 207922 330970 207978
rect 331026 207922 331094 207978
rect 331150 207922 331218 207978
rect 331274 207922 331342 207978
rect 331398 207922 342758 207978
rect 342814 207922 342882 207978
rect 342938 207922 348970 207978
rect 349026 207922 349094 207978
rect 349150 207922 349218 207978
rect 349274 207922 349342 207978
rect 349398 207922 366970 207978
rect 367026 207922 367094 207978
rect 367150 207922 367218 207978
rect 367274 207922 367342 207978
rect 367398 207922 373478 207978
rect 373534 207922 373602 207978
rect 373658 207922 384970 207978
rect 385026 207922 385094 207978
rect 385150 207922 385218 207978
rect 385274 207922 385342 207978
rect 385398 207922 402970 207978
rect 403026 207922 403094 207978
rect 403150 207922 403218 207978
rect 403274 207922 403342 207978
rect 403398 207922 404198 207978
rect 404254 207922 404322 207978
rect 404378 207922 420970 207978
rect 421026 207922 421094 207978
rect 421150 207922 421218 207978
rect 421274 207922 421342 207978
rect 421398 207922 434918 207978
rect 434974 207922 435042 207978
rect 435098 207922 438970 207978
rect 439026 207922 439094 207978
rect 439150 207922 439218 207978
rect 439274 207922 439342 207978
rect 439398 207922 456970 207978
rect 457026 207922 457094 207978
rect 457150 207922 457218 207978
rect 457274 207922 457342 207978
rect 457398 207922 465638 207978
rect 465694 207922 465762 207978
rect 465818 207922 474970 207978
rect 475026 207922 475094 207978
rect 475150 207922 475218 207978
rect 475274 207922 475342 207978
rect 475398 207922 492970 207978
rect 493026 207922 493094 207978
rect 493150 207922 493218 207978
rect 493274 207922 493342 207978
rect 493398 207922 496358 207978
rect 496414 207922 496482 207978
rect 496538 207922 510970 207978
rect 511026 207922 511094 207978
rect 511150 207922 511218 207978
rect 511274 207922 511342 207978
rect 511398 207922 528970 207978
rect 529026 207922 529094 207978
rect 529150 207922 529218 207978
rect 529274 207922 529342 207978
rect 529398 207922 546970 207978
rect 547026 207922 547094 207978
rect 547150 207922 547218 207978
rect 547274 207922 547342 207978
rect 547398 207922 564970 207978
rect 565026 207922 565094 207978
rect 565150 207922 565218 207978
rect 565274 207922 565342 207978
rect 565398 207922 582970 207978
rect 583026 207922 583094 207978
rect 583150 207922 583218 207978
rect 583274 207922 583342 207978
rect 583398 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 3250 202350
rect 3306 202294 3374 202350
rect 3430 202294 3498 202350
rect 3554 202294 3622 202350
rect 3678 202294 21250 202350
rect 21306 202294 21374 202350
rect 21430 202294 21498 202350
rect 21554 202294 21622 202350
rect 21678 202294 39250 202350
rect 39306 202294 39374 202350
rect 39430 202294 39498 202350
rect 39554 202294 39622 202350
rect 39678 202294 57250 202350
rect 57306 202294 57374 202350
rect 57430 202294 57498 202350
rect 57554 202294 57622 202350
rect 57678 202294 75250 202350
rect 75306 202294 75374 202350
rect 75430 202294 75498 202350
rect 75554 202294 75622 202350
rect 75678 202294 93250 202350
rect 93306 202294 93374 202350
rect 93430 202294 93498 202350
rect 93554 202294 93622 202350
rect 93678 202294 111250 202350
rect 111306 202294 111374 202350
rect 111430 202294 111498 202350
rect 111554 202294 111622 202350
rect 111678 202294 129250 202350
rect 129306 202294 129374 202350
rect 129430 202294 129498 202350
rect 129554 202294 129622 202350
rect 129678 202294 147250 202350
rect 147306 202294 147374 202350
rect 147430 202294 147498 202350
rect 147554 202294 147622 202350
rect 147678 202294 165250 202350
rect 165306 202294 165374 202350
rect 165430 202294 165498 202350
rect 165554 202294 165622 202350
rect 165678 202294 183250 202350
rect 183306 202294 183374 202350
rect 183430 202294 183498 202350
rect 183554 202294 183622 202350
rect 183678 202294 201250 202350
rect 201306 202294 201374 202350
rect 201430 202294 201498 202350
rect 201554 202294 201622 202350
rect 201678 202294 237250 202350
rect 237306 202294 237374 202350
rect 237430 202294 237498 202350
rect 237554 202294 237622 202350
rect 237678 202294 255250 202350
rect 255306 202294 255374 202350
rect 255430 202294 255498 202350
rect 255554 202294 255622 202350
rect 255678 202294 273250 202350
rect 273306 202294 273374 202350
rect 273430 202294 273498 202350
rect 273554 202294 273622 202350
rect 273678 202294 291250 202350
rect 291306 202294 291374 202350
rect 291430 202294 291498 202350
rect 291554 202294 291622 202350
rect 291678 202294 309250 202350
rect 309306 202294 309374 202350
rect 309430 202294 309498 202350
rect 309554 202294 309622 202350
rect 309678 202294 345250 202350
rect 345306 202294 345374 202350
rect 345430 202294 345498 202350
rect 345554 202294 345622 202350
rect 345678 202294 363250 202350
rect 363306 202294 363374 202350
rect 363430 202294 363498 202350
rect 363554 202294 363622 202350
rect 363678 202294 381250 202350
rect 381306 202294 381374 202350
rect 381430 202294 381498 202350
rect 381554 202294 381622 202350
rect 381678 202294 399250 202350
rect 399306 202294 399374 202350
rect 399430 202294 399498 202350
rect 399554 202294 399622 202350
rect 399678 202294 417250 202350
rect 417306 202294 417374 202350
rect 417430 202294 417498 202350
rect 417554 202294 417622 202350
rect 417678 202294 453250 202350
rect 453306 202294 453374 202350
rect 453430 202294 453498 202350
rect 453554 202294 453622 202350
rect 453678 202294 471250 202350
rect 471306 202294 471374 202350
rect 471430 202294 471498 202350
rect 471554 202294 471622 202350
rect 471678 202294 489250 202350
rect 489306 202294 489374 202350
rect 489430 202294 489498 202350
rect 489554 202294 489622 202350
rect 489678 202294 507250 202350
rect 507306 202294 507374 202350
rect 507430 202294 507498 202350
rect 507554 202294 507622 202350
rect 507678 202294 525250 202350
rect 525306 202294 525374 202350
rect 525430 202294 525498 202350
rect 525554 202294 525622 202350
rect 525678 202294 543250 202350
rect 543306 202294 543374 202350
rect 543430 202294 543498 202350
rect 543554 202294 543622 202350
rect 543678 202294 561250 202350
rect 561306 202294 561374 202350
rect 561430 202294 561498 202350
rect 561554 202294 561622 202350
rect 561678 202294 579250 202350
rect 579306 202294 579374 202350
rect 579430 202294 579498 202350
rect 579554 202294 579622 202350
rect 579678 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 3250 202226
rect 3306 202170 3374 202226
rect 3430 202170 3498 202226
rect 3554 202170 3622 202226
rect 3678 202170 21250 202226
rect 21306 202170 21374 202226
rect 21430 202170 21498 202226
rect 21554 202170 21622 202226
rect 21678 202170 39250 202226
rect 39306 202170 39374 202226
rect 39430 202170 39498 202226
rect 39554 202170 39622 202226
rect 39678 202170 57250 202226
rect 57306 202170 57374 202226
rect 57430 202170 57498 202226
rect 57554 202170 57622 202226
rect 57678 202170 75250 202226
rect 75306 202170 75374 202226
rect 75430 202170 75498 202226
rect 75554 202170 75622 202226
rect 75678 202170 93250 202226
rect 93306 202170 93374 202226
rect 93430 202170 93498 202226
rect 93554 202170 93622 202226
rect 93678 202170 111250 202226
rect 111306 202170 111374 202226
rect 111430 202170 111498 202226
rect 111554 202170 111622 202226
rect 111678 202170 129250 202226
rect 129306 202170 129374 202226
rect 129430 202170 129498 202226
rect 129554 202170 129622 202226
rect 129678 202170 147250 202226
rect 147306 202170 147374 202226
rect 147430 202170 147498 202226
rect 147554 202170 147622 202226
rect 147678 202170 165250 202226
rect 165306 202170 165374 202226
rect 165430 202170 165498 202226
rect 165554 202170 165622 202226
rect 165678 202170 183250 202226
rect 183306 202170 183374 202226
rect 183430 202170 183498 202226
rect 183554 202170 183622 202226
rect 183678 202170 201250 202226
rect 201306 202170 201374 202226
rect 201430 202170 201498 202226
rect 201554 202170 201622 202226
rect 201678 202170 237250 202226
rect 237306 202170 237374 202226
rect 237430 202170 237498 202226
rect 237554 202170 237622 202226
rect 237678 202170 255250 202226
rect 255306 202170 255374 202226
rect 255430 202170 255498 202226
rect 255554 202170 255622 202226
rect 255678 202170 273250 202226
rect 273306 202170 273374 202226
rect 273430 202170 273498 202226
rect 273554 202170 273622 202226
rect 273678 202170 291250 202226
rect 291306 202170 291374 202226
rect 291430 202170 291498 202226
rect 291554 202170 291622 202226
rect 291678 202170 309250 202226
rect 309306 202170 309374 202226
rect 309430 202170 309498 202226
rect 309554 202170 309622 202226
rect 309678 202170 345250 202226
rect 345306 202170 345374 202226
rect 345430 202170 345498 202226
rect 345554 202170 345622 202226
rect 345678 202170 363250 202226
rect 363306 202170 363374 202226
rect 363430 202170 363498 202226
rect 363554 202170 363622 202226
rect 363678 202170 381250 202226
rect 381306 202170 381374 202226
rect 381430 202170 381498 202226
rect 381554 202170 381622 202226
rect 381678 202170 399250 202226
rect 399306 202170 399374 202226
rect 399430 202170 399498 202226
rect 399554 202170 399622 202226
rect 399678 202170 417250 202226
rect 417306 202170 417374 202226
rect 417430 202170 417498 202226
rect 417554 202170 417622 202226
rect 417678 202170 453250 202226
rect 453306 202170 453374 202226
rect 453430 202170 453498 202226
rect 453554 202170 453622 202226
rect 453678 202170 471250 202226
rect 471306 202170 471374 202226
rect 471430 202170 471498 202226
rect 471554 202170 471622 202226
rect 471678 202170 489250 202226
rect 489306 202170 489374 202226
rect 489430 202170 489498 202226
rect 489554 202170 489622 202226
rect 489678 202170 507250 202226
rect 507306 202170 507374 202226
rect 507430 202170 507498 202226
rect 507554 202170 507622 202226
rect 507678 202170 525250 202226
rect 525306 202170 525374 202226
rect 525430 202170 525498 202226
rect 525554 202170 525622 202226
rect 525678 202170 543250 202226
rect 543306 202170 543374 202226
rect 543430 202170 543498 202226
rect 543554 202170 543622 202226
rect 543678 202170 561250 202226
rect 561306 202170 561374 202226
rect 561430 202170 561498 202226
rect 561554 202170 561622 202226
rect 561678 202170 579250 202226
rect 579306 202170 579374 202226
rect 579430 202170 579498 202226
rect 579554 202170 579622 202226
rect 579678 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 3250 202102
rect 3306 202046 3374 202102
rect 3430 202046 3498 202102
rect 3554 202046 3622 202102
rect 3678 202046 21250 202102
rect 21306 202046 21374 202102
rect 21430 202046 21498 202102
rect 21554 202046 21622 202102
rect 21678 202046 39250 202102
rect 39306 202046 39374 202102
rect 39430 202046 39498 202102
rect 39554 202046 39622 202102
rect 39678 202046 57250 202102
rect 57306 202046 57374 202102
rect 57430 202046 57498 202102
rect 57554 202046 57622 202102
rect 57678 202046 75250 202102
rect 75306 202046 75374 202102
rect 75430 202046 75498 202102
rect 75554 202046 75622 202102
rect 75678 202046 93250 202102
rect 93306 202046 93374 202102
rect 93430 202046 93498 202102
rect 93554 202046 93622 202102
rect 93678 202046 111250 202102
rect 111306 202046 111374 202102
rect 111430 202046 111498 202102
rect 111554 202046 111622 202102
rect 111678 202046 129250 202102
rect 129306 202046 129374 202102
rect 129430 202046 129498 202102
rect 129554 202046 129622 202102
rect 129678 202046 147250 202102
rect 147306 202046 147374 202102
rect 147430 202046 147498 202102
rect 147554 202046 147622 202102
rect 147678 202046 165250 202102
rect 165306 202046 165374 202102
rect 165430 202046 165498 202102
rect 165554 202046 165622 202102
rect 165678 202046 183250 202102
rect 183306 202046 183374 202102
rect 183430 202046 183498 202102
rect 183554 202046 183622 202102
rect 183678 202046 201250 202102
rect 201306 202046 201374 202102
rect 201430 202046 201498 202102
rect 201554 202046 201622 202102
rect 201678 202046 237250 202102
rect 237306 202046 237374 202102
rect 237430 202046 237498 202102
rect 237554 202046 237622 202102
rect 237678 202046 255250 202102
rect 255306 202046 255374 202102
rect 255430 202046 255498 202102
rect 255554 202046 255622 202102
rect 255678 202046 273250 202102
rect 273306 202046 273374 202102
rect 273430 202046 273498 202102
rect 273554 202046 273622 202102
rect 273678 202046 291250 202102
rect 291306 202046 291374 202102
rect 291430 202046 291498 202102
rect 291554 202046 291622 202102
rect 291678 202046 309250 202102
rect 309306 202046 309374 202102
rect 309430 202046 309498 202102
rect 309554 202046 309622 202102
rect 309678 202046 345250 202102
rect 345306 202046 345374 202102
rect 345430 202046 345498 202102
rect 345554 202046 345622 202102
rect 345678 202046 363250 202102
rect 363306 202046 363374 202102
rect 363430 202046 363498 202102
rect 363554 202046 363622 202102
rect 363678 202046 381250 202102
rect 381306 202046 381374 202102
rect 381430 202046 381498 202102
rect 381554 202046 381622 202102
rect 381678 202046 399250 202102
rect 399306 202046 399374 202102
rect 399430 202046 399498 202102
rect 399554 202046 399622 202102
rect 399678 202046 417250 202102
rect 417306 202046 417374 202102
rect 417430 202046 417498 202102
rect 417554 202046 417622 202102
rect 417678 202046 453250 202102
rect 453306 202046 453374 202102
rect 453430 202046 453498 202102
rect 453554 202046 453622 202102
rect 453678 202046 471250 202102
rect 471306 202046 471374 202102
rect 471430 202046 471498 202102
rect 471554 202046 471622 202102
rect 471678 202046 489250 202102
rect 489306 202046 489374 202102
rect 489430 202046 489498 202102
rect 489554 202046 489622 202102
rect 489678 202046 507250 202102
rect 507306 202046 507374 202102
rect 507430 202046 507498 202102
rect 507554 202046 507622 202102
rect 507678 202046 525250 202102
rect 525306 202046 525374 202102
rect 525430 202046 525498 202102
rect 525554 202046 525622 202102
rect 525678 202046 543250 202102
rect 543306 202046 543374 202102
rect 543430 202046 543498 202102
rect 543554 202046 543622 202102
rect 543678 202046 561250 202102
rect 561306 202046 561374 202102
rect 561430 202046 561498 202102
rect 561554 202046 561622 202102
rect 561678 202046 579250 202102
rect 579306 202046 579374 202102
rect 579430 202046 579498 202102
rect 579554 202046 579622 202102
rect 579678 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 3250 201978
rect 3306 201922 3374 201978
rect 3430 201922 3498 201978
rect 3554 201922 3622 201978
rect 3678 201922 21250 201978
rect 21306 201922 21374 201978
rect 21430 201922 21498 201978
rect 21554 201922 21622 201978
rect 21678 201922 39250 201978
rect 39306 201922 39374 201978
rect 39430 201922 39498 201978
rect 39554 201922 39622 201978
rect 39678 201922 57250 201978
rect 57306 201922 57374 201978
rect 57430 201922 57498 201978
rect 57554 201922 57622 201978
rect 57678 201922 75250 201978
rect 75306 201922 75374 201978
rect 75430 201922 75498 201978
rect 75554 201922 75622 201978
rect 75678 201922 93250 201978
rect 93306 201922 93374 201978
rect 93430 201922 93498 201978
rect 93554 201922 93622 201978
rect 93678 201922 111250 201978
rect 111306 201922 111374 201978
rect 111430 201922 111498 201978
rect 111554 201922 111622 201978
rect 111678 201922 129250 201978
rect 129306 201922 129374 201978
rect 129430 201922 129498 201978
rect 129554 201922 129622 201978
rect 129678 201922 147250 201978
rect 147306 201922 147374 201978
rect 147430 201922 147498 201978
rect 147554 201922 147622 201978
rect 147678 201922 165250 201978
rect 165306 201922 165374 201978
rect 165430 201922 165498 201978
rect 165554 201922 165622 201978
rect 165678 201922 183250 201978
rect 183306 201922 183374 201978
rect 183430 201922 183498 201978
rect 183554 201922 183622 201978
rect 183678 201922 201250 201978
rect 201306 201922 201374 201978
rect 201430 201922 201498 201978
rect 201554 201922 201622 201978
rect 201678 201922 237250 201978
rect 237306 201922 237374 201978
rect 237430 201922 237498 201978
rect 237554 201922 237622 201978
rect 237678 201922 255250 201978
rect 255306 201922 255374 201978
rect 255430 201922 255498 201978
rect 255554 201922 255622 201978
rect 255678 201922 273250 201978
rect 273306 201922 273374 201978
rect 273430 201922 273498 201978
rect 273554 201922 273622 201978
rect 273678 201922 291250 201978
rect 291306 201922 291374 201978
rect 291430 201922 291498 201978
rect 291554 201922 291622 201978
rect 291678 201922 309250 201978
rect 309306 201922 309374 201978
rect 309430 201922 309498 201978
rect 309554 201922 309622 201978
rect 309678 201922 345250 201978
rect 345306 201922 345374 201978
rect 345430 201922 345498 201978
rect 345554 201922 345622 201978
rect 345678 201922 363250 201978
rect 363306 201922 363374 201978
rect 363430 201922 363498 201978
rect 363554 201922 363622 201978
rect 363678 201922 381250 201978
rect 381306 201922 381374 201978
rect 381430 201922 381498 201978
rect 381554 201922 381622 201978
rect 381678 201922 399250 201978
rect 399306 201922 399374 201978
rect 399430 201922 399498 201978
rect 399554 201922 399622 201978
rect 399678 201922 417250 201978
rect 417306 201922 417374 201978
rect 417430 201922 417498 201978
rect 417554 201922 417622 201978
rect 417678 201922 453250 201978
rect 453306 201922 453374 201978
rect 453430 201922 453498 201978
rect 453554 201922 453622 201978
rect 453678 201922 471250 201978
rect 471306 201922 471374 201978
rect 471430 201922 471498 201978
rect 471554 201922 471622 201978
rect 471678 201922 489250 201978
rect 489306 201922 489374 201978
rect 489430 201922 489498 201978
rect 489554 201922 489622 201978
rect 489678 201922 507250 201978
rect 507306 201922 507374 201978
rect 507430 201922 507498 201978
rect 507554 201922 507622 201978
rect 507678 201922 525250 201978
rect 525306 201922 525374 201978
rect 525430 201922 525498 201978
rect 525554 201922 525622 201978
rect 525678 201922 543250 201978
rect 543306 201922 543374 201978
rect 543430 201922 543498 201978
rect 543554 201922 543622 201978
rect 543678 201922 561250 201978
rect 561306 201922 561374 201978
rect 561430 201922 561498 201978
rect 561554 201922 561622 201978
rect 561678 201922 579250 201978
rect 579306 201922 579374 201978
rect 579430 201922 579498 201978
rect 579554 201922 579622 201978
rect 579678 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 6970 190350
rect 7026 190294 7094 190350
rect 7150 190294 7218 190350
rect 7274 190294 7342 190350
rect 7398 190294 24970 190350
rect 25026 190294 25094 190350
rect 25150 190294 25218 190350
rect 25274 190294 25342 190350
rect 25398 190294 42970 190350
rect 43026 190294 43094 190350
rect 43150 190294 43218 190350
rect 43274 190294 43342 190350
rect 43398 190294 60970 190350
rect 61026 190294 61094 190350
rect 61150 190294 61218 190350
rect 61274 190294 61342 190350
rect 61398 190294 78970 190350
rect 79026 190294 79094 190350
rect 79150 190294 79218 190350
rect 79274 190294 79342 190350
rect 79398 190294 96970 190350
rect 97026 190294 97094 190350
rect 97150 190294 97218 190350
rect 97274 190294 97342 190350
rect 97398 190294 114970 190350
rect 115026 190294 115094 190350
rect 115150 190294 115218 190350
rect 115274 190294 115342 190350
rect 115398 190294 132970 190350
rect 133026 190294 133094 190350
rect 133150 190294 133218 190350
rect 133274 190294 133342 190350
rect 133398 190294 150970 190350
rect 151026 190294 151094 190350
rect 151150 190294 151218 190350
rect 151274 190294 151342 190350
rect 151398 190294 168970 190350
rect 169026 190294 169094 190350
rect 169150 190294 169218 190350
rect 169274 190294 169342 190350
rect 169398 190294 186970 190350
rect 187026 190294 187094 190350
rect 187150 190294 187218 190350
rect 187274 190294 187342 190350
rect 187398 190294 204970 190350
rect 205026 190294 205094 190350
rect 205150 190294 205218 190350
rect 205274 190294 205342 190350
rect 205398 190294 222970 190350
rect 223026 190294 223094 190350
rect 223150 190294 223218 190350
rect 223274 190294 223342 190350
rect 223398 190294 240970 190350
rect 241026 190294 241094 190350
rect 241150 190294 241218 190350
rect 241274 190294 241342 190350
rect 241398 190294 258970 190350
rect 259026 190294 259094 190350
rect 259150 190294 259218 190350
rect 259274 190294 259342 190350
rect 259398 190294 276970 190350
rect 277026 190294 277094 190350
rect 277150 190294 277218 190350
rect 277274 190294 277342 190350
rect 277398 190294 294970 190350
rect 295026 190294 295094 190350
rect 295150 190294 295218 190350
rect 295274 190294 295342 190350
rect 295398 190294 312970 190350
rect 313026 190294 313094 190350
rect 313150 190294 313218 190350
rect 313274 190294 313342 190350
rect 313398 190294 330970 190350
rect 331026 190294 331094 190350
rect 331150 190294 331218 190350
rect 331274 190294 331342 190350
rect 331398 190294 348970 190350
rect 349026 190294 349094 190350
rect 349150 190294 349218 190350
rect 349274 190294 349342 190350
rect 349398 190294 366970 190350
rect 367026 190294 367094 190350
rect 367150 190294 367218 190350
rect 367274 190294 367342 190350
rect 367398 190294 384970 190350
rect 385026 190294 385094 190350
rect 385150 190294 385218 190350
rect 385274 190294 385342 190350
rect 385398 190294 402970 190350
rect 403026 190294 403094 190350
rect 403150 190294 403218 190350
rect 403274 190294 403342 190350
rect 403398 190294 420970 190350
rect 421026 190294 421094 190350
rect 421150 190294 421218 190350
rect 421274 190294 421342 190350
rect 421398 190294 438970 190350
rect 439026 190294 439094 190350
rect 439150 190294 439218 190350
rect 439274 190294 439342 190350
rect 439398 190294 456970 190350
rect 457026 190294 457094 190350
rect 457150 190294 457218 190350
rect 457274 190294 457342 190350
rect 457398 190294 474970 190350
rect 475026 190294 475094 190350
rect 475150 190294 475218 190350
rect 475274 190294 475342 190350
rect 475398 190294 492970 190350
rect 493026 190294 493094 190350
rect 493150 190294 493218 190350
rect 493274 190294 493342 190350
rect 493398 190294 510970 190350
rect 511026 190294 511094 190350
rect 511150 190294 511218 190350
rect 511274 190294 511342 190350
rect 511398 190294 528970 190350
rect 529026 190294 529094 190350
rect 529150 190294 529218 190350
rect 529274 190294 529342 190350
rect 529398 190294 546970 190350
rect 547026 190294 547094 190350
rect 547150 190294 547218 190350
rect 547274 190294 547342 190350
rect 547398 190294 564970 190350
rect 565026 190294 565094 190350
rect 565150 190294 565218 190350
rect 565274 190294 565342 190350
rect 565398 190294 582970 190350
rect 583026 190294 583094 190350
rect 583150 190294 583218 190350
rect 583274 190294 583342 190350
rect 583398 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 6970 190226
rect 7026 190170 7094 190226
rect 7150 190170 7218 190226
rect 7274 190170 7342 190226
rect 7398 190170 24970 190226
rect 25026 190170 25094 190226
rect 25150 190170 25218 190226
rect 25274 190170 25342 190226
rect 25398 190170 42970 190226
rect 43026 190170 43094 190226
rect 43150 190170 43218 190226
rect 43274 190170 43342 190226
rect 43398 190170 60970 190226
rect 61026 190170 61094 190226
rect 61150 190170 61218 190226
rect 61274 190170 61342 190226
rect 61398 190170 78970 190226
rect 79026 190170 79094 190226
rect 79150 190170 79218 190226
rect 79274 190170 79342 190226
rect 79398 190170 96970 190226
rect 97026 190170 97094 190226
rect 97150 190170 97218 190226
rect 97274 190170 97342 190226
rect 97398 190170 114970 190226
rect 115026 190170 115094 190226
rect 115150 190170 115218 190226
rect 115274 190170 115342 190226
rect 115398 190170 132970 190226
rect 133026 190170 133094 190226
rect 133150 190170 133218 190226
rect 133274 190170 133342 190226
rect 133398 190170 150970 190226
rect 151026 190170 151094 190226
rect 151150 190170 151218 190226
rect 151274 190170 151342 190226
rect 151398 190170 168970 190226
rect 169026 190170 169094 190226
rect 169150 190170 169218 190226
rect 169274 190170 169342 190226
rect 169398 190170 186970 190226
rect 187026 190170 187094 190226
rect 187150 190170 187218 190226
rect 187274 190170 187342 190226
rect 187398 190170 204970 190226
rect 205026 190170 205094 190226
rect 205150 190170 205218 190226
rect 205274 190170 205342 190226
rect 205398 190170 222970 190226
rect 223026 190170 223094 190226
rect 223150 190170 223218 190226
rect 223274 190170 223342 190226
rect 223398 190170 240970 190226
rect 241026 190170 241094 190226
rect 241150 190170 241218 190226
rect 241274 190170 241342 190226
rect 241398 190170 258970 190226
rect 259026 190170 259094 190226
rect 259150 190170 259218 190226
rect 259274 190170 259342 190226
rect 259398 190170 276970 190226
rect 277026 190170 277094 190226
rect 277150 190170 277218 190226
rect 277274 190170 277342 190226
rect 277398 190170 294970 190226
rect 295026 190170 295094 190226
rect 295150 190170 295218 190226
rect 295274 190170 295342 190226
rect 295398 190170 312970 190226
rect 313026 190170 313094 190226
rect 313150 190170 313218 190226
rect 313274 190170 313342 190226
rect 313398 190170 330970 190226
rect 331026 190170 331094 190226
rect 331150 190170 331218 190226
rect 331274 190170 331342 190226
rect 331398 190170 348970 190226
rect 349026 190170 349094 190226
rect 349150 190170 349218 190226
rect 349274 190170 349342 190226
rect 349398 190170 366970 190226
rect 367026 190170 367094 190226
rect 367150 190170 367218 190226
rect 367274 190170 367342 190226
rect 367398 190170 384970 190226
rect 385026 190170 385094 190226
rect 385150 190170 385218 190226
rect 385274 190170 385342 190226
rect 385398 190170 402970 190226
rect 403026 190170 403094 190226
rect 403150 190170 403218 190226
rect 403274 190170 403342 190226
rect 403398 190170 420970 190226
rect 421026 190170 421094 190226
rect 421150 190170 421218 190226
rect 421274 190170 421342 190226
rect 421398 190170 438970 190226
rect 439026 190170 439094 190226
rect 439150 190170 439218 190226
rect 439274 190170 439342 190226
rect 439398 190170 456970 190226
rect 457026 190170 457094 190226
rect 457150 190170 457218 190226
rect 457274 190170 457342 190226
rect 457398 190170 474970 190226
rect 475026 190170 475094 190226
rect 475150 190170 475218 190226
rect 475274 190170 475342 190226
rect 475398 190170 492970 190226
rect 493026 190170 493094 190226
rect 493150 190170 493218 190226
rect 493274 190170 493342 190226
rect 493398 190170 510970 190226
rect 511026 190170 511094 190226
rect 511150 190170 511218 190226
rect 511274 190170 511342 190226
rect 511398 190170 528970 190226
rect 529026 190170 529094 190226
rect 529150 190170 529218 190226
rect 529274 190170 529342 190226
rect 529398 190170 546970 190226
rect 547026 190170 547094 190226
rect 547150 190170 547218 190226
rect 547274 190170 547342 190226
rect 547398 190170 564970 190226
rect 565026 190170 565094 190226
rect 565150 190170 565218 190226
rect 565274 190170 565342 190226
rect 565398 190170 582970 190226
rect 583026 190170 583094 190226
rect 583150 190170 583218 190226
rect 583274 190170 583342 190226
rect 583398 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 6970 190102
rect 7026 190046 7094 190102
rect 7150 190046 7218 190102
rect 7274 190046 7342 190102
rect 7398 190046 24970 190102
rect 25026 190046 25094 190102
rect 25150 190046 25218 190102
rect 25274 190046 25342 190102
rect 25398 190046 42970 190102
rect 43026 190046 43094 190102
rect 43150 190046 43218 190102
rect 43274 190046 43342 190102
rect 43398 190046 60970 190102
rect 61026 190046 61094 190102
rect 61150 190046 61218 190102
rect 61274 190046 61342 190102
rect 61398 190046 78970 190102
rect 79026 190046 79094 190102
rect 79150 190046 79218 190102
rect 79274 190046 79342 190102
rect 79398 190046 96970 190102
rect 97026 190046 97094 190102
rect 97150 190046 97218 190102
rect 97274 190046 97342 190102
rect 97398 190046 114970 190102
rect 115026 190046 115094 190102
rect 115150 190046 115218 190102
rect 115274 190046 115342 190102
rect 115398 190046 132970 190102
rect 133026 190046 133094 190102
rect 133150 190046 133218 190102
rect 133274 190046 133342 190102
rect 133398 190046 150970 190102
rect 151026 190046 151094 190102
rect 151150 190046 151218 190102
rect 151274 190046 151342 190102
rect 151398 190046 168970 190102
rect 169026 190046 169094 190102
rect 169150 190046 169218 190102
rect 169274 190046 169342 190102
rect 169398 190046 186970 190102
rect 187026 190046 187094 190102
rect 187150 190046 187218 190102
rect 187274 190046 187342 190102
rect 187398 190046 204970 190102
rect 205026 190046 205094 190102
rect 205150 190046 205218 190102
rect 205274 190046 205342 190102
rect 205398 190046 222970 190102
rect 223026 190046 223094 190102
rect 223150 190046 223218 190102
rect 223274 190046 223342 190102
rect 223398 190046 240970 190102
rect 241026 190046 241094 190102
rect 241150 190046 241218 190102
rect 241274 190046 241342 190102
rect 241398 190046 258970 190102
rect 259026 190046 259094 190102
rect 259150 190046 259218 190102
rect 259274 190046 259342 190102
rect 259398 190046 276970 190102
rect 277026 190046 277094 190102
rect 277150 190046 277218 190102
rect 277274 190046 277342 190102
rect 277398 190046 294970 190102
rect 295026 190046 295094 190102
rect 295150 190046 295218 190102
rect 295274 190046 295342 190102
rect 295398 190046 312970 190102
rect 313026 190046 313094 190102
rect 313150 190046 313218 190102
rect 313274 190046 313342 190102
rect 313398 190046 330970 190102
rect 331026 190046 331094 190102
rect 331150 190046 331218 190102
rect 331274 190046 331342 190102
rect 331398 190046 348970 190102
rect 349026 190046 349094 190102
rect 349150 190046 349218 190102
rect 349274 190046 349342 190102
rect 349398 190046 366970 190102
rect 367026 190046 367094 190102
rect 367150 190046 367218 190102
rect 367274 190046 367342 190102
rect 367398 190046 384970 190102
rect 385026 190046 385094 190102
rect 385150 190046 385218 190102
rect 385274 190046 385342 190102
rect 385398 190046 402970 190102
rect 403026 190046 403094 190102
rect 403150 190046 403218 190102
rect 403274 190046 403342 190102
rect 403398 190046 420970 190102
rect 421026 190046 421094 190102
rect 421150 190046 421218 190102
rect 421274 190046 421342 190102
rect 421398 190046 438970 190102
rect 439026 190046 439094 190102
rect 439150 190046 439218 190102
rect 439274 190046 439342 190102
rect 439398 190046 456970 190102
rect 457026 190046 457094 190102
rect 457150 190046 457218 190102
rect 457274 190046 457342 190102
rect 457398 190046 474970 190102
rect 475026 190046 475094 190102
rect 475150 190046 475218 190102
rect 475274 190046 475342 190102
rect 475398 190046 492970 190102
rect 493026 190046 493094 190102
rect 493150 190046 493218 190102
rect 493274 190046 493342 190102
rect 493398 190046 510970 190102
rect 511026 190046 511094 190102
rect 511150 190046 511218 190102
rect 511274 190046 511342 190102
rect 511398 190046 528970 190102
rect 529026 190046 529094 190102
rect 529150 190046 529218 190102
rect 529274 190046 529342 190102
rect 529398 190046 546970 190102
rect 547026 190046 547094 190102
rect 547150 190046 547218 190102
rect 547274 190046 547342 190102
rect 547398 190046 564970 190102
rect 565026 190046 565094 190102
rect 565150 190046 565218 190102
rect 565274 190046 565342 190102
rect 565398 190046 582970 190102
rect 583026 190046 583094 190102
rect 583150 190046 583218 190102
rect 583274 190046 583342 190102
rect 583398 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 6970 189978
rect 7026 189922 7094 189978
rect 7150 189922 7218 189978
rect 7274 189922 7342 189978
rect 7398 189922 24970 189978
rect 25026 189922 25094 189978
rect 25150 189922 25218 189978
rect 25274 189922 25342 189978
rect 25398 189922 42970 189978
rect 43026 189922 43094 189978
rect 43150 189922 43218 189978
rect 43274 189922 43342 189978
rect 43398 189922 60970 189978
rect 61026 189922 61094 189978
rect 61150 189922 61218 189978
rect 61274 189922 61342 189978
rect 61398 189922 78970 189978
rect 79026 189922 79094 189978
rect 79150 189922 79218 189978
rect 79274 189922 79342 189978
rect 79398 189922 96970 189978
rect 97026 189922 97094 189978
rect 97150 189922 97218 189978
rect 97274 189922 97342 189978
rect 97398 189922 114970 189978
rect 115026 189922 115094 189978
rect 115150 189922 115218 189978
rect 115274 189922 115342 189978
rect 115398 189922 132970 189978
rect 133026 189922 133094 189978
rect 133150 189922 133218 189978
rect 133274 189922 133342 189978
rect 133398 189922 150970 189978
rect 151026 189922 151094 189978
rect 151150 189922 151218 189978
rect 151274 189922 151342 189978
rect 151398 189922 168970 189978
rect 169026 189922 169094 189978
rect 169150 189922 169218 189978
rect 169274 189922 169342 189978
rect 169398 189922 186970 189978
rect 187026 189922 187094 189978
rect 187150 189922 187218 189978
rect 187274 189922 187342 189978
rect 187398 189922 204970 189978
rect 205026 189922 205094 189978
rect 205150 189922 205218 189978
rect 205274 189922 205342 189978
rect 205398 189922 222970 189978
rect 223026 189922 223094 189978
rect 223150 189922 223218 189978
rect 223274 189922 223342 189978
rect 223398 189922 240970 189978
rect 241026 189922 241094 189978
rect 241150 189922 241218 189978
rect 241274 189922 241342 189978
rect 241398 189922 258970 189978
rect 259026 189922 259094 189978
rect 259150 189922 259218 189978
rect 259274 189922 259342 189978
rect 259398 189922 276970 189978
rect 277026 189922 277094 189978
rect 277150 189922 277218 189978
rect 277274 189922 277342 189978
rect 277398 189922 294970 189978
rect 295026 189922 295094 189978
rect 295150 189922 295218 189978
rect 295274 189922 295342 189978
rect 295398 189922 312970 189978
rect 313026 189922 313094 189978
rect 313150 189922 313218 189978
rect 313274 189922 313342 189978
rect 313398 189922 330970 189978
rect 331026 189922 331094 189978
rect 331150 189922 331218 189978
rect 331274 189922 331342 189978
rect 331398 189922 348970 189978
rect 349026 189922 349094 189978
rect 349150 189922 349218 189978
rect 349274 189922 349342 189978
rect 349398 189922 366970 189978
rect 367026 189922 367094 189978
rect 367150 189922 367218 189978
rect 367274 189922 367342 189978
rect 367398 189922 384970 189978
rect 385026 189922 385094 189978
rect 385150 189922 385218 189978
rect 385274 189922 385342 189978
rect 385398 189922 402970 189978
rect 403026 189922 403094 189978
rect 403150 189922 403218 189978
rect 403274 189922 403342 189978
rect 403398 189922 420970 189978
rect 421026 189922 421094 189978
rect 421150 189922 421218 189978
rect 421274 189922 421342 189978
rect 421398 189922 438970 189978
rect 439026 189922 439094 189978
rect 439150 189922 439218 189978
rect 439274 189922 439342 189978
rect 439398 189922 456970 189978
rect 457026 189922 457094 189978
rect 457150 189922 457218 189978
rect 457274 189922 457342 189978
rect 457398 189922 474970 189978
rect 475026 189922 475094 189978
rect 475150 189922 475218 189978
rect 475274 189922 475342 189978
rect 475398 189922 492970 189978
rect 493026 189922 493094 189978
rect 493150 189922 493218 189978
rect 493274 189922 493342 189978
rect 493398 189922 510970 189978
rect 511026 189922 511094 189978
rect 511150 189922 511218 189978
rect 511274 189922 511342 189978
rect 511398 189922 528970 189978
rect 529026 189922 529094 189978
rect 529150 189922 529218 189978
rect 529274 189922 529342 189978
rect 529398 189922 546970 189978
rect 547026 189922 547094 189978
rect 547150 189922 547218 189978
rect 547274 189922 547342 189978
rect 547398 189922 564970 189978
rect 565026 189922 565094 189978
rect 565150 189922 565218 189978
rect 565274 189922 565342 189978
rect 565398 189922 582970 189978
rect 583026 189922 583094 189978
rect 583150 189922 583218 189978
rect 583274 189922 583342 189978
rect 583398 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 3250 184350
rect 3306 184294 3374 184350
rect 3430 184294 3498 184350
rect 3554 184294 3622 184350
rect 3678 184294 21250 184350
rect 21306 184294 21374 184350
rect 21430 184294 21498 184350
rect 21554 184294 21622 184350
rect 21678 184294 39250 184350
rect 39306 184294 39374 184350
rect 39430 184294 39498 184350
rect 39554 184294 39622 184350
rect 39678 184294 57250 184350
rect 57306 184294 57374 184350
rect 57430 184294 57498 184350
rect 57554 184294 57622 184350
rect 57678 184294 75250 184350
rect 75306 184294 75374 184350
rect 75430 184294 75498 184350
rect 75554 184294 75622 184350
rect 75678 184294 93250 184350
rect 93306 184294 93374 184350
rect 93430 184294 93498 184350
rect 93554 184294 93622 184350
rect 93678 184294 111250 184350
rect 111306 184294 111374 184350
rect 111430 184294 111498 184350
rect 111554 184294 111622 184350
rect 111678 184294 129250 184350
rect 129306 184294 129374 184350
rect 129430 184294 129498 184350
rect 129554 184294 129622 184350
rect 129678 184294 147250 184350
rect 147306 184294 147374 184350
rect 147430 184294 147498 184350
rect 147554 184294 147622 184350
rect 147678 184294 165250 184350
rect 165306 184294 165374 184350
rect 165430 184294 165498 184350
rect 165554 184294 165622 184350
rect 165678 184294 183250 184350
rect 183306 184294 183374 184350
rect 183430 184294 183498 184350
rect 183554 184294 183622 184350
rect 183678 184294 201250 184350
rect 201306 184294 201374 184350
rect 201430 184294 201498 184350
rect 201554 184294 201622 184350
rect 201678 184294 219250 184350
rect 219306 184294 219374 184350
rect 219430 184294 219498 184350
rect 219554 184294 219622 184350
rect 219678 184294 237250 184350
rect 237306 184294 237374 184350
rect 237430 184294 237498 184350
rect 237554 184294 237622 184350
rect 237678 184294 255250 184350
rect 255306 184294 255374 184350
rect 255430 184294 255498 184350
rect 255554 184294 255622 184350
rect 255678 184294 273250 184350
rect 273306 184294 273374 184350
rect 273430 184294 273498 184350
rect 273554 184294 273622 184350
rect 273678 184294 291250 184350
rect 291306 184294 291374 184350
rect 291430 184294 291498 184350
rect 291554 184294 291622 184350
rect 291678 184294 309250 184350
rect 309306 184294 309374 184350
rect 309430 184294 309498 184350
rect 309554 184294 309622 184350
rect 309678 184294 327250 184350
rect 327306 184294 327374 184350
rect 327430 184294 327498 184350
rect 327554 184294 327622 184350
rect 327678 184294 345250 184350
rect 345306 184294 345374 184350
rect 345430 184294 345498 184350
rect 345554 184294 345622 184350
rect 345678 184294 363250 184350
rect 363306 184294 363374 184350
rect 363430 184294 363498 184350
rect 363554 184294 363622 184350
rect 363678 184294 381250 184350
rect 381306 184294 381374 184350
rect 381430 184294 381498 184350
rect 381554 184294 381622 184350
rect 381678 184294 399250 184350
rect 399306 184294 399374 184350
rect 399430 184294 399498 184350
rect 399554 184294 399622 184350
rect 399678 184294 417250 184350
rect 417306 184294 417374 184350
rect 417430 184294 417498 184350
rect 417554 184294 417622 184350
rect 417678 184294 435250 184350
rect 435306 184294 435374 184350
rect 435430 184294 435498 184350
rect 435554 184294 435622 184350
rect 435678 184294 453250 184350
rect 453306 184294 453374 184350
rect 453430 184294 453498 184350
rect 453554 184294 453622 184350
rect 453678 184294 471250 184350
rect 471306 184294 471374 184350
rect 471430 184294 471498 184350
rect 471554 184294 471622 184350
rect 471678 184294 489250 184350
rect 489306 184294 489374 184350
rect 489430 184294 489498 184350
rect 489554 184294 489622 184350
rect 489678 184294 507250 184350
rect 507306 184294 507374 184350
rect 507430 184294 507498 184350
rect 507554 184294 507622 184350
rect 507678 184294 525250 184350
rect 525306 184294 525374 184350
rect 525430 184294 525498 184350
rect 525554 184294 525622 184350
rect 525678 184294 543250 184350
rect 543306 184294 543374 184350
rect 543430 184294 543498 184350
rect 543554 184294 543622 184350
rect 543678 184294 561250 184350
rect 561306 184294 561374 184350
rect 561430 184294 561498 184350
rect 561554 184294 561622 184350
rect 561678 184294 579250 184350
rect 579306 184294 579374 184350
rect 579430 184294 579498 184350
rect 579554 184294 579622 184350
rect 579678 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 3250 184226
rect 3306 184170 3374 184226
rect 3430 184170 3498 184226
rect 3554 184170 3622 184226
rect 3678 184170 21250 184226
rect 21306 184170 21374 184226
rect 21430 184170 21498 184226
rect 21554 184170 21622 184226
rect 21678 184170 39250 184226
rect 39306 184170 39374 184226
rect 39430 184170 39498 184226
rect 39554 184170 39622 184226
rect 39678 184170 57250 184226
rect 57306 184170 57374 184226
rect 57430 184170 57498 184226
rect 57554 184170 57622 184226
rect 57678 184170 75250 184226
rect 75306 184170 75374 184226
rect 75430 184170 75498 184226
rect 75554 184170 75622 184226
rect 75678 184170 93250 184226
rect 93306 184170 93374 184226
rect 93430 184170 93498 184226
rect 93554 184170 93622 184226
rect 93678 184170 111250 184226
rect 111306 184170 111374 184226
rect 111430 184170 111498 184226
rect 111554 184170 111622 184226
rect 111678 184170 129250 184226
rect 129306 184170 129374 184226
rect 129430 184170 129498 184226
rect 129554 184170 129622 184226
rect 129678 184170 147250 184226
rect 147306 184170 147374 184226
rect 147430 184170 147498 184226
rect 147554 184170 147622 184226
rect 147678 184170 165250 184226
rect 165306 184170 165374 184226
rect 165430 184170 165498 184226
rect 165554 184170 165622 184226
rect 165678 184170 183250 184226
rect 183306 184170 183374 184226
rect 183430 184170 183498 184226
rect 183554 184170 183622 184226
rect 183678 184170 201250 184226
rect 201306 184170 201374 184226
rect 201430 184170 201498 184226
rect 201554 184170 201622 184226
rect 201678 184170 219250 184226
rect 219306 184170 219374 184226
rect 219430 184170 219498 184226
rect 219554 184170 219622 184226
rect 219678 184170 237250 184226
rect 237306 184170 237374 184226
rect 237430 184170 237498 184226
rect 237554 184170 237622 184226
rect 237678 184170 255250 184226
rect 255306 184170 255374 184226
rect 255430 184170 255498 184226
rect 255554 184170 255622 184226
rect 255678 184170 273250 184226
rect 273306 184170 273374 184226
rect 273430 184170 273498 184226
rect 273554 184170 273622 184226
rect 273678 184170 291250 184226
rect 291306 184170 291374 184226
rect 291430 184170 291498 184226
rect 291554 184170 291622 184226
rect 291678 184170 309250 184226
rect 309306 184170 309374 184226
rect 309430 184170 309498 184226
rect 309554 184170 309622 184226
rect 309678 184170 327250 184226
rect 327306 184170 327374 184226
rect 327430 184170 327498 184226
rect 327554 184170 327622 184226
rect 327678 184170 345250 184226
rect 345306 184170 345374 184226
rect 345430 184170 345498 184226
rect 345554 184170 345622 184226
rect 345678 184170 363250 184226
rect 363306 184170 363374 184226
rect 363430 184170 363498 184226
rect 363554 184170 363622 184226
rect 363678 184170 381250 184226
rect 381306 184170 381374 184226
rect 381430 184170 381498 184226
rect 381554 184170 381622 184226
rect 381678 184170 399250 184226
rect 399306 184170 399374 184226
rect 399430 184170 399498 184226
rect 399554 184170 399622 184226
rect 399678 184170 417250 184226
rect 417306 184170 417374 184226
rect 417430 184170 417498 184226
rect 417554 184170 417622 184226
rect 417678 184170 435250 184226
rect 435306 184170 435374 184226
rect 435430 184170 435498 184226
rect 435554 184170 435622 184226
rect 435678 184170 453250 184226
rect 453306 184170 453374 184226
rect 453430 184170 453498 184226
rect 453554 184170 453622 184226
rect 453678 184170 471250 184226
rect 471306 184170 471374 184226
rect 471430 184170 471498 184226
rect 471554 184170 471622 184226
rect 471678 184170 489250 184226
rect 489306 184170 489374 184226
rect 489430 184170 489498 184226
rect 489554 184170 489622 184226
rect 489678 184170 507250 184226
rect 507306 184170 507374 184226
rect 507430 184170 507498 184226
rect 507554 184170 507622 184226
rect 507678 184170 525250 184226
rect 525306 184170 525374 184226
rect 525430 184170 525498 184226
rect 525554 184170 525622 184226
rect 525678 184170 543250 184226
rect 543306 184170 543374 184226
rect 543430 184170 543498 184226
rect 543554 184170 543622 184226
rect 543678 184170 561250 184226
rect 561306 184170 561374 184226
rect 561430 184170 561498 184226
rect 561554 184170 561622 184226
rect 561678 184170 579250 184226
rect 579306 184170 579374 184226
rect 579430 184170 579498 184226
rect 579554 184170 579622 184226
rect 579678 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 3250 184102
rect 3306 184046 3374 184102
rect 3430 184046 3498 184102
rect 3554 184046 3622 184102
rect 3678 184046 21250 184102
rect 21306 184046 21374 184102
rect 21430 184046 21498 184102
rect 21554 184046 21622 184102
rect 21678 184046 39250 184102
rect 39306 184046 39374 184102
rect 39430 184046 39498 184102
rect 39554 184046 39622 184102
rect 39678 184046 57250 184102
rect 57306 184046 57374 184102
rect 57430 184046 57498 184102
rect 57554 184046 57622 184102
rect 57678 184046 75250 184102
rect 75306 184046 75374 184102
rect 75430 184046 75498 184102
rect 75554 184046 75622 184102
rect 75678 184046 93250 184102
rect 93306 184046 93374 184102
rect 93430 184046 93498 184102
rect 93554 184046 93622 184102
rect 93678 184046 111250 184102
rect 111306 184046 111374 184102
rect 111430 184046 111498 184102
rect 111554 184046 111622 184102
rect 111678 184046 129250 184102
rect 129306 184046 129374 184102
rect 129430 184046 129498 184102
rect 129554 184046 129622 184102
rect 129678 184046 147250 184102
rect 147306 184046 147374 184102
rect 147430 184046 147498 184102
rect 147554 184046 147622 184102
rect 147678 184046 165250 184102
rect 165306 184046 165374 184102
rect 165430 184046 165498 184102
rect 165554 184046 165622 184102
rect 165678 184046 183250 184102
rect 183306 184046 183374 184102
rect 183430 184046 183498 184102
rect 183554 184046 183622 184102
rect 183678 184046 201250 184102
rect 201306 184046 201374 184102
rect 201430 184046 201498 184102
rect 201554 184046 201622 184102
rect 201678 184046 219250 184102
rect 219306 184046 219374 184102
rect 219430 184046 219498 184102
rect 219554 184046 219622 184102
rect 219678 184046 237250 184102
rect 237306 184046 237374 184102
rect 237430 184046 237498 184102
rect 237554 184046 237622 184102
rect 237678 184046 255250 184102
rect 255306 184046 255374 184102
rect 255430 184046 255498 184102
rect 255554 184046 255622 184102
rect 255678 184046 273250 184102
rect 273306 184046 273374 184102
rect 273430 184046 273498 184102
rect 273554 184046 273622 184102
rect 273678 184046 291250 184102
rect 291306 184046 291374 184102
rect 291430 184046 291498 184102
rect 291554 184046 291622 184102
rect 291678 184046 309250 184102
rect 309306 184046 309374 184102
rect 309430 184046 309498 184102
rect 309554 184046 309622 184102
rect 309678 184046 327250 184102
rect 327306 184046 327374 184102
rect 327430 184046 327498 184102
rect 327554 184046 327622 184102
rect 327678 184046 345250 184102
rect 345306 184046 345374 184102
rect 345430 184046 345498 184102
rect 345554 184046 345622 184102
rect 345678 184046 363250 184102
rect 363306 184046 363374 184102
rect 363430 184046 363498 184102
rect 363554 184046 363622 184102
rect 363678 184046 381250 184102
rect 381306 184046 381374 184102
rect 381430 184046 381498 184102
rect 381554 184046 381622 184102
rect 381678 184046 399250 184102
rect 399306 184046 399374 184102
rect 399430 184046 399498 184102
rect 399554 184046 399622 184102
rect 399678 184046 417250 184102
rect 417306 184046 417374 184102
rect 417430 184046 417498 184102
rect 417554 184046 417622 184102
rect 417678 184046 435250 184102
rect 435306 184046 435374 184102
rect 435430 184046 435498 184102
rect 435554 184046 435622 184102
rect 435678 184046 453250 184102
rect 453306 184046 453374 184102
rect 453430 184046 453498 184102
rect 453554 184046 453622 184102
rect 453678 184046 471250 184102
rect 471306 184046 471374 184102
rect 471430 184046 471498 184102
rect 471554 184046 471622 184102
rect 471678 184046 489250 184102
rect 489306 184046 489374 184102
rect 489430 184046 489498 184102
rect 489554 184046 489622 184102
rect 489678 184046 507250 184102
rect 507306 184046 507374 184102
rect 507430 184046 507498 184102
rect 507554 184046 507622 184102
rect 507678 184046 525250 184102
rect 525306 184046 525374 184102
rect 525430 184046 525498 184102
rect 525554 184046 525622 184102
rect 525678 184046 543250 184102
rect 543306 184046 543374 184102
rect 543430 184046 543498 184102
rect 543554 184046 543622 184102
rect 543678 184046 561250 184102
rect 561306 184046 561374 184102
rect 561430 184046 561498 184102
rect 561554 184046 561622 184102
rect 561678 184046 579250 184102
rect 579306 184046 579374 184102
rect 579430 184046 579498 184102
rect 579554 184046 579622 184102
rect 579678 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 3250 183978
rect 3306 183922 3374 183978
rect 3430 183922 3498 183978
rect 3554 183922 3622 183978
rect 3678 183922 21250 183978
rect 21306 183922 21374 183978
rect 21430 183922 21498 183978
rect 21554 183922 21622 183978
rect 21678 183922 39250 183978
rect 39306 183922 39374 183978
rect 39430 183922 39498 183978
rect 39554 183922 39622 183978
rect 39678 183922 57250 183978
rect 57306 183922 57374 183978
rect 57430 183922 57498 183978
rect 57554 183922 57622 183978
rect 57678 183922 75250 183978
rect 75306 183922 75374 183978
rect 75430 183922 75498 183978
rect 75554 183922 75622 183978
rect 75678 183922 93250 183978
rect 93306 183922 93374 183978
rect 93430 183922 93498 183978
rect 93554 183922 93622 183978
rect 93678 183922 111250 183978
rect 111306 183922 111374 183978
rect 111430 183922 111498 183978
rect 111554 183922 111622 183978
rect 111678 183922 129250 183978
rect 129306 183922 129374 183978
rect 129430 183922 129498 183978
rect 129554 183922 129622 183978
rect 129678 183922 147250 183978
rect 147306 183922 147374 183978
rect 147430 183922 147498 183978
rect 147554 183922 147622 183978
rect 147678 183922 165250 183978
rect 165306 183922 165374 183978
rect 165430 183922 165498 183978
rect 165554 183922 165622 183978
rect 165678 183922 183250 183978
rect 183306 183922 183374 183978
rect 183430 183922 183498 183978
rect 183554 183922 183622 183978
rect 183678 183922 201250 183978
rect 201306 183922 201374 183978
rect 201430 183922 201498 183978
rect 201554 183922 201622 183978
rect 201678 183922 219250 183978
rect 219306 183922 219374 183978
rect 219430 183922 219498 183978
rect 219554 183922 219622 183978
rect 219678 183922 237250 183978
rect 237306 183922 237374 183978
rect 237430 183922 237498 183978
rect 237554 183922 237622 183978
rect 237678 183922 255250 183978
rect 255306 183922 255374 183978
rect 255430 183922 255498 183978
rect 255554 183922 255622 183978
rect 255678 183922 273250 183978
rect 273306 183922 273374 183978
rect 273430 183922 273498 183978
rect 273554 183922 273622 183978
rect 273678 183922 291250 183978
rect 291306 183922 291374 183978
rect 291430 183922 291498 183978
rect 291554 183922 291622 183978
rect 291678 183922 309250 183978
rect 309306 183922 309374 183978
rect 309430 183922 309498 183978
rect 309554 183922 309622 183978
rect 309678 183922 327250 183978
rect 327306 183922 327374 183978
rect 327430 183922 327498 183978
rect 327554 183922 327622 183978
rect 327678 183922 345250 183978
rect 345306 183922 345374 183978
rect 345430 183922 345498 183978
rect 345554 183922 345622 183978
rect 345678 183922 363250 183978
rect 363306 183922 363374 183978
rect 363430 183922 363498 183978
rect 363554 183922 363622 183978
rect 363678 183922 381250 183978
rect 381306 183922 381374 183978
rect 381430 183922 381498 183978
rect 381554 183922 381622 183978
rect 381678 183922 399250 183978
rect 399306 183922 399374 183978
rect 399430 183922 399498 183978
rect 399554 183922 399622 183978
rect 399678 183922 417250 183978
rect 417306 183922 417374 183978
rect 417430 183922 417498 183978
rect 417554 183922 417622 183978
rect 417678 183922 435250 183978
rect 435306 183922 435374 183978
rect 435430 183922 435498 183978
rect 435554 183922 435622 183978
rect 435678 183922 453250 183978
rect 453306 183922 453374 183978
rect 453430 183922 453498 183978
rect 453554 183922 453622 183978
rect 453678 183922 471250 183978
rect 471306 183922 471374 183978
rect 471430 183922 471498 183978
rect 471554 183922 471622 183978
rect 471678 183922 489250 183978
rect 489306 183922 489374 183978
rect 489430 183922 489498 183978
rect 489554 183922 489622 183978
rect 489678 183922 507250 183978
rect 507306 183922 507374 183978
rect 507430 183922 507498 183978
rect 507554 183922 507622 183978
rect 507678 183922 525250 183978
rect 525306 183922 525374 183978
rect 525430 183922 525498 183978
rect 525554 183922 525622 183978
rect 525678 183922 543250 183978
rect 543306 183922 543374 183978
rect 543430 183922 543498 183978
rect 543554 183922 543622 183978
rect 543678 183922 561250 183978
rect 561306 183922 561374 183978
rect 561430 183922 561498 183978
rect 561554 183922 561622 183978
rect 561678 183922 579250 183978
rect 579306 183922 579374 183978
rect 579430 183922 579498 183978
rect 579554 183922 579622 183978
rect 579678 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 6970 172350
rect 7026 172294 7094 172350
rect 7150 172294 7218 172350
rect 7274 172294 7342 172350
rect 7398 172294 24970 172350
rect 25026 172294 25094 172350
rect 25150 172294 25218 172350
rect 25274 172294 25342 172350
rect 25398 172294 42970 172350
rect 43026 172294 43094 172350
rect 43150 172294 43218 172350
rect 43274 172294 43342 172350
rect 43398 172294 60970 172350
rect 61026 172294 61094 172350
rect 61150 172294 61218 172350
rect 61274 172294 61342 172350
rect 61398 172294 78970 172350
rect 79026 172294 79094 172350
rect 79150 172294 79218 172350
rect 79274 172294 79342 172350
rect 79398 172294 96970 172350
rect 97026 172294 97094 172350
rect 97150 172294 97218 172350
rect 97274 172294 97342 172350
rect 97398 172294 114970 172350
rect 115026 172294 115094 172350
rect 115150 172294 115218 172350
rect 115274 172294 115342 172350
rect 115398 172294 132970 172350
rect 133026 172294 133094 172350
rect 133150 172294 133218 172350
rect 133274 172294 133342 172350
rect 133398 172294 150970 172350
rect 151026 172294 151094 172350
rect 151150 172294 151218 172350
rect 151274 172294 151342 172350
rect 151398 172294 168970 172350
rect 169026 172294 169094 172350
rect 169150 172294 169218 172350
rect 169274 172294 169342 172350
rect 169398 172294 186970 172350
rect 187026 172294 187094 172350
rect 187150 172294 187218 172350
rect 187274 172294 187342 172350
rect 187398 172294 204970 172350
rect 205026 172294 205094 172350
rect 205150 172294 205218 172350
rect 205274 172294 205342 172350
rect 205398 172294 222970 172350
rect 223026 172294 223094 172350
rect 223150 172294 223218 172350
rect 223274 172294 223342 172350
rect 223398 172294 240970 172350
rect 241026 172294 241094 172350
rect 241150 172294 241218 172350
rect 241274 172294 241342 172350
rect 241398 172294 258970 172350
rect 259026 172294 259094 172350
rect 259150 172294 259218 172350
rect 259274 172294 259342 172350
rect 259398 172294 276970 172350
rect 277026 172294 277094 172350
rect 277150 172294 277218 172350
rect 277274 172294 277342 172350
rect 277398 172294 294970 172350
rect 295026 172294 295094 172350
rect 295150 172294 295218 172350
rect 295274 172294 295342 172350
rect 295398 172294 312970 172350
rect 313026 172294 313094 172350
rect 313150 172294 313218 172350
rect 313274 172294 313342 172350
rect 313398 172294 330970 172350
rect 331026 172294 331094 172350
rect 331150 172294 331218 172350
rect 331274 172294 331342 172350
rect 331398 172294 348970 172350
rect 349026 172294 349094 172350
rect 349150 172294 349218 172350
rect 349274 172294 349342 172350
rect 349398 172294 366970 172350
rect 367026 172294 367094 172350
rect 367150 172294 367218 172350
rect 367274 172294 367342 172350
rect 367398 172294 384970 172350
rect 385026 172294 385094 172350
rect 385150 172294 385218 172350
rect 385274 172294 385342 172350
rect 385398 172294 402970 172350
rect 403026 172294 403094 172350
rect 403150 172294 403218 172350
rect 403274 172294 403342 172350
rect 403398 172294 420970 172350
rect 421026 172294 421094 172350
rect 421150 172294 421218 172350
rect 421274 172294 421342 172350
rect 421398 172294 438970 172350
rect 439026 172294 439094 172350
rect 439150 172294 439218 172350
rect 439274 172294 439342 172350
rect 439398 172294 456970 172350
rect 457026 172294 457094 172350
rect 457150 172294 457218 172350
rect 457274 172294 457342 172350
rect 457398 172294 474970 172350
rect 475026 172294 475094 172350
rect 475150 172294 475218 172350
rect 475274 172294 475342 172350
rect 475398 172294 492970 172350
rect 493026 172294 493094 172350
rect 493150 172294 493218 172350
rect 493274 172294 493342 172350
rect 493398 172294 510970 172350
rect 511026 172294 511094 172350
rect 511150 172294 511218 172350
rect 511274 172294 511342 172350
rect 511398 172294 528970 172350
rect 529026 172294 529094 172350
rect 529150 172294 529218 172350
rect 529274 172294 529342 172350
rect 529398 172294 546970 172350
rect 547026 172294 547094 172350
rect 547150 172294 547218 172350
rect 547274 172294 547342 172350
rect 547398 172294 564970 172350
rect 565026 172294 565094 172350
rect 565150 172294 565218 172350
rect 565274 172294 565342 172350
rect 565398 172294 582970 172350
rect 583026 172294 583094 172350
rect 583150 172294 583218 172350
rect 583274 172294 583342 172350
rect 583398 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 6970 172226
rect 7026 172170 7094 172226
rect 7150 172170 7218 172226
rect 7274 172170 7342 172226
rect 7398 172170 24970 172226
rect 25026 172170 25094 172226
rect 25150 172170 25218 172226
rect 25274 172170 25342 172226
rect 25398 172170 42970 172226
rect 43026 172170 43094 172226
rect 43150 172170 43218 172226
rect 43274 172170 43342 172226
rect 43398 172170 60970 172226
rect 61026 172170 61094 172226
rect 61150 172170 61218 172226
rect 61274 172170 61342 172226
rect 61398 172170 78970 172226
rect 79026 172170 79094 172226
rect 79150 172170 79218 172226
rect 79274 172170 79342 172226
rect 79398 172170 96970 172226
rect 97026 172170 97094 172226
rect 97150 172170 97218 172226
rect 97274 172170 97342 172226
rect 97398 172170 114970 172226
rect 115026 172170 115094 172226
rect 115150 172170 115218 172226
rect 115274 172170 115342 172226
rect 115398 172170 132970 172226
rect 133026 172170 133094 172226
rect 133150 172170 133218 172226
rect 133274 172170 133342 172226
rect 133398 172170 150970 172226
rect 151026 172170 151094 172226
rect 151150 172170 151218 172226
rect 151274 172170 151342 172226
rect 151398 172170 168970 172226
rect 169026 172170 169094 172226
rect 169150 172170 169218 172226
rect 169274 172170 169342 172226
rect 169398 172170 186970 172226
rect 187026 172170 187094 172226
rect 187150 172170 187218 172226
rect 187274 172170 187342 172226
rect 187398 172170 204970 172226
rect 205026 172170 205094 172226
rect 205150 172170 205218 172226
rect 205274 172170 205342 172226
rect 205398 172170 222970 172226
rect 223026 172170 223094 172226
rect 223150 172170 223218 172226
rect 223274 172170 223342 172226
rect 223398 172170 240970 172226
rect 241026 172170 241094 172226
rect 241150 172170 241218 172226
rect 241274 172170 241342 172226
rect 241398 172170 258970 172226
rect 259026 172170 259094 172226
rect 259150 172170 259218 172226
rect 259274 172170 259342 172226
rect 259398 172170 276970 172226
rect 277026 172170 277094 172226
rect 277150 172170 277218 172226
rect 277274 172170 277342 172226
rect 277398 172170 294970 172226
rect 295026 172170 295094 172226
rect 295150 172170 295218 172226
rect 295274 172170 295342 172226
rect 295398 172170 312970 172226
rect 313026 172170 313094 172226
rect 313150 172170 313218 172226
rect 313274 172170 313342 172226
rect 313398 172170 330970 172226
rect 331026 172170 331094 172226
rect 331150 172170 331218 172226
rect 331274 172170 331342 172226
rect 331398 172170 348970 172226
rect 349026 172170 349094 172226
rect 349150 172170 349218 172226
rect 349274 172170 349342 172226
rect 349398 172170 366970 172226
rect 367026 172170 367094 172226
rect 367150 172170 367218 172226
rect 367274 172170 367342 172226
rect 367398 172170 384970 172226
rect 385026 172170 385094 172226
rect 385150 172170 385218 172226
rect 385274 172170 385342 172226
rect 385398 172170 402970 172226
rect 403026 172170 403094 172226
rect 403150 172170 403218 172226
rect 403274 172170 403342 172226
rect 403398 172170 420970 172226
rect 421026 172170 421094 172226
rect 421150 172170 421218 172226
rect 421274 172170 421342 172226
rect 421398 172170 438970 172226
rect 439026 172170 439094 172226
rect 439150 172170 439218 172226
rect 439274 172170 439342 172226
rect 439398 172170 456970 172226
rect 457026 172170 457094 172226
rect 457150 172170 457218 172226
rect 457274 172170 457342 172226
rect 457398 172170 474970 172226
rect 475026 172170 475094 172226
rect 475150 172170 475218 172226
rect 475274 172170 475342 172226
rect 475398 172170 492970 172226
rect 493026 172170 493094 172226
rect 493150 172170 493218 172226
rect 493274 172170 493342 172226
rect 493398 172170 510970 172226
rect 511026 172170 511094 172226
rect 511150 172170 511218 172226
rect 511274 172170 511342 172226
rect 511398 172170 528970 172226
rect 529026 172170 529094 172226
rect 529150 172170 529218 172226
rect 529274 172170 529342 172226
rect 529398 172170 546970 172226
rect 547026 172170 547094 172226
rect 547150 172170 547218 172226
rect 547274 172170 547342 172226
rect 547398 172170 564970 172226
rect 565026 172170 565094 172226
rect 565150 172170 565218 172226
rect 565274 172170 565342 172226
rect 565398 172170 582970 172226
rect 583026 172170 583094 172226
rect 583150 172170 583218 172226
rect 583274 172170 583342 172226
rect 583398 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 6970 172102
rect 7026 172046 7094 172102
rect 7150 172046 7218 172102
rect 7274 172046 7342 172102
rect 7398 172046 24970 172102
rect 25026 172046 25094 172102
rect 25150 172046 25218 172102
rect 25274 172046 25342 172102
rect 25398 172046 42970 172102
rect 43026 172046 43094 172102
rect 43150 172046 43218 172102
rect 43274 172046 43342 172102
rect 43398 172046 60970 172102
rect 61026 172046 61094 172102
rect 61150 172046 61218 172102
rect 61274 172046 61342 172102
rect 61398 172046 78970 172102
rect 79026 172046 79094 172102
rect 79150 172046 79218 172102
rect 79274 172046 79342 172102
rect 79398 172046 96970 172102
rect 97026 172046 97094 172102
rect 97150 172046 97218 172102
rect 97274 172046 97342 172102
rect 97398 172046 114970 172102
rect 115026 172046 115094 172102
rect 115150 172046 115218 172102
rect 115274 172046 115342 172102
rect 115398 172046 132970 172102
rect 133026 172046 133094 172102
rect 133150 172046 133218 172102
rect 133274 172046 133342 172102
rect 133398 172046 150970 172102
rect 151026 172046 151094 172102
rect 151150 172046 151218 172102
rect 151274 172046 151342 172102
rect 151398 172046 168970 172102
rect 169026 172046 169094 172102
rect 169150 172046 169218 172102
rect 169274 172046 169342 172102
rect 169398 172046 186970 172102
rect 187026 172046 187094 172102
rect 187150 172046 187218 172102
rect 187274 172046 187342 172102
rect 187398 172046 204970 172102
rect 205026 172046 205094 172102
rect 205150 172046 205218 172102
rect 205274 172046 205342 172102
rect 205398 172046 222970 172102
rect 223026 172046 223094 172102
rect 223150 172046 223218 172102
rect 223274 172046 223342 172102
rect 223398 172046 240970 172102
rect 241026 172046 241094 172102
rect 241150 172046 241218 172102
rect 241274 172046 241342 172102
rect 241398 172046 258970 172102
rect 259026 172046 259094 172102
rect 259150 172046 259218 172102
rect 259274 172046 259342 172102
rect 259398 172046 276970 172102
rect 277026 172046 277094 172102
rect 277150 172046 277218 172102
rect 277274 172046 277342 172102
rect 277398 172046 294970 172102
rect 295026 172046 295094 172102
rect 295150 172046 295218 172102
rect 295274 172046 295342 172102
rect 295398 172046 312970 172102
rect 313026 172046 313094 172102
rect 313150 172046 313218 172102
rect 313274 172046 313342 172102
rect 313398 172046 330970 172102
rect 331026 172046 331094 172102
rect 331150 172046 331218 172102
rect 331274 172046 331342 172102
rect 331398 172046 348970 172102
rect 349026 172046 349094 172102
rect 349150 172046 349218 172102
rect 349274 172046 349342 172102
rect 349398 172046 366970 172102
rect 367026 172046 367094 172102
rect 367150 172046 367218 172102
rect 367274 172046 367342 172102
rect 367398 172046 384970 172102
rect 385026 172046 385094 172102
rect 385150 172046 385218 172102
rect 385274 172046 385342 172102
rect 385398 172046 402970 172102
rect 403026 172046 403094 172102
rect 403150 172046 403218 172102
rect 403274 172046 403342 172102
rect 403398 172046 420970 172102
rect 421026 172046 421094 172102
rect 421150 172046 421218 172102
rect 421274 172046 421342 172102
rect 421398 172046 438970 172102
rect 439026 172046 439094 172102
rect 439150 172046 439218 172102
rect 439274 172046 439342 172102
rect 439398 172046 456970 172102
rect 457026 172046 457094 172102
rect 457150 172046 457218 172102
rect 457274 172046 457342 172102
rect 457398 172046 474970 172102
rect 475026 172046 475094 172102
rect 475150 172046 475218 172102
rect 475274 172046 475342 172102
rect 475398 172046 492970 172102
rect 493026 172046 493094 172102
rect 493150 172046 493218 172102
rect 493274 172046 493342 172102
rect 493398 172046 510970 172102
rect 511026 172046 511094 172102
rect 511150 172046 511218 172102
rect 511274 172046 511342 172102
rect 511398 172046 528970 172102
rect 529026 172046 529094 172102
rect 529150 172046 529218 172102
rect 529274 172046 529342 172102
rect 529398 172046 546970 172102
rect 547026 172046 547094 172102
rect 547150 172046 547218 172102
rect 547274 172046 547342 172102
rect 547398 172046 564970 172102
rect 565026 172046 565094 172102
rect 565150 172046 565218 172102
rect 565274 172046 565342 172102
rect 565398 172046 582970 172102
rect 583026 172046 583094 172102
rect 583150 172046 583218 172102
rect 583274 172046 583342 172102
rect 583398 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 6970 171978
rect 7026 171922 7094 171978
rect 7150 171922 7218 171978
rect 7274 171922 7342 171978
rect 7398 171922 24970 171978
rect 25026 171922 25094 171978
rect 25150 171922 25218 171978
rect 25274 171922 25342 171978
rect 25398 171922 42970 171978
rect 43026 171922 43094 171978
rect 43150 171922 43218 171978
rect 43274 171922 43342 171978
rect 43398 171922 60970 171978
rect 61026 171922 61094 171978
rect 61150 171922 61218 171978
rect 61274 171922 61342 171978
rect 61398 171922 78970 171978
rect 79026 171922 79094 171978
rect 79150 171922 79218 171978
rect 79274 171922 79342 171978
rect 79398 171922 96970 171978
rect 97026 171922 97094 171978
rect 97150 171922 97218 171978
rect 97274 171922 97342 171978
rect 97398 171922 114970 171978
rect 115026 171922 115094 171978
rect 115150 171922 115218 171978
rect 115274 171922 115342 171978
rect 115398 171922 132970 171978
rect 133026 171922 133094 171978
rect 133150 171922 133218 171978
rect 133274 171922 133342 171978
rect 133398 171922 150970 171978
rect 151026 171922 151094 171978
rect 151150 171922 151218 171978
rect 151274 171922 151342 171978
rect 151398 171922 168970 171978
rect 169026 171922 169094 171978
rect 169150 171922 169218 171978
rect 169274 171922 169342 171978
rect 169398 171922 186970 171978
rect 187026 171922 187094 171978
rect 187150 171922 187218 171978
rect 187274 171922 187342 171978
rect 187398 171922 204970 171978
rect 205026 171922 205094 171978
rect 205150 171922 205218 171978
rect 205274 171922 205342 171978
rect 205398 171922 222970 171978
rect 223026 171922 223094 171978
rect 223150 171922 223218 171978
rect 223274 171922 223342 171978
rect 223398 171922 240970 171978
rect 241026 171922 241094 171978
rect 241150 171922 241218 171978
rect 241274 171922 241342 171978
rect 241398 171922 258970 171978
rect 259026 171922 259094 171978
rect 259150 171922 259218 171978
rect 259274 171922 259342 171978
rect 259398 171922 276970 171978
rect 277026 171922 277094 171978
rect 277150 171922 277218 171978
rect 277274 171922 277342 171978
rect 277398 171922 294970 171978
rect 295026 171922 295094 171978
rect 295150 171922 295218 171978
rect 295274 171922 295342 171978
rect 295398 171922 312970 171978
rect 313026 171922 313094 171978
rect 313150 171922 313218 171978
rect 313274 171922 313342 171978
rect 313398 171922 330970 171978
rect 331026 171922 331094 171978
rect 331150 171922 331218 171978
rect 331274 171922 331342 171978
rect 331398 171922 348970 171978
rect 349026 171922 349094 171978
rect 349150 171922 349218 171978
rect 349274 171922 349342 171978
rect 349398 171922 366970 171978
rect 367026 171922 367094 171978
rect 367150 171922 367218 171978
rect 367274 171922 367342 171978
rect 367398 171922 384970 171978
rect 385026 171922 385094 171978
rect 385150 171922 385218 171978
rect 385274 171922 385342 171978
rect 385398 171922 402970 171978
rect 403026 171922 403094 171978
rect 403150 171922 403218 171978
rect 403274 171922 403342 171978
rect 403398 171922 420970 171978
rect 421026 171922 421094 171978
rect 421150 171922 421218 171978
rect 421274 171922 421342 171978
rect 421398 171922 438970 171978
rect 439026 171922 439094 171978
rect 439150 171922 439218 171978
rect 439274 171922 439342 171978
rect 439398 171922 456970 171978
rect 457026 171922 457094 171978
rect 457150 171922 457218 171978
rect 457274 171922 457342 171978
rect 457398 171922 474970 171978
rect 475026 171922 475094 171978
rect 475150 171922 475218 171978
rect 475274 171922 475342 171978
rect 475398 171922 492970 171978
rect 493026 171922 493094 171978
rect 493150 171922 493218 171978
rect 493274 171922 493342 171978
rect 493398 171922 510970 171978
rect 511026 171922 511094 171978
rect 511150 171922 511218 171978
rect 511274 171922 511342 171978
rect 511398 171922 528970 171978
rect 529026 171922 529094 171978
rect 529150 171922 529218 171978
rect 529274 171922 529342 171978
rect 529398 171922 546970 171978
rect 547026 171922 547094 171978
rect 547150 171922 547218 171978
rect 547274 171922 547342 171978
rect 547398 171922 564970 171978
rect 565026 171922 565094 171978
rect 565150 171922 565218 171978
rect 565274 171922 565342 171978
rect 565398 171922 582970 171978
rect 583026 171922 583094 171978
rect 583150 171922 583218 171978
rect 583274 171922 583342 171978
rect 583398 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 3250 166350
rect 3306 166294 3374 166350
rect 3430 166294 3498 166350
rect 3554 166294 3622 166350
rect 3678 166294 21250 166350
rect 21306 166294 21374 166350
rect 21430 166294 21498 166350
rect 21554 166294 21622 166350
rect 21678 166294 39250 166350
rect 39306 166294 39374 166350
rect 39430 166294 39498 166350
rect 39554 166294 39622 166350
rect 39678 166294 57250 166350
rect 57306 166294 57374 166350
rect 57430 166294 57498 166350
rect 57554 166294 57622 166350
rect 57678 166294 75250 166350
rect 75306 166294 75374 166350
rect 75430 166294 75498 166350
rect 75554 166294 75622 166350
rect 75678 166294 93250 166350
rect 93306 166294 93374 166350
rect 93430 166294 93498 166350
rect 93554 166294 93622 166350
rect 93678 166294 111250 166350
rect 111306 166294 111374 166350
rect 111430 166294 111498 166350
rect 111554 166294 111622 166350
rect 111678 166294 129250 166350
rect 129306 166294 129374 166350
rect 129430 166294 129498 166350
rect 129554 166294 129622 166350
rect 129678 166294 147250 166350
rect 147306 166294 147374 166350
rect 147430 166294 147498 166350
rect 147554 166294 147622 166350
rect 147678 166294 165250 166350
rect 165306 166294 165374 166350
rect 165430 166294 165498 166350
rect 165554 166294 165622 166350
rect 165678 166294 183250 166350
rect 183306 166294 183374 166350
rect 183430 166294 183498 166350
rect 183554 166294 183622 166350
rect 183678 166294 201250 166350
rect 201306 166294 201374 166350
rect 201430 166294 201498 166350
rect 201554 166294 201622 166350
rect 201678 166294 219250 166350
rect 219306 166294 219374 166350
rect 219430 166294 219498 166350
rect 219554 166294 219622 166350
rect 219678 166294 237250 166350
rect 237306 166294 237374 166350
rect 237430 166294 237498 166350
rect 237554 166294 237622 166350
rect 237678 166294 255250 166350
rect 255306 166294 255374 166350
rect 255430 166294 255498 166350
rect 255554 166294 255622 166350
rect 255678 166294 273250 166350
rect 273306 166294 273374 166350
rect 273430 166294 273498 166350
rect 273554 166294 273622 166350
rect 273678 166294 291250 166350
rect 291306 166294 291374 166350
rect 291430 166294 291498 166350
rect 291554 166294 291622 166350
rect 291678 166294 309250 166350
rect 309306 166294 309374 166350
rect 309430 166294 309498 166350
rect 309554 166294 309622 166350
rect 309678 166294 327250 166350
rect 327306 166294 327374 166350
rect 327430 166294 327498 166350
rect 327554 166294 327622 166350
rect 327678 166294 345250 166350
rect 345306 166294 345374 166350
rect 345430 166294 345498 166350
rect 345554 166294 345622 166350
rect 345678 166294 363250 166350
rect 363306 166294 363374 166350
rect 363430 166294 363498 166350
rect 363554 166294 363622 166350
rect 363678 166294 381250 166350
rect 381306 166294 381374 166350
rect 381430 166294 381498 166350
rect 381554 166294 381622 166350
rect 381678 166294 399250 166350
rect 399306 166294 399374 166350
rect 399430 166294 399498 166350
rect 399554 166294 399622 166350
rect 399678 166294 417250 166350
rect 417306 166294 417374 166350
rect 417430 166294 417498 166350
rect 417554 166294 417622 166350
rect 417678 166294 435250 166350
rect 435306 166294 435374 166350
rect 435430 166294 435498 166350
rect 435554 166294 435622 166350
rect 435678 166294 453250 166350
rect 453306 166294 453374 166350
rect 453430 166294 453498 166350
rect 453554 166294 453622 166350
rect 453678 166294 471250 166350
rect 471306 166294 471374 166350
rect 471430 166294 471498 166350
rect 471554 166294 471622 166350
rect 471678 166294 489250 166350
rect 489306 166294 489374 166350
rect 489430 166294 489498 166350
rect 489554 166294 489622 166350
rect 489678 166294 507250 166350
rect 507306 166294 507374 166350
rect 507430 166294 507498 166350
rect 507554 166294 507622 166350
rect 507678 166294 525250 166350
rect 525306 166294 525374 166350
rect 525430 166294 525498 166350
rect 525554 166294 525622 166350
rect 525678 166294 543250 166350
rect 543306 166294 543374 166350
rect 543430 166294 543498 166350
rect 543554 166294 543622 166350
rect 543678 166294 561250 166350
rect 561306 166294 561374 166350
rect 561430 166294 561498 166350
rect 561554 166294 561622 166350
rect 561678 166294 579250 166350
rect 579306 166294 579374 166350
rect 579430 166294 579498 166350
rect 579554 166294 579622 166350
rect 579678 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 3250 166226
rect 3306 166170 3374 166226
rect 3430 166170 3498 166226
rect 3554 166170 3622 166226
rect 3678 166170 21250 166226
rect 21306 166170 21374 166226
rect 21430 166170 21498 166226
rect 21554 166170 21622 166226
rect 21678 166170 39250 166226
rect 39306 166170 39374 166226
rect 39430 166170 39498 166226
rect 39554 166170 39622 166226
rect 39678 166170 57250 166226
rect 57306 166170 57374 166226
rect 57430 166170 57498 166226
rect 57554 166170 57622 166226
rect 57678 166170 75250 166226
rect 75306 166170 75374 166226
rect 75430 166170 75498 166226
rect 75554 166170 75622 166226
rect 75678 166170 93250 166226
rect 93306 166170 93374 166226
rect 93430 166170 93498 166226
rect 93554 166170 93622 166226
rect 93678 166170 111250 166226
rect 111306 166170 111374 166226
rect 111430 166170 111498 166226
rect 111554 166170 111622 166226
rect 111678 166170 129250 166226
rect 129306 166170 129374 166226
rect 129430 166170 129498 166226
rect 129554 166170 129622 166226
rect 129678 166170 147250 166226
rect 147306 166170 147374 166226
rect 147430 166170 147498 166226
rect 147554 166170 147622 166226
rect 147678 166170 165250 166226
rect 165306 166170 165374 166226
rect 165430 166170 165498 166226
rect 165554 166170 165622 166226
rect 165678 166170 183250 166226
rect 183306 166170 183374 166226
rect 183430 166170 183498 166226
rect 183554 166170 183622 166226
rect 183678 166170 201250 166226
rect 201306 166170 201374 166226
rect 201430 166170 201498 166226
rect 201554 166170 201622 166226
rect 201678 166170 219250 166226
rect 219306 166170 219374 166226
rect 219430 166170 219498 166226
rect 219554 166170 219622 166226
rect 219678 166170 237250 166226
rect 237306 166170 237374 166226
rect 237430 166170 237498 166226
rect 237554 166170 237622 166226
rect 237678 166170 255250 166226
rect 255306 166170 255374 166226
rect 255430 166170 255498 166226
rect 255554 166170 255622 166226
rect 255678 166170 273250 166226
rect 273306 166170 273374 166226
rect 273430 166170 273498 166226
rect 273554 166170 273622 166226
rect 273678 166170 291250 166226
rect 291306 166170 291374 166226
rect 291430 166170 291498 166226
rect 291554 166170 291622 166226
rect 291678 166170 309250 166226
rect 309306 166170 309374 166226
rect 309430 166170 309498 166226
rect 309554 166170 309622 166226
rect 309678 166170 327250 166226
rect 327306 166170 327374 166226
rect 327430 166170 327498 166226
rect 327554 166170 327622 166226
rect 327678 166170 345250 166226
rect 345306 166170 345374 166226
rect 345430 166170 345498 166226
rect 345554 166170 345622 166226
rect 345678 166170 363250 166226
rect 363306 166170 363374 166226
rect 363430 166170 363498 166226
rect 363554 166170 363622 166226
rect 363678 166170 381250 166226
rect 381306 166170 381374 166226
rect 381430 166170 381498 166226
rect 381554 166170 381622 166226
rect 381678 166170 399250 166226
rect 399306 166170 399374 166226
rect 399430 166170 399498 166226
rect 399554 166170 399622 166226
rect 399678 166170 417250 166226
rect 417306 166170 417374 166226
rect 417430 166170 417498 166226
rect 417554 166170 417622 166226
rect 417678 166170 435250 166226
rect 435306 166170 435374 166226
rect 435430 166170 435498 166226
rect 435554 166170 435622 166226
rect 435678 166170 453250 166226
rect 453306 166170 453374 166226
rect 453430 166170 453498 166226
rect 453554 166170 453622 166226
rect 453678 166170 471250 166226
rect 471306 166170 471374 166226
rect 471430 166170 471498 166226
rect 471554 166170 471622 166226
rect 471678 166170 489250 166226
rect 489306 166170 489374 166226
rect 489430 166170 489498 166226
rect 489554 166170 489622 166226
rect 489678 166170 507250 166226
rect 507306 166170 507374 166226
rect 507430 166170 507498 166226
rect 507554 166170 507622 166226
rect 507678 166170 525250 166226
rect 525306 166170 525374 166226
rect 525430 166170 525498 166226
rect 525554 166170 525622 166226
rect 525678 166170 543250 166226
rect 543306 166170 543374 166226
rect 543430 166170 543498 166226
rect 543554 166170 543622 166226
rect 543678 166170 561250 166226
rect 561306 166170 561374 166226
rect 561430 166170 561498 166226
rect 561554 166170 561622 166226
rect 561678 166170 579250 166226
rect 579306 166170 579374 166226
rect 579430 166170 579498 166226
rect 579554 166170 579622 166226
rect 579678 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 3250 166102
rect 3306 166046 3374 166102
rect 3430 166046 3498 166102
rect 3554 166046 3622 166102
rect 3678 166046 21250 166102
rect 21306 166046 21374 166102
rect 21430 166046 21498 166102
rect 21554 166046 21622 166102
rect 21678 166046 39250 166102
rect 39306 166046 39374 166102
rect 39430 166046 39498 166102
rect 39554 166046 39622 166102
rect 39678 166046 57250 166102
rect 57306 166046 57374 166102
rect 57430 166046 57498 166102
rect 57554 166046 57622 166102
rect 57678 166046 75250 166102
rect 75306 166046 75374 166102
rect 75430 166046 75498 166102
rect 75554 166046 75622 166102
rect 75678 166046 93250 166102
rect 93306 166046 93374 166102
rect 93430 166046 93498 166102
rect 93554 166046 93622 166102
rect 93678 166046 111250 166102
rect 111306 166046 111374 166102
rect 111430 166046 111498 166102
rect 111554 166046 111622 166102
rect 111678 166046 129250 166102
rect 129306 166046 129374 166102
rect 129430 166046 129498 166102
rect 129554 166046 129622 166102
rect 129678 166046 147250 166102
rect 147306 166046 147374 166102
rect 147430 166046 147498 166102
rect 147554 166046 147622 166102
rect 147678 166046 165250 166102
rect 165306 166046 165374 166102
rect 165430 166046 165498 166102
rect 165554 166046 165622 166102
rect 165678 166046 183250 166102
rect 183306 166046 183374 166102
rect 183430 166046 183498 166102
rect 183554 166046 183622 166102
rect 183678 166046 201250 166102
rect 201306 166046 201374 166102
rect 201430 166046 201498 166102
rect 201554 166046 201622 166102
rect 201678 166046 219250 166102
rect 219306 166046 219374 166102
rect 219430 166046 219498 166102
rect 219554 166046 219622 166102
rect 219678 166046 237250 166102
rect 237306 166046 237374 166102
rect 237430 166046 237498 166102
rect 237554 166046 237622 166102
rect 237678 166046 255250 166102
rect 255306 166046 255374 166102
rect 255430 166046 255498 166102
rect 255554 166046 255622 166102
rect 255678 166046 273250 166102
rect 273306 166046 273374 166102
rect 273430 166046 273498 166102
rect 273554 166046 273622 166102
rect 273678 166046 291250 166102
rect 291306 166046 291374 166102
rect 291430 166046 291498 166102
rect 291554 166046 291622 166102
rect 291678 166046 309250 166102
rect 309306 166046 309374 166102
rect 309430 166046 309498 166102
rect 309554 166046 309622 166102
rect 309678 166046 327250 166102
rect 327306 166046 327374 166102
rect 327430 166046 327498 166102
rect 327554 166046 327622 166102
rect 327678 166046 345250 166102
rect 345306 166046 345374 166102
rect 345430 166046 345498 166102
rect 345554 166046 345622 166102
rect 345678 166046 363250 166102
rect 363306 166046 363374 166102
rect 363430 166046 363498 166102
rect 363554 166046 363622 166102
rect 363678 166046 381250 166102
rect 381306 166046 381374 166102
rect 381430 166046 381498 166102
rect 381554 166046 381622 166102
rect 381678 166046 399250 166102
rect 399306 166046 399374 166102
rect 399430 166046 399498 166102
rect 399554 166046 399622 166102
rect 399678 166046 417250 166102
rect 417306 166046 417374 166102
rect 417430 166046 417498 166102
rect 417554 166046 417622 166102
rect 417678 166046 435250 166102
rect 435306 166046 435374 166102
rect 435430 166046 435498 166102
rect 435554 166046 435622 166102
rect 435678 166046 453250 166102
rect 453306 166046 453374 166102
rect 453430 166046 453498 166102
rect 453554 166046 453622 166102
rect 453678 166046 471250 166102
rect 471306 166046 471374 166102
rect 471430 166046 471498 166102
rect 471554 166046 471622 166102
rect 471678 166046 489250 166102
rect 489306 166046 489374 166102
rect 489430 166046 489498 166102
rect 489554 166046 489622 166102
rect 489678 166046 507250 166102
rect 507306 166046 507374 166102
rect 507430 166046 507498 166102
rect 507554 166046 507622 166102
rect 507678 166046 525250 166102
rect 525306 166046 525374 166102
rect 525430 166046 525498 166102
rect 525554 166046 525622 166102
rect 525678 166046 543250 166102
rect 543306 166046 543374 166102
rect 543430 166046 543498 166102
rect 543554 166046 543622 166102
rect 543678 166046 561250 166102
rect 561306 166046 561374 166102
rect 561430 166046 561498 166102
rect 561554 166046 561622 166102
rect 561678 166046 579250 166102
rect 579306 166046 579374 166102
rect 579430 166046 579498 166102
rect 579554 166046 579622 166102
rect 579678 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 3250 165978
rect 3306 165922 3374 165978
rect 3430 165922 3498 165978
rect 3554 165922 3622 165978
rect 3678 165922 21250 165978
rect 21306 165922 21374 165978
rect 21430 165922 21498 165978
rect 21554 165922 21622 165978
rect 21678 165922 39250 165978
rect 39306 165922 39374 165978
rect 39430 165922 39498 165978
rect 39554 165922 39622 165978
rect 39678 165922 57250 165978
rect 57306 165922 57374 165978
rect 57430 165922 57498 165978
rect 57554 165922 57622 165978
rect 57678 165922 75250 165978
rect 75306 165922 75374 165978
rect 75430 165922 75498 165978
rect 75554 165922 75622 165978
rect 75678 165922 93250 165978
rect 93306 165922 93374 165978
rect 93430 165922 93498 165978
rect 93554 165922 93622 165978
rect 93678 165922 111250 165978
rect 111306 165922 111374 165978
rect 111430 165922 111498 165978
rect 111554 165922 111622 165978
rect 111678 165922 129250 165978
rect 129306 165922 129374 165978
rect 129430 165922 129498 165978
rect 129554 165922 129622 165978
rect 129678 165922 147250 165978
rect 147306 165922 147374 165978
rect 147430 165922 147498 165978
rect 147554 165922 147622 165978
rect 147678 165922 165250 165978
rect 165306 165922 165374 165978
rect 165430 165922 165498 165978
rect 165554 165922 165622 165978
rect 165678 165922 183250 165978
rect 183306 165922 183374 165978
rect 183430 165922 183498 165978
rect 183554 165922 183622 165978
rect 183678 165922 201250 165978
rect 201306 165922 201374 165978
rect 201430 165922 201498 165978
rect 201554 165922 201622 165978
rect 201678 165922 219250 165978
rect 219306 165922 219374 165978
rect 219430 165922 219498 165978
rect 219554 165922 219622 165978
rect 219678 165922 237250 165978
rect 237306 165922 237374 165978
rect 237430 165922 237498 165978
rect 237554 165922 237622 165978
rect 237678 165922 255250 165978
rect 255306 165922 255374 165978
rect 255430 165922 255498 165978
rect 255554 165922 255622 165978
rect 255678 165922 273250 165978
rect 273306 165922 273374 165978
rect 273430 165922 273498 165978
rect 273554 165922 273622 165978
rect 273678 165922 291250 165978
rect 291306 165922 291374 165978
rect 291430 165922 291498 165978
rect 291554 165922 291622 165978
rect 291678 165922 309250 165978
rect 309306 165922 309374 165978
rect 309430 165922 309498 165978
rect 309554 165922 309622 165978
rect 309678 165922 327250 165978
rect 327306 165922 327374 165978
rect 327430 165922 327498 165978
rect 327554 165922 327622 165978
rect 327678 165922 345250 165978
rect 345306 165922 345374 165978
rect 345430 165922 345498 165978
rect 345554 165922 345622 165978
rect 345678 165922 363250 165978
rect 363306 165922 363374 165978
rect 363430 165922 363498 165978
rect 363554 165922 363622 165978
rect 363678 165922 381250 165978
rect 381306 165922 381374 165978
rect 381430 165922 381498 165978
rect 381554 165922 381622 165978
rect 381678 165922 399250 165978
rect 399306 165922 399374 165978
rect 399430 165922 399498 165978
rect 399554 165922 399622 165978
rect 399678 165922 417250 165978
rect 417306 165922 417374 165978
rect 417430 165922 417498 165978
rect 417554 165922 417622 165978
rect 417678 165922 435250 165978
rect 435306 165922 435374 165978
rect 435430 165922 435498 165978
rect 435554 165922 435622 165978
rect 435678 165922 453250 165978
rect 453306 165922 453374 165978
rect 453430 165922 453498 165978
rect 453554 165922 453622 165978
rect 453678 165922 471250 165978
rect 471306 165922 471374 165978
rect 471430 165922 471498 165978
rect 471554 165922 471622 165978
rect 471678 165922 489250 165978
rect 489306 165922 489374 165978
rect 489430 165922 489498 165978
rect 489554 165922 489622 165978
rect 489678 165922 507250 165978
rect 507306 165922 507374 165978
rect 507430 165922 507498 165978
rect 507554 165922 507622 165978
rect 507678 165922 525250 165978
rect 525306 165922 525374 165978
rect 525430 165922 525498 165978
rect 525554 165922 525622 165978
rect 525678 165922 543250 165978
rect 543306 165922 543374 165978
rect 543430 165922 543498 165978
rect 543554 165922 543622 165978
rect 543678 165922 561250 165978
rect 561306 165922 561374 165978
rect 561430 165922 561498 165978
rect 561554 165922 561622 165978
rect 561678 165922 579250 165978
rect 579306 165922 579374 165978
rect 579430 165922 579498 165978
rect 579554 165922 579622 165978
rect 579678 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 6970 154350
rect 7026 154294 7094 154350
rect 7150 154294 7218 154350
rect 7274 154294 7342 154350
rect 7398 154294 24970 154350
rect 25026 154294 25094 154350
rect 25150 154294 25218 154350
rect 25274 154294 25342 154350
rect 25398 154294 42970 154350
rect 43026 154294 43094 154350
rect 43150 154294 43218 154350
rect 43274 154294 43342 154350
rect 43398 154294 60970 154350
rect 61026 154294 61094 154350
rect 61150 154294 61218 154350
rect 61274 154294 61342 154350
rect 61398 154294 78970 154350
rect 79026 154294 79094 154350
rect 79150 154294 79218 154350
rect 79274 154294 79342 154350
rect 79398 154294 96970 154350
rect 97026 154294 97094 154350
rect 97150 154294 97218 154350
rect 97274 154294 97342 154350
rect 97398 154294 114970 154350
rect 115026 154294 115094 154350
rect 115150 154294 115218 154350
rect 115274 154294 115342 154350
rect 115398 154294 132970 154350
rect 133026 154294 133094 154350
rect 133150 154294 133218 154350
rect 133274 154294 133342 154350
rect 133398 154294 150970 154350
rect 151026 154294 151094 154350
rect 151150 154294 151218 154350
rect 151274 154294 151342 154350
rect 151398 154294 168970 154350
rect 169026 154294 169094 154350
rect 169150 154294 169218 154350
rect 169274 154294 169342 154350
rect 169398 154294 186970 154350
rect 187026 154294 187094 154350
rect 187150 154294 187218 154350
rect 187274 154294 187342 154350
rect 187398 154294 204970 154350
rect 205026 154294 205094 154350
rect 205150 154294 205218 154350
rect 205274 154294 205342 154350
rect 205398 154294 222970 154350
rect 223026 154294 223094 154350
rect 223150 154294 223218 154350
rect 223274 154294 223342 154350
rect 223398 154294 240970 154350
rect 241026 154294 241094 154350
rect 241150 154294 241218 154350
rect 241274 154294 241342 154350
rect 241398 154294 258970 154350
rect 259026 154294 259094 154350
rect 259150 154294 259218 154350
rect 259274 154294 259342 154350
rect 259398 154294 276970 154350
rect 277026 154294 277094 154350
rect 277150 154294 277218 154350
rect 277274 154294 277342 154350
rect 277398 154294 294970 154350
rect 295026 154294 295094 154350
rect 295150 154294 295218 154350
rect 295274 154294 295342 154350
rect 295398 154294 312970 154350
rect 313026 154294 313094 154350
rect 313150 154294 313218 154350
rect 313274 154294 313342 154350
rect 313398 154294 330970 154350
rect 331026 154294 331094 154350
rect 331150 154294 331218 154350
rect 331274 154294 331342 154350
rect 331398 154294 348970 154350
rect 349026 154294 349094 154350
rect 349150 154294 349218 154350
rect 349274 154294 349342 154350
rect 349398 154294 366970 154350
rect 367026 154294 367094 154350
rect 367150 154294 367218 154350
rect 367274 154294 367342 154350
rect 367398 154294 384970 154350
rect 385026 154294 385094 154350
rect 385150 154294 385218 154350
rect 385274 154294 385342 154350
rect 385398 154294 402970 154350
rect 403026 154294 403094 154350
rect 403150 154294 403218 154350
rect 403274 154294 403342 154350
rect 403398 154294 420970 154350
rect 421026 154294 421094 154350
rect 421150 154294 421218 154350
rect 421274 154294 421342 154350
rect 421398 154294 438970 154350
rect 439026 154294 439094 154350
rect 439150 154294 439218 154350
rect 439274 154294 439342 154350
rect 439398 154294 456970 154350
rect 457026 154294 457094 154350
rect 457150 154294 457218 154350
rect 457274 154294 457342 154350
rect 457398 154294 474970 154350
rect 475026 154294 475094 154350
rect 475150 154294 475218 154350
rect 475274 154294 475342 154350
rect 475398 154294 492970 154350
rect 493026 154294 493094 154350
rect 493150 154294 493218 154350
rect 493274 154294 493342 154350
rect 493398 154294 510970 154350
rect 511026 154294 511094 154350
rect 511150 154294 511218 154350
rect 511274 154294 511342 154350
rect 511398 154294 528970 154350
rect 529026 154294 529094 154350
rect 529150 154294 529218 154350
rect 529274 154294 529342 154350
rect 529398 154294 546970 154350
rect 547026 154294 547094 154350
rect 547150 154294 547218 154350
rect 547274 154294 547342 154350
rect 547398 154294 564970 154350
rect 565026 154294 565094 154350
rect 565150 154294 565218 154350
rect 565274 154294 565342 154350
rect 565398 154294 582970 154350
rect 583026 154294 583094 154350
rect 583150 154294 583218 154350
rect 583274 154294 583342 154350
rect 583398 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 6970 154226
rect 7026 154170 7094 154226
rect 7150 154170 7218 154226
rect 7274 154170 7342 154226
rect 7398 154170 24970 154226
rect 25026 154170 25094 154226
rect 25150 154170 25218 154226
rect 25274 154170 25342 154226
rect 25398 154170 42970 154226
rect 43026 154170 43094 154226
rect 43150 154170 43218 154226
rect 43274 154170 43342 154226
rect 43398 154170 60970 154226
rect 61026 154170 61094 154226
rect 61150 154170 61218 154226
rect 61274 154170 61342 154226
rect 61398 154170 78970 154226
rect 79026 154170 79094 154226
rect 79150 154170 79218 154226
rect 79274 154170 79342 154226
rect 79398 154170 96970 154226
rect 97026 154170 97094 154226
rect 97150 154170 97218 154226
rect 97274 154170 97342 154226
rect 97398 154170 114970 154226
rect 115026 154170 115094 154226
rect 115150 154170 115218 154226
rect 115274 154170 115342 154226
rect 115398 154170 132970 154226
rect 133026 154170 133094 154226
rect 133150 154170 133218 154226
rect 133274 154170 133342 154226
rect 133398 154170 150970 154226
rect 151026 154170 151094 154226
rect 151150 154170 151218 154226
rect 151274 154170 151342 154226
rect 151398 154170 168970 154226
rect 169026 154170 169094 154226
rect 169150 154170 169218 154226
rect 169274 154170 169342 154226
rect 169398 154170 186970 154226
rect 187026 154170 187094 154226
rect 187150 154170 187218 154226
rect 187274 154170 187342 154226
rect 187398 154170 204970 154226
rect 205026 154170 205094 154226
rect 205150 154170 205218 154226
rect 205274 154170 205342 154226
rect 205398 154170 222970 154226
rect 223026 154170 223094 154226
rect 223150 154170 223218 154226
rect 223274 154170 223342 154226
rect 223398 154170 240970 154226
rect 241026 154170 241094 154226
rect 241150 154170 241218 154226
rect 241274 154170 241342 154226
rect 241398 154170 258970 154226
rect 259026 154170 259094 154226
rect 259150 154170 259218 154226
rect 259274 154170 259342 154226
rect 259398 154170 276970 154226
rect 277026 154170 277094 154226
rect 277150 154170 277218 154226
rect 277274 154170 277342 154226
rect 277398 154170 294970 154226
rect 295026 154170 295094 154226
rect 295150 154170 295218 154226
rect 295274 154170 295342 154226
rect 295398 154170 312970 154226
rect 313026 154170 313094 154226
rect 313150 154170 313218 154226
rect 313274 154170 313342 154226
rect 313398 154170 330970 154226
rect 331026 154170 331094 154226
rect 331150 154170 331218 154226
rect 331274 154170 331342 154226
rect 331398 154170 348970 154226
rect 349026 154170 349094 154226
rect 349150 154170 349218 154226
rect 349274 154170 349342 154226
rect 349398 154170 366970 154226
rect 367026 154170 367094 154226
rect 367150 154170 367218 154226
rect 367274 154170 367342 154226
rect 367398 154170 384970 154226
rect 385026 154170 385094 154226
rect 385150 154170 385218 154226
rect 385274 154170 385342 154226
rect 385398 154170 402970 154226
rect 403026 154170 403094 154226
rect 403150 154170 403218 154226
rect 403274 154170 403342 154226
rect 403398 154170 420970 154226
rect 421026 154170 421094 154226
rect 421150 154170 421218 154226
rect 421274 154170 421342 154226
rect 421398 154170 438970 154226
rect 439026 154170 439094 154226
rect 439150 154170 439218 154226
rect 439274 154170 439342 154226
rect 439398 154170 456970 154226
rect 457026 154170 457094 154226
rect 457150 154170 457218 154226
rect 457274 154170 457342 154226
rect 457398 154170 474970 154226
rect 475026 154170 475094 154226
rect 475150 154170 475218 154226
rect 475274 154170 475342 154226
rect 475398 154170 492970 154226
rect 493026 154170 493094 154226
rect 493150 154170 493218 154226
rect 493274 154170 493342 154226
rect 493398 154170 510970 154226
rect 511026 154170 511094 154226
rect 511150 154170 511218 154226
rect 511274 154170 511342 154226
rect 511398 154170 528970 154226
rect 529026 154170 529094 154226
rect 529150 154170 529218 154226
rect 529274 154170 529342 154226
rect 529398 154170 546970 154226
rect 547026 154170 547094 154226
rect 547150 154170 547218 154226
rect 547274 154170 547342 154226
rect 547398 154170 564970 154226
rect 565026 154170 565094 154226
rect 565150 154170 565218 154226
rect 565274 154170 565342 154226
rect 565398 154170 582970 154226
rect 583026 154170 583094 154226
rect 583150 154170 583218 154226
rect 583274 154170 583342 154226
rect 583398 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 6970 154102
rect 7026 154046 7094 154102
rect 7150 154046 7218 154102
rect 7274 154046 7342 154102
rect 7398 154046 24970 154102
rect 25026 154046 25094 154102
rect 25150 154046 25218 154102
rect 25274 154046 25342 154102
rect 25398 154046 42970 154102
rect 43026 154046 43094 154102
rect 43150 154046 43218 154102
rect 43274 154046 43342 154102
rect 43398 154046 60970 154102
rect 61026 154046 61094 154102
rect 61150 154046 61218 154102
rect 61274 154046 61342 154102
rect 61398 154046 78970 154102
rect 79026 154046 79094 154102
rect 79150 154046 79218 154102
rect 79274 154046 79342 154102
rect 79398 154046 96970 154102
rect 97026 154046 97094 154102
rect 97150 154046 97218 154102
rect 97274 154046 97342 154102
rect 97398 154046 114970 154102
rect 115026 154046 115094 154102
rect 115150 154046 115218 154102
rect 115274 154046 115342 154102
rect 115398 154046 132970 154102
rect 133026 154046 133094 154102
rect 133150 154046 133218 154102
rect 133274 154046 133342 154102
rect 133398 154046 150970 154102
rect 151026 154046 151094 154102
rect 151150 154046 151218 154102
rect 151274 154046 151342 154102
rect 151398 154046 168970 154102
rect 169026 154046 169094 154102
rect 169150 154046 169218 154102
rect 169274 154046 169342 154102
rect 169398 154046 186970 154102
rect 187026 154046 187094 154102
rect 187150 154046 187218 154102
rect 187274 154046 187342 154102
rect 187398 154046 204970 154102
rect 205026 154046 205094 154102
rect 205150 154046 205218 154102
rect 205274 154046 205342 154102
rect 205398 154046 222970 154102
rect 223026 154046 223094 154102
rect 223150 154046 223218 154102
rect 223274 154046 223342 154102
rect 223398 154046 240970 154102
rect 241026 154046 241094 154102
rect 241150 154046 241218 154102
rect 241274 154046 241342 154102
rect 241398 154046 258970 154102
rect 259026 154046 259094 154102
rect 259150 154046 259218 154102
rect 259274 154046 259342 154102
rect 259398 154046 276970 154102
rect 277026 154046 277094 154102
rect 277150 154046 277218 154102
rect 277274 154046 277342 154102
rect 277398 154046 294970 154102
rect 295026 154046 295094 154102
rect 295150 154046 295218 154102
rect 295274 154046 295342 154102
rect 295398 154046 312970 154102
rect 313026 154046 313094 154102
rect 313150 154046 313218 154102
rect 313274 154046 313342 154102
rect 313398 154046 330970 154102
rect 331026 154046 331094 154102
rect 331150 154046 331218 154102
rect 331274 154046 331342 154102
rect 331398 154046 348970 154102
rect 349026 154046 349094 154102
rect 349150 154046 349218 154102
rect 349274 154046 349342 154102
rect 349398 154046 366970 154102
rect 367026 154046 367094 154102
rect 367150 154046 367218 154102
rect 367274 154046 367342 154102
rect 367398 154046 384970 154102
rect 385026 154046 385094 154102
rect 385150 154046 385218 154102
rect 385274 154046 385342 154102
rect 385398 154046 402970 154102
rect 403026 154046 403094 154102
rect 403150 154046 403218 154102
rect 403274 154046 403342 154102
rect 403398 154046 420970 154102
rect 421026 154046 421094 154102
rect 421150 154046 421218 154102
rect 421274 154046 421342 154102
rect 421398 154046 438970 154102
rect 439026 154046 439094 154102
rect 439150 154046 439218 154102
rect 439274 154046 439342 154102
rect 439398 154046 456970 154102
rect 457026 154046 457094 154102
rect 457150 154046 457218 154102
rect 457274 154046 457342 154102
rect 457398 154046 474970 154102
rect 475026 154046 475094 154102
rect 475150 154046 475218 154102
rect 475274 154046 475342 154102
rect 475398 154046 492970 154102
rect 493026 154046 493094 154102
rect 493150 154046 493218 154102
rect 493274 154046 493342 154102
rect 493398 154046 510970 154102
rect 511026 154046 511094 154102
rect 511150 154046 511218 154102
rect 511274 154046 511342 154102
rect 511398 154046 528970 154102
rect 529026 154046 529094 154102
rect 529150 154046 529218 154102
rect 529274 154046 529342 154102
rect 529398 154046 546970 154102
rect 547026 154046 547094 154102
rect 547150 154046 547218 154102
rect 547274 154046 547342 154102
rect 547398 154046 564970 154102
rect 565026 154046 565094 154102
rect 565150 154046 565218 154102
rect 565274 154046 565342 154102
rect 565398 154046 582970 154102
rect 583026 154046 583094 154102
rect 583150 154046 583218 154102
rect 583274 154046 583342 154102
rect 583398 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 6970 153978
rect 7026 153922 7094 153978
rect 7150 153922 7218 153978
rect 7274 153922 7342 153978
rect 7398 153922 24970 153978
rect 25026 153922 25094 153978
rect 25150 153922 25218 153978
rect 25274 153922 25342 153978
rect 25398 153922 42970 153978
rect 43026 153922 43094 153978
rect 43150 153922 43218 153978
rect 43274 153922 43342 153978
rect 43398 153922 60970 153978
rect 61026 153922 61094 153978
rect 61150 153922 61218 153978
rect 61274 153922 61342 153978
rect 61398 153922 78970 153978
rect 79026 153922 79094 153978
rect 79150 153922 79218 153978
rect 79274 153922 79342 153978
rect 79398 153922 96970 153978
rect 97026 153922 97094 153978
rect 97150 153922 97218 153978
rect 97274 153922 97342 153978
rect 97398 153922 114970 153978
rect 115026 153922 115094 153978
rect 115150 153922 115218 153978
rect 115274 153922 115342 153978
rect 115398 153922 132970 153978
rect 133026 153922 133094 153978
rect 133150 153922 133218 153978
rect 133274 153922 133342 153978
rect 133398 153922 150970 153978
rect 151026 153922 151094 153978
rect 151150 153922 151218 153978
rect 151274 153922 151342 153978
rect 151398 153922 168970 153978
rect 169026 153922 169094 153978
rect 169150 153922 169218 153978
rect 169274 153922 169342 153978
rect 169398 153922 186970 153978
rect 187026 153922 187094 153978
rect 187150 153922 187218 153978
rect 187274 153922 187342 153978
rect 187398 153922 204970 153978
rect 205026 153922 205094 153978
rect 205150 153922 205218 153978
rect 205274 153922 205342 153978
rect 205398 153922 222970 153978
rect 223026 153922 223094 153978
rect 223150 153922 223218 153978
rect 223274 153922 223342 153978
rect 223398 153922 240970 153978
rect 241026 153922 241094 153978
rect 241150 153922 241218 153978
rect 241274 153922 241342 153978
rect 241398 153922 258970 153978
rect 259026 153922 259094 153978
rect 259150 153922 259218 153978
rect 259274 153922 259342 153978
rect 259398 153922 276970 153978
rect 277026 153922 277094 153978
rect 277150 153922 277218 153978
rect 277274 153922 277342 153978
rect 277398 153922 294970 153978
rect 295026 153922 295094 153978
rect 295150 153922 295218 153978
rect 295274 153922 295342 153978
rect 295398 153922 312970 153978
rect 313026 153922 313094 153978
rect 313150 153922 313218 153978
rect 313274 153922 313342 153978
rect 313398 153922 330970 153978
rect 331026 153922 331094 153978
rect 331150 153922 331218 153978
rect 331274 153922 331342 153978
rect 331398 153922 348970 153978
rect 349026 153922 349094 153978
rect 349150 153922 349218 153978
rect 349274 153922 349342 153978
rect 349398 153922 366970 153978
rect 367026 153922 367094 153978
rect 367150 153922 367218 153978
rect 367274 153922 367342 153978
rect 367398 153922 384970 153978
rect 385026 153922 385094 153978
rect 385150 153922 385218 153978
rect 385274 153922 385342 153978
rect 385398 153922 402970 153978
rect 403026 153922 403094 153978
rect 403150 153922 403218 153978
rect 403274 153922 403342 153978
rect 403398 153922 420970 153978
rect 421026 153922 421094 153978
rect 421150 153922 421218 153978
rect 421274 153922 421342 153978
rect 421398 153922 438970 153978
rect 439026 153922 439094 153978
rect 439150 153922 439218 153978
rect 439274 153922 439342 153978
rect 439398 153922 456970 153978
rect 457026 153922 457094 153978
rect 457150 153922 457218 153978
rect 457274 153922 457342 153978
rect 457398 153922 474970 153978
rect 475026 153922 475094 153978
rect 475150 153922 475218 153978
rect 475274 153922 475342 153978
rect 475398 153922 492970 153978
rect 493026 153922 493094 153978
rect 493150 153922 493218 153978
rect 493274 153922 493342 153978
rect 493398 153922 510970 153978
rect 511026 153922 511094 153978
rect 511150 153922 511218 153978
rect 511274 153922 511342 153978
rect 511398 153922 528970 153978
rect 529026 153922 529094 153978
rect 529150 153922 529218 153978
rect 529274 153922 529342 153978
rect 529398 153922 546970 153978
rect 547026 153922 547094 153978
rect 547150 153922 547218 153978
rect 547274 153922 547342 153978
rect 547398 153922 564970 153978
rect 565026 153922 565094 153978
rect 565150 153922 565218 153978
rect 565274 153922 565342 153978
rect 565398 153922 582970 153978
rect 583026 153922 583094 153978
rect 583150 153922 583218 153978
rect 583274 153922 583342 153978
rect 583398 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 3250 148350
rect 3306 148294 3374 148350
rect 3430 148294 3498 148350
rect 3554 148294 3622 148350
rect 3678 148294 21250 148350
rect 21306 148294 21374 148350
rect 21430 148294 21498 148350
rect 21554 148294 21622 148350
rect 21678 148294 39250 148350
rect 39306 148294 39374 148350
rect 39430 148294 39498 148350
rect 39554 148294 39622 148350
rect 39678 148294 57250 148350
rect 57306 148294 57374 148350
rect 57430 148294 57498 148350
rect 57554 148294 57622 148350
rect 57678 148294 75250 148350
rect 75306 148294 75374 148350
rect 75430 148294 75498 148350
rect 75554 148294 75622 148350
rect 75678 148294 93250 148350
rect 93306 148294 93374 148350
rect 93430 148294 93498 148350
rect 93554 148294 93622 148350
rect 93678 148294 111250 148350
rect 111306 148294 111374 148350
rect 111430 148294 111498 148350
rect 111554 148294 111622 148350
rect 111678 148294 129250 148350
rect 129306 148294 129374 148350
rect 129430 148294 129498 148350
rect 129554 148294 129622 148350
rect 129678 148294 147250 148350
rect 147306 148294 147374 148350
rect 147430 148294 147498 148350
rect 147554 148294 147622 148350
rect 147678 148294 165250 148350
rect 165306 148294 165374 148350
rect 165430 148294 165498 148350
rect 165554 148294 165622 148350
rect 165678 148294 183250 148350
rect 183306 148294 183374 148350
rect 183430 148294 183498 148350
rect 183554 148294 183622 148350
rect 183678 148294 201250 148350
rect 201306 148294 201374 148350
rect 201430 148294 201498 148350
rect 201554 148294 201622 148350
rect 201678 148294 219250 148350
rect 219306 148294 219374 148350
rect 219430 148294 219498 148350
rect 219554 148294 219622 148350
rect 219678 148294 237250 148350
rect 237306 148294 237374 148350
rect 237430 148294 237498 148350
rect 237554 148294 237622 148350
rect 237678 148294 255250 148350
rect 255306 148294 255374 148350
rect 255430 148294 255498 148350
rect 255554 148294 255622 148350
rect 255678 148294 273250 148350
rect 273306 148294 273374 148350
rect 273430 148294 273498 148350
rect 273554 148294 273622 148350
rect 273678 148294 291250 148350
rect 291306 148294 291374 148350
rect 291430 148294 291498 148350
rect 291554 148294 291622 148350
rect 291678 148294 309250 148350
rect 309306 148294 309374 148350
rect 309430 148294 309498 148350
rect 309554 148294 309622 148350
rect 309678 148294 327250 148350
rect 327306 148294 327374 148350
rect 327430 148294 327498 148350
rect 327554 148294 327622 148350
rect 327678 148294 345250 148350
rect 345306 148294 345374 148350
rect 345430 148294 345498 148350
rect 345554 148294 345622 148350
rect 345678 148294 363250 148350
rect 363306 148294 363374 148350
rect 363430 148294 363498 148350
rect 363554 148294 363622 148350
rect 363678 148294 381250 148350
rect 381306 148294 381374 148350
rect 381430 148294 381498 148350
rect 381554 148294 381622 148350
rect 381678 148294 399250 148350
rect 399306 148294 399374 148350
rect 399430 148294 399498 148350
rect 399554 148294 399622 148350
rect 399678 148294 417250 148350
rect 417306 148294 417374 148350
rect 417430 148294 417498 148350
rect 417554 148294 417622 148350
rect 417678 148294 435250 148350
rect 435306 148294 435374 148350
rect 435430 148294 435498 148350
rect 435554 148294 435622 148350
rect 435678 148294 453250 148350
rect 453306 148294 453374 148350
rect 453430 148294 453498 148350
rect 453554 148294 453622 148350
rect 453678 148294 471250 148350
rect 471306 148294 471374 148350
rect 471430 148294 471498 148350
rect 471554 148294 471622 148350
rect 471678 148294 489250 148350
rect 489306 148294 489374 148350
rect 489430 148294 489498 148350
rect 489554 148294 489622 148350
rect 489678 148294 507250 148350
rect 507306 148294 507374 148350
rect 507430 148294 507498 148350
rect 507554 148294 507622 148350
rect 507678 148294 525250 148350
rect 525306 148294 525374 148350
rect 525430 148294 525498 148350
rect 525554 148294 525622 148350
rect 525678 148294 543250 148350
rect 543306 148294 543374 148350
rect 543430 148294 543498 148350
rect 543554 148294 543622 148350
rect 543678 148294 561250 148350
rect 561306 148294 561374 148350
rect 561430 148294 561498 148350
rect 561554 148294 561622 148350
rect 561678 148294 579250 148350
rect 579306 148294 579374 148350
rect 579430 148294 579498 148350
rect 579554 148294 579622 148350
rect 579678 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 3250 148226
rect 3306 148170 3374 148226
rect 3430 148170 3498 148226
rect 3554 148170 3622 148226
rect 3678 148170 21250 148226
rect 21306 148170 21374 148226
rect 21430 148170 21498 148226
rect 21554 148170 21622 148226
rect 21678 148170 39250 148226
rect 39306 148170 39374 148226
rect 39430 148170 39498 148226
rect 39554 148170 39622 148226
rect 39678 148170 57250 148226
rect 57306 148170 57374 148226
rect 57430 148170 57498 148226
rect 57554 148170 57622 148226
rect 57678 148170 75250 148226
rect 75306 148170 75374 148226
rect 75430 148170 75498 148226
rect 75554 148170 75622 148226
rect 75678 148170 93250 148226
rect 93306 148170 93374 148226
rect 93430 148170 93498 148226
rect 93554 148170 93622 148226
rect 93678 148170 111250 148226
rect 111306 148170 111374 148226
rect 111430 148170 111498 148226
rect 111554 148170 111622 148226
rect 111678 148170 129250 148226
rect 129306 148170 129374 148226
rect 129430 148170 129498 148226
rect 129554 148170 129622 148226
rect 129678 148170 147250 148226
rect 147306 148170 147374 148226
rect 147430 148170 147498 148226
rect 147554 148170 147622 148226
rect 147678 148170 165250 148226
rect 165306 148170 165374 148226
rect 165430 148170 165498 148226
rect 165554 148170 165622 148226
rect 165678 148170 183250 148226
rect 183306 148170 183374 148226
rect 183430 148170 183498 148226
rect 183554 148170 183622 148226
rect 183678 148170 201250 148226
rect 201306 148170 201374 148226
rect 201430 148170 201498 148226
rect 201554 148170 201622 148226
rect 201678 148170 219250 148226
rect 219306 148170 219374 148226
rect 219430 148170 219498 148226
rect 219554 148170 219622 148226
rect 219678 148170 237250 148226
rect 237306 148170 237374 148226
rect 237430 148170 237498 148226
rect 237554 148170 237622 148226
rect 237678 148170 255250 148226
rect 255306 148170 255374 148226
rect 255430 148170 255498 148226
rect 255554 148170 255622 148226
rect 255678 148170 273250 148226
rect 273306 148170 273374 148226
rect 273430 148170 273498 148226
rect 273554 148170 273622 148226
rect 273678 148170 291250 148226
rect 291306 148170 291374 148226
rect 291430 148170 291498 148226
rect 291554 148170 291622 148226
rect 291678 148170 309250 148226
rect 309306 148170 309374 148226
rect 309430 148170 309498 148226
rect 309554 148170 309622 148226
rect 309678 148170 327250 148226
rect 327306 148170 327374 148226
rect 327430 148170 327498 148226
rect 327554 148170 327622 148226
rect 327678 148170 345250 148226
rect 345306 148170 345374 148226
rect 345430 148170 345498 148226
rect 345554 148170 345622 148226
rect 345678 148170 363250 148226
rect 363306 148170 363374 148226
rect 363430 148170 363498 148226
rect 363554 148170 363622 148226
rect 363678 148170 381250 148226
rect 381306 148170 381374 148226
rect 381430 148170 381498 148226
rect 381554 148170 381622 148226
rect 381678 148170 399250 148226
rect 399306 148170 399374 148226
rect 399430 148170 399498 148226
rect 399554 148170 399622 148226
rect 399678 148170 417250 148226
rect 417306 148170 417374 148226
rect 417430 148170 417498 148226
rect 417554 148170 417622 148226
rect 417678 148170 435250 148226
rect 435306 148170 435374 148226
rect 435430 148170 435498 148226
rect 435554 148170 435622 148226
rect 435678 148170 453250 148226
rect 453306 148170 453374 148226
rect 453430 148170 453498 148226
rect 453554 148170 453622 148226
rect 453678 148170 471250 148226
rect 471306 148170 471374 148226
rect 471430 148170 471498 148226
rect 471554 148170 471622 148226
rect 471678 148170 489250 148226
rect 489306 148170 489374 148226
rect 489430 148170 489498 148226
rect 489554 148170 489622 148226
rect 489678 148170 507250 148226
rect 507306 148170 507374 148226
rect 507430 148170 507498 148226
rect 507554 148170 507622 148226
rect 507678 148170 525250 148226
rect 525306 148170 525374 148226
rect 525430 148170 525498 148226
rect 525554 148170 525622 148226
rect 525678 148170 543250 148226
rect 543306 148170 543374 148226
rect 543430 148170 543498 148226
rect 543554 148170 543622 148226
rect 543678 148170 561250 148226
rect 561306 148170 561374 148226
rect 561430 148170 561498 148226
rect 561554 148170 561622 148226
rect 561678 148170 579250 148226
rect 579306 148170 579374 148226
rect 579430 148170 579498 148226
rect 579554 148170 579622 148226
rect 579678 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 3250 148102
rect 3306 148046 3374 148102
rect 3430 148046 3498 148102
rect 3554 148046 3622 148102
rect 3678 148046 21250 148102
rect 21306 148046 21374 148102
rect 21430 148046 21498 148102
rect 21554 148046 21622 148102
rect 21678 148046 39250 148102
rect 39306 148046 39374 148102
rect 39430 148046 39498 148102
rect 39554 148046 39622 148102
rect 39678 148046 57250 148102
rect 57306 148046 57374 148102
rect 57430 148046 57498 148102
rect 57554 148046 57622 148102
rect 57678 148046 75250 148102
rect 75306 148046 75374 148102
rect 75430 148046 75498 148102
rect 75554 148046 75622 148102
rect 75678 148046 93250 148102
rect 93306 148046 93374 148102
rect 93430 148046 93498 148102
rect 93554 148046 93622 148102
rect 93678 148046 111250 148102
rect 111306 148046 111374 148102
rect 111430 148046 111498 148102
rect 111554 148046 111622 148102
rect 111678 148046 129250 148102
rect 129306 148046 129374 148102
rect 129430 148046 129498 148102
rect 129554 148046 129622 148102
rect 129678 148046 147250 148102
rect 147306 148046 147374 148102
rect 147430 148046 147498 148102
rect 147554 148046 147622 148102
rect 147678 148046 165250 148102
rect 165306 148046 165374 148102
rect 165430 148046 165498 148102
rect 165554 148046 165622 148102
rect 165678 148046 183250 148102
rect 183306 148046 183374 148102
rect 183430 148046 183498 148102
rect 183554 148046 183622 148102
rect 183678 148046 201250 148102
rect 201306 148046 201374 148102
rect 201430 148046 201498 148102
rect 201554 148046 201622 148102
rect 201678 148046 219250 148102
rect 219306 148046 219374 148102
rect 219430 148046 219498 148102
rect 219554 148046 219622 148102
rect 219678 148046 237250 148102
rect 237306 148046 237374 148102
rect 237430 148046 237498 148102
rect 237554 148046 237622 148102
rect 237678 148046 255250 148102
rect 255306 148046 255374 148102
rect 255430 148046 255498 148102
rect 255554 148046 255622 148102
rect 255678 148046 273250 148102
rect 273306 148046 273374 148102
rect 273430 148046 273498 148102
rect 273554 148046 273622 148102
rect 273678 148046 291250 148102
rect 291306 148046 291374 148102
rect 291430 148046 291498 148102
rect 291554 148046 291622 148102
rect 291678 148046 309250 148102
rect 309306 148046 309374 148102
rect 309430 148046 309498 148102
rect 309554 148046 309622 148102
rect 309678 148046 327250 148102
rect 327306 148046 327374 148102
rect 327430 148046 327498 148102
rect 327554 148046 327622 148102
rect 327678 148046 345250 148102
rect 345306 148046 345374 148102
rect 345430 148046 345498 148102
rect 345554 148046 345622 148102
rect 345678 148046 363250 148102
rect 363306 148046 363374 148102
rect 363430 148046 363498 148102
rect 363554 148046 363622 148102
rect 363678 148046 381250 148102
rect 381306 148046 381374 148102
rect 381430 148046 381498 148102
rect 381554 148046 381622 148102
rect 381678 148046 399250 148102
rect 399306 148046 399374 148102
rect 399430 148046 399498 148102
rect 399554 148046 399622 148102
rect 399678 148046 417250 148102
rect 417306 148046 417374 148102
rect 417430 148046 417498 148102
rect 417554 148046 417622 148102
rect 417678 148046 435250 148102
rect 435306 148046 435374 148102
rect 435430 148046 435498 148102
rect 435554 148046 435622 148102
rect 435678 148046 453250 148102
rect 453306 148046 453374 148102
rect 453430 148046 453498 148102
rect 453554 148046 453622 148102
rect 453678 148046 471250 148102
rect 471306 148046 471374 148102
rect 471430 148046 471498 148102
rect 471554 148046 471622 148102
rect 471678 148046 489250 148102
rect 489306 148046 489374 148102
rect 489430 148046 489498 148102
rect 489554 148046 489622 148102
rect 489678 148046 507250 148102
rect 507306 148046 507374 148102
rect 507430 148046 507498 148102
rect 507554 148046 507622 148102
rect 507678 148046 525250 148102
rect 525306 148046 525374 148102
rect 525430 148046 525498 148102
rect 525554 148046 525622 148102
rect 525678 148046 543250 148102
rect 543306 148046 543374 148102
rect 543430 148046 543498 148102
rect 543554 148046 543622 148102
rect 543678 148046 561250 148102
rect 561306 148046 561374 148102
rect 561430 148046 561498 148102
rect 561554 148046 561622 148102
rect 561678 148046 579250 148102
rect 579306 148046 579374 148102
rect 579430 148046 579498 148102
rect 579554 148046 579622 148102
rect 579678 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 3250 147978
rect 3306 147922 3374 147978
rect 3430 147922 3498 147978
rect 3554 147922 3622 147978
rect 3678 147922 21250 147978
rect 21306 147922 21374 147978
rect 21430 147922 21498 147978
rect 21554 147922 21622 147978
rect 21678 147922 39250 147978
rect 39306 147922 39374 147978
rect 39430 147922 39498 147978
rect 39554 147922 39622 147978
rect 39678 147922 57250 147978
rect 57306 147922 57374 147978
rect 57430 147922 57498 147978
rect 57554 147922 57622 147978
rect 57678 147922 75250 147978
rect 75306 147922 75374 147978
rect 75430 147922 75498 147978
rect 75554 147922 75622 147978
rect 75678 147922 93250 147978
rect 93306 147922 93374 147978
rect 93430 147922 93498 147978
rect 93554 147922 93622 147978
rect 93678 147922 111250 147978
rect 111306 147922 111374 147978
rect 111430 147922 111498 147978
rect 111554 147922 111622 147978
rect 111678 147922 129250 147978
rect 129306 147922 129374 147978
rect 129430 147922 129498 147978
rect 129554 147922 129622 147978
rect 129678 147922 147250 147978
rect 147306 147922 147374 147978
rect 147430 147922 147498 147978
rect 147554 147922 147622 147978
rect 147678 147922 165250 147978
rect 165306 147922 165374 147978
rect 165430 147922 165498 147978
rect 165554 147922 165622 147978
rect 165678 147922 183250 147978
rect 183306 147922 183374 147978
rect 183430 147922 183498 147978
rect 183554 147922 183622 147978
rect 183678 147922 201250 147978
rect 201306 147922 201374 147978
rect 201430 147922 201498 147978
rect 201554 147922 201622 147978
rect 201678 147922 219250 147978
rect 219306 147922 219374 147978
rect 219430 147922 219498 147978
rect 219554 147922 219622 147978
rect 219678 147922 237250 147978
rect 237306 147922 237374 147978
rect 237430 147922 237498 147978
rect 237554 147922 237622 147978
rect 237678 147922 255250 147978
rect 255306 147922 255374 147978
rect 255430 147922 255498 147978
rect 255554 147922 255622 147978
rect 255678 147922 273250 147978
rect 273306 147922 273374 147978
rect 273430 147922 273498 147978
rect 273554 147922 273622 147978
rect 273678 147922 291250 147978
rect 291306 147922 291374 147978
rect 291430 147922 291498 147978
rect 291554 147922 291622 147978
rect 291678 147922 309250 147978
rect 309306 147922 309374 147978
rect 309430 147922 309498 147978
rect 309554 147922 309622 147978
rect 309678 147922 327250 147978
rect 327306 147922 327374 147978
rect 327430 147922 327498 147978
rect 327554 147922 327622 147978
rect 327678 147922 345250 147978
rect 345306 147922 345374 147978
rect 345430 147922 345498 147978
rect 345554 147922 345622 147978
rect 345678 147922 363250 147978
rect 363306 147922 363374 147978
rect 363430 147922 363498 147978
rect 363554 147922 363622 147978
rect 363678 147922 381250 147978
rect 381306 147922 381374 147978
rect 381430 147922 381498 147978
rect 381554 147922 381622 147978
rect 381678 147922 399250 147978
rect 399306 147922 399374 147978
rect 399430 147922 399498 147978
rect 399554 147922 399622 147978
rect 399678 147922 417250 147978
rect 417306 147922 417374 147978
rect 417430 147922 417498 147978
rect 417554 147922 417622 147978
rect 417678 147922 435250 147978
rect 435306 147922 435374 147978
rect 435430 147922 435498 147978
rect 435554 147922 435622 147978
rect 435678 147922 453250 147978
rect 453306 147922 453374 147978
rect 453430 147922 453498 147978
rect 453554 147922 453622 147978
rect 453678 147922 471250 147978
rect 471306 147922 471374 147978
rect 471430 147922 471498 147978
rect 471554 147922 471622 147978
rect 471678 147922 489250 147978
rect 489306 147922 489374 147978
rect 489430 147922 489498 147978
rect 489554 147922 489622 147978
rect 489678 147922 507250 147978
rect 507306 147922 507374 147978
rect 507430 147922 507498 147978
rect 507554 147922 507622 147978
rect 507678 147922 525250 147978
rect 525306 147922 525374 147978
rect 525430 147922 525498 147978
rect 525554 147922 525622 147978
rect 525678 147922 543250 147978
rect 543306 147922 543374 147978
rect 543430 147922 543498 147978
rect 543554 147922 543622 147978
rect 543678 147922 561250 147978
rect 561306 147922 561374 147978
rect 561430 147922 561498 147978
rect 561554 147922 561622 147978
rect 561678 147922 579250 147978
rect 579306 147922 579374 147978
rect 579430 147922 579498 147978
rect 579554 147922 579622 147978
rect 579678 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 6970 136350
rect 7026 136294 7094 136350
rect 7150 136294 7218 136350
rect 7274 136294 7342 136350
rect 7398 136294 24970 136350
rect 25026 136294 25094 136350
rect 25150 136294 25218 136350
rect 25274 136294 25342 136350
rect 25398 136294 42970 136350
rect 43026 136294 43094 136350
rect 43150 136294 43218 136350
rect 43274 136294 43342 136350
rect 43398 136294 60970 136350
rect 61026 136294 61094 136350
rect 61150 136294 61218 136350
rect 61274 136294 61342 136350
rect 61398 136294 78970 136350
rect 79026 136294 79094 136350
rect 79150 136294 79218 136350
rect 79274 136294 79342 136350
rect 79398 136294 96970 136350
rect 97026 136294 97094 136350
rect 97150 136294 97218 136350
rect 97274 136294 97342 136350
rect 97398 136294 114970 136350
rect 115026 136294 115094 136350
rect 115150 136294 115218 136350
rect 115274 136294 115342 136350
rect 115398 136294 132970 136350
rect 133026 136294 133094 136350
rect 133150 136294 133218 136350
rect 133274 136294 133342 136350
rect 133398 136294 150970 136350
rect 151026 136294 151094 136350
rect 151150 136294 151218 136350
rect 151274 136294 151342 136350
rect 151398 136294 168970 136350
rect 169026 136294 169094 136350
rect 169150 136294 169218 136350
rect 169274 136294 169342 136350
rect 169398 136294 186970 136350
rect 187026 136294 187094 136350
rect 187150 136294 187218 136350
rect 187274 136294 187342 136350
rect 187398 136294 204970 136350
rect 205026 136294 205094 136350
rect 205150 136294 205218 136350
rect 205274 136294 205342 136350
rect 205398 136294 222970 136350
rect 223026 136294 223094 136350
rect 223150 136294 223218 136350
rect 223274 136294 223342 136350
rect 223398 136294 240970 136350
rect 241026 136294 241094 136350
rect 241150 136294 241218 136350
rect 241274 136294 241342 136350
rect 241398 136294 258970 136350
rect 259026 136294 259094 136350
rect 259150 136294 259218 136350
rect 259274 136294 259342 136350
rect 259398 136294 276970 136350
rect 277026 136294 277094 136350
rect 277150 136294 277218 136350
rect 277274 136294 277342 136350
rect 277398 136294 294970 136350
rect 295026 136294 295094 136350
rect 295150 136294 295218 136350
rect 295274 136294 295342 136350
rect 295398 136294 312970 136350
rect 313026 136294 313094 136350
rect 313150 136294 313218 136350
rect 313274 136294 313342 136350
rect 313398 136294 330970 136350
rect 331026 136294 331094 136350
rect 331150 136294 331218 136350
rect 331274 136294 331342 136350
rect 331398 136294 348970 136350
rect 349026 136294 349094 136350
rect 349150 136294 349218 136350
rect 349274 136294 349342 136350
rect 349398 136294 366970 136350
rect 367026 136294 367094 136350
rect 367150 136294 367218 136350
rect 367274 136294 367342 136350
rect 367398 136294 384970 136350
rect 385026 136294 385094 136350
rect 385150 136294 385218 136350
rect 385274 136294 385342 136350
rect 385398 136294 402970 136350
rect 403026 136294 403094 136350
rect 403150 136294 403218 136350
rect 403274 136294 403342 136350
rect 403398 136294 420970 136350
rect 421026 136294 421094 136350
rect 421150 136294 421218 136350
rect 421274 136294 421342 136350
rect 421398 136294 438970 136350
rect 439026 136294 439094 136350
rect 439150 136294 439218 136350
rect 439274 136294 439342 136350
rect 439398 136294 456970 136350
rect 457026 136294 457094 136350
rect 457150 136294 457218 136350
rect 457274 136294 457342 136350
rect 457398 136294 474970 136350
rect 475026 136294 475094 136350
rect 475150 136294 475218 136350
rect 475274 136294 475342 136350
rect 475398 136294 492970 136350
rect 493026 136294 493094 136350
rect 493150 136294 493218 136350
rect 493274 136294 493342 136350
rect 493398 136294 510970 136350
rect 511026 136294 511094 136350
rect 511150 136294 511218 136350
rect 511274 136294 511342 136350
rect 511398 136294 528970 136350
rect 529026 136294 529094 136350
rect 529150 136294 529218 136350
rect 529274 136294 529342 136350
rect 529398 136294 546970 136350
rect 547026 136294 547094 136350
rect 547150 136294 547218 136350
rect 547274 136294 547342 136350
rect 547398 136294 564970 136350
rect 565026 136294 565094 136350
rect 565150 136294 565218 136350
rect 565274 136294 565342 136350
rect 565398 136294 582970 136350
rect 583026 136294 583094 136350
rect 583150 136294 583218 136350
rect 583274 136294 583342 136350
rect 583398 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 6970 136226
rect 7026 136170 7094 136226
rect 7150 136170 7218 136226
rect 7274 136170 7342 136226
rect 7398 136170 24970 136226
rect 25026 136170 25094 136226
rect 25150 136170 25218 136226
rect 25274 136170 25342 136226
rect 25398 136170 42970 136226
rect 43026 136170 43094 136226
rect 43150 136170 43218 136226
rect 43274 136170 43342 136226
rect 43398 136170 60970 136226
rect 61026 136170 61094 136226
rect 61150 136170 61218 136226
rect 61274 136170 61342 136226
rect 61398 136170 78970 136226
rect 79026 136170 79094 136226
rect 79150 136170 79218 136226
rect 79274 136170 79342 136226
rect 79398 136170 96970 136226
rect 97026 136170 97094 136226
rect 97150 136170 97218 136226
rect 97274 136170 97342 136226
rect 97398 136170 114970 136226
rect 115026 136170 115094 136226
rect 115150 136170 115218 136226
rect 115274 136170 115342 136226
rect 115398 136170 132970 136226
rect 133026 136170 133094 136226
rect 133150 136170 133218 136226
rect 133274 136170 133342 136226
rect 133398 136170 150970 136226
rect 151026 136170 151094 136226
rect 151150 136170 151218 136226
rect 151274 136170 151342 136226
rect 151398 136170 168970 136226
rect 169026 136170 169094 136226
rect 169150 136170 169218 136226
rect 169274 136170 169342 136226
rect 169398 136170 186970 136226
rect 187026 136170 187094 136226
rect 187150 136170 187218 136226
rect 187274 136170 187342 136226
rect 187398 136170 204970 136226
rect 205026 136170 205094 136226
rect 205150 136170 205218 136226
rect 205274 136170 205342 136226
rect 205398 136170 222970 136226
rect 223026 136170 223094 136226
rect 223150 136170 223218 136226
rect 223274 136170 223342 136226
rect 223398 136170 240970 136226
rect 241026 136170 241094 136226
rect 241150 136170 241218 136226
rect 241274 136170 241342 136226
rect 241398 136170 258970 136226
rect 259026 136170 259094 136226
rect 259150 136170 259218 136226
rect 259274 136170 259342 136226
rect 259398 136170 276970 136226
rect 277026 136170 277094 136226
rect 277150 136170 277218 136226
rect 277274 136170 277342 136226
rect 277398 136170 294970 136226
rect 295026 136170 295094 136226
rect 295150 136170 295218 136226
rect 295274 136170 295342 136226
rect 295398 136170 312970 136226
rect 313026 136170 313094 136226
rect 313150 136170 313218 136226
rect 313274 136170 313342 136226
rect 313398 136170 330970 136226
rect 331026 136170 331094 136226
rect 331150 136170 331218 136226
rect 331274 136170 331342 136226
rect 331398 136170 348970 136226
rect 349026 136170 349094 136226
rect 349150 136170 349218 136226
rect 349274 136170 349342 136226
rect 349398 136170 366970 136226
rect 367026 136170 367094 136226
rect 367150 136170 367218 136226
rect 367274 136170 367342 136226
rect 367398 136170 384970 136226
rect 385026 136170 385094 136226
rect 385150 136170 385218 136226
rect 385274 136170 385342 136226
rect 385398 136170 402970 136226
rect 403026 136170 403094 136226
rect 403150 136170 403218 136226
rect 403274 136170 403342 136226
rect 403398 136170 420970 136226
rect 421026 136170 421094 136226
rect 421150 136170 421218 136226
rect 421274 136170 421342 136226
rect 421398 136170 438970 136226
rect 439026 136170 439094 136226
rect 439150 136170 439218 136226
rect 439274 136170 439342 136226
rect 439398 136170 456970 136226
rect 457026 136170 457094 136226
rect 457150 136170 457218 136226
rect 457274 136170 457342 136226
rect 457398 136170 474970 136226
rect 475026 136170 475094 136226
rect 475150 136170 475218 136226
rect 475274 136170 475342 136226
rect 475398 136170 492970 136226
rect 493026 136170 493094 136226
rect 493150 136170 493218 136226
rect 493274 136170 493342 136226
rect 493398 136170 510970 136226
rect 511026 136170 511094 136226
rect 511150 136170 511218 136226
rect 511274 136170 511342 136226
rect 511398 136170 528970 136226
rect 529026 136170 529094 136226
rect 529150 136170 529218 136226
rect 529274 136170 529342 136226
rect 529398 136170 546970 136226
rect 547026 136170 547094 136226
rect 547150 136170 547218 136226
rect 547274 136170 547342 136226
rect 547398 136170 564970 136226
rect 565026 136170 565094 136226
rect 565150 136170 565218 136226
rect 565274 136170 565342 136226
rect 565398 136170 582970 136226
rect 583026 136170 583094 136226
rect 583150 136170 583218 136226
rect 583274 136170 583342 136226
rect 583398 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 6970 136102
rect 7026 136046 7094 136102
rect 7150 136046 7218 136102
rect 7274 136046 7342 136102
rect 7398 136046 24970 136102
rect 25026 136046 25094 136102
rect 25150 136046 25218 136102
rect 25274 136046 25342 136102
rect 25398 136046 42970 136102
rect 43026 136046 43094 136102
rect 43150 136046 43218 136102
rect 43274 136046 43342 136102
rect 43398 136046 60970 136102
rect 61026 136046 61094 136102
rect 61150 136046 61218 136102
rect 61274 136046 61342 136102
rect 61398 136046 78970 136102
rect 79026 136046 79094 136102
rect 79150 136046 79218 136102
rect 79274 136046 79342 136102
rect 79398 136046 96970 136102
rect 97026 136046 97094 136102
rect 97150 136046 97218 136102
rect 97274 136046 97342 136102
rect 97398 136046 114970 136102
rect 115026 136046 115094 136102
rect 115150 136046 115218 136102
rect 115274 136046 115342 136102
rect 115398 136046 132970 136102
rect 133026 136046 133094 136102
rect 133150 136046 133218 136102
rect 133274 136046 133342 136102
rect 133398 136046 150970 136102
rect 151026 136046 151094 136102
rect 151150 136046 151218 136102
rect 151274 136046 151342 136102
rect 151398 136046 168970 136102
rect 169026 136046 169094 136102
rect 169150 136046 169218 136102
rect 169274 136046 169342 136102
rect 169398 136046 186970 136102
rect 187026 136046 187094 136102
rect 187150 136046 187218 136102
rect 187274 136046 187342 136102
rect 187398 136046 204970 136102
rect 205026 136046 205094 136102
rect 205150 136046 205218 136102
rect 205274 136046 205342 136102
rect 205398 136046 222970 136102
rect 223026 136046 223094 136102
rect 223150 136046 223218 136102
rect 223274 136046 223342 136102
rect 223398 136046 240970 136102
rect 241026 136046 241094 136102
rect 241150 136046 241218 136102
rect 241274 136046 241342 136102
rect 241398 136046 258970 136102
rect 259026 136046 259094 136102
rect 259150 136046 259218 136102
rect 259274 136046 259342 136102
rect 259398 136046 276970 136102
rect 277026 136046 277094 136102
rect 277150 136046 277218 136102
rect 277274 136046 277342 136102
rect 277398 136046 294970 136102
rect 295026 136046 295094 136102
rect 295150 136046 295218 136102
rect 295274 136046 295342 136102
rect 295398 136046 312970 136102
rect 313026 136046 313094 136102
rect 313150 136046 313218 136102
rect 313274 136046 313342 136102
rect 313398 136046 330970 136102
rect 331026 136046 331094 136102
rect 331150 136046 331218 136102
rect 331274 136046 331342 136102
rect 331398 136046 348970 136102
rect 349026 136046 349094 136102
rect 349150 136046 349218 136102
rect 349274 136046 349342 136102
rect 349398 136046 366970 136102
rect 367026 136046 367094 136102
rect 367150 136046 367218 136102
rect 367274 136046 367342 136102
rect 367398 136046 384970 136102
rect 385026 136046 385094 136102
rect 385150 136046 385218 136102
rect 385274 136046 385342 136102
rect 385398 136046 402970 136102
rect 403026 136046 403094 136102
rect 403150 136046 403218 136102
rect 403274 136046 403342 136102
rect 403398 136046 420970 136102
rect 421026 136046 421094 136102
rect 421150 136046 421218 136102
rect 421274 136046 421342 136102
rect 421398 136046 438970 136102
rect 439026 136046 439094 136102
rect 439150 136046 439218 136102
rect 439274 136046 439342 136102
rect 439398 136046 456970 136102
rect 457026 136046 457094 136102
rect 457150 136046 457218 136102
rect 457274 136046 457342 136102
rect 457398 136046 474970 136102
rect 475026 136046 475094 136102
rect 475150 136046 475218 136102
rect 475274 136046 475342 136102
rect 475398 136046 492970 136102
rect 493026 136046 493094 136102
rect 493150 136046 493218 136102
rect 493274 136046 493342 136102
rect 493398 136046 510970 136102
rect 511026 136046 511094 136102
rect 511150 136046 511218 136102
rect 511274 136046 511342 136102
rect 511398 136046 528970 136102
rect 529026 136046 529094 136102
rect 529150 136046 529218 136102
rect 529274 136046 529342 136102
rect 529398 136046 546970 136102
rect 547026 136046 547094 136102
rect 547150 136046 547218 136102
rect 547274 136046 547342 136102
rect 547398 136046 564970 136102
rect 565026 136046 565094 136102
rect 565150 136046 565218 136102
rect 565274 136046 565342 136102
rect 565398 136046 582970 136102
rect 583026 136046 583094 136102
rect 583150 136046 583218 136102
rect 583274 136046 583342 136102
rect 583398 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 6970 135978
rect 7026 135922 7094 135978
rect 7150 135922 7218 135978
rect 7274 135922 7342 135978
rect 7398 135922 24970 135978
rect 25026 135922 25094 135978
rect 25150 135922 25218 135978
rect 25274 135922 25342 135978
rect 25398 135922 42970 135978
rect 43026 135922 43094 135978
rect 43150 135922 43218 135978
rect 43274 135922 43342 135978
rect 43398 135922 60970 135978
rect 61026 135922 61094 135978
rect 61150 135922 61218 135978
rect 61274 135922 61342 135978
rect 61398 135922 78970 135978
rect 79026 135922 79094 135978
rect 79150 135922 79218 135978
rect 79274 135922 79342 135978
rect 79398 135922 96970 135978
rect 97026 135922 97094 135978
rect 97150 135922 97218 135978
rect 97274 135922 97342 135978
rect 97398 135922 114970 135978
rect 115026 135922 115094 135978
rect 115150 135922 115218 135978
rect 115274 135922 115342 135978
rect 115398 135922 132970 135978
rect 133026 135922 133094 135978
rect 133150 135922 133218 135978
rect 133274 135922 133342 135978
rect 133398 135922 150970 135978
rect 151026 135922 151094 135978
rect 151150 135922 151218 135978
rect 151274 135922 151342 135978
rect 151398 135922 168970 135978
rect 169026 135922 169094 135978
rect 169150 135922 169218 135978
rect 169274 135922 169342 135978
rect 169398 135922 186970 135978
rect 187026 135922 187094 135978
rect 187150 135922 187218 135978
rect 187274 135922 187342 135978
rect 187398 135922 204970 135978
rect 205026 135922 205094 135978
rect 205150 135922 205218 135978
rect 205274 135922 205342 135978
rect 205398 135922 222970 135978
rect 223026 135922 223094 135978
rect 223150 135922 223218 135978
rect 223274 135922 223342 135978
rect 223398 135922 240970 135978
rect 241026 135922 241094 135978
rect 241150 135922 241218 135978
rect 241274 135922 241342 135978
rect 241398 135922 258970 135978
rect 259026 135922 259094 135978
rect 259150 135922 259218 135978
rect 259274 135922 259342 135978
rect 259398 135922 276970 135978
rect 277026 135922 277094 135978
rect 277150 135922 277218 135978
rect 277274 135922 277342 135978
rect 277398 135922 294970 135978
rect 295026 135922 295094 135978
rect 295150 135922 295218 135978
rect 295274 135922 295342 135978
rect 295398 135922 312970 135978
rect 313026 135922 313094 135978
rect 313150 135922 313218 135978
rect 313274 135922 313342 135978
rect 313398 135922 330970 135978
rect 331026 135922 331094 135978
rect 331150 135922 331218 135978
rect 331274 135922 331342 135978
rect 331398 135922 348970 135978
rect 349026 135922 349094 135978
rect 349150 135922 349218 135978
rect 349274 135922 349342 135978
rect 349398 135922 366970 135978
rect 367026 135922 367094 135978
rect 367150 135922 367218 135978
rect 367274 135922 367342 135978
rect 367398 135922 384970 135978
rect 385026 135922 385094 135978
rect 385150 135922 385218 135978
rect 385274 135922 385342 135978
rect 385398 135922 402970 135978
rect 403026 135922 403094 135978
rect 403150 135922 403218 135978
rect 403274 135922 403342 135978
rect 403398 135922 420970 135978
rect 421026 135922 421094 135978
rect 421150 135922 421218 135978
rect 421274 135922 421342 135978
rect 421398 135922 438970 135978
rect 439026 135922 439094 135978
rect 439150 135922 439218 135978
rect 439274 135922 439342 135978
rect 439398 135922 456970 135978
rect 457026 135922 457094 135978
rect 457150 135922 457218 135978
rect 457274 135922 457342 135978
rect 457398 135922 474970 135978
rect 475026 135922 475094 135978
rect 475150 135922 475218 135978
rect 475274 135922 475342 135978
rect 475398 135922 492970 135978
rect 493026 135922 493094 135978
rect 493150 135922 493218 135978
rect 493274 135922 493342 135978
rect 493398 135922 510970 135978
rect 511026 135922 511094 135978
rect 511150 135922 511218 135978
rect 511274 135922 511342 135978
rect 511398 135922 528970 135978
rect 529026 135922 529094 135978
rect 529150 135922 529218 135978
rect 529274 135922 529342 135978
rect 529398 135922 546970 135978
rect 547026 135922 547094 135978
rect 547150 135922 547218 135978
rect 547274 135922 547342 135978
rect 547398 135922 564970 135978
rect 565026 135922 565094 135978
rect 565150 135922 565218 135978
rect 565274 135922 565342 135978
rect 565398 135922 582970 135978
rect 583026 135922 583094 135978
rect 583150 135922 583218 135978
rect 583274 135922 583342 135978
rect 583398 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 3250 130350
rect 3306 130294 3374 130350
rect 3430 130294 3498 130350
rect 3554 130294 3622 130350
rect 3678 130294 21250 130350
rect 21306 130294 21374 130350
rect 21430 130294 21498 130350
rect 21554 130294 21622 130350
rect 21678 130294 39250 130350
rect 39306 130294 39374 130350
rect 39430 130294 39498 130350
rect 39554 130294 39622 130350
rect 39678 130294 57250 130350
rect 57306 130294 57374 130350
rect 57430 130294 57498 130350
rect 57554 130294 57622 130350
rect 57678 130294 75250 130350
rect 75306 130294 75374 130350
rect 75430 130294 75498 130350
rect 75554 130294 75622 130350
rect 75678 130294 93250 130350
rect 93306 130294 93374 130350
rect 93430 130294 93498 130350
rect 93554 130294 93622 130350
rect 93678 130294 111250 130350
rect 111306 130294 111374 130350
rect 111430 130294 111498 130350
rect 111554 130294 111622 130350
rect 111678 130294 129250 130350
rect 129306 130294 129374 130350
rect 129430 130294 129498 130350
rect 129554 130294 129622 130350
rect 129678 130294 147250 130350
rect 147306 130294 147374 130350
rect 147430 130294 147498 130350
rect 147554 130294 147622 130350
rect 147678 130294 165250 130350
rect 165306 130294 165374 130350
rect 165430 130294 165498 130350
rect 165554 130294 165622 130350
rect 165678 130294 183250 130350
rect 183306 130294 183374 130350
rect 183430 130294 183498 130350
rect 183554 130294 183622 130350
rect 183678 130294 201250 130350
rect 201306 130294 201374 130350
rect 201430 130294 201498 130350
rect 201554 130294 201622 130350
rect 201678 130294 219250 130350
rect 219306 130294 219374 130350
rect 219430 130294 219498 130350
rect 219554 130294 219622 130350
rect 219678 130294 237250 130350
rect 237306 130294 237374 130350
rect 237430 130294 237498 130350
rect 237554 130294 237622 130350
rect 237678 130294 255250 130350
rect 255306 130294 255374 130350
rect 255430 130294 255498 130350
rect 255554 130294 255622 130350
rect 255678 130294 273250 130350
rect 273306 130294 273374 130350
rect 273430 130294 273498 130350
rect 273554 130294 273622 130350
rect 273678 130294 291250 130350
rect 291306 130294 291374 130350
rect 291430 130294 291498 130350
rect 291554 130294 291622 130350
rect 291678 130294 309250 130350
rect 309306 130294 309374 130350
rect 309430 130294 309498 130350
rect 309554 130294 309622 130350
rect 309678 130294 327250 130350
rect 327306 130294 327374 130350
rect 327430 130294 327498 130350
rect 327554 130294 327622 130350
rect 327678 130294 345250 130350
rect 345306 130294 345374 130350
rect 345430 130294 345498 130350
rect 345554 130294 345622 130350
rect 345678 130294 363250 130350
rect 363306 130294 363374 130350
rect 363430 130294 363498 130350
rect 363554 130294 363622 130350
rect 363678 130294 381250 130350
rect 381306 130294 381374 130350
rect 381430 130294 381498 130350
rect 381554 130294 381622 130350
rect 381678 130294 399250 130350
rect 399306 130294 399374 130350
rect 399430 130294 399498 130350
rect 399554 130294 399622 130350
rect 399678 130294 417250 130350
rect 417306 130294 417374 130350
rect 417430 130294 417498 130350
rect 417554 130294 417622 130350
rect 417678 130294 435250 130350
rect 435306 130294 435374 130350
rect 435430 130294 435498 130350
rect 435554 130294 435622 130350
rect 435678 130294 453250 130350
rect 453306 130294 453374 130350
rect 453430 130294 453498 130350
rect 453554 130294 453622 130350
rect 453678 130294 471250 130350
rect 471306 130294 471374 130350
rect 471430 130294 471498 130350
rect 471554 130294 471622 130350
rect 471678 130294 489250 130350
rect 489306 130294 489374 130350
rect 489430 130294 489498 130350
rect 489554 130294 489622 130350
rect 489678 130294 507250 130350
rect 507306 130294 507374 130350
rect 507430 130294 507498 130350
rect 507554 130294 507622 130350
rect 507678 130294 525250 130350
rect 525306 130294 525374 130350
rect 525430 130294 525498 130350
rect 525554 130294 525622 130350
rect 525678 130294 543250 130350
rect 543306 130294 543374 130350
rect 543430 130294 543498 130350
rect 543554 130294 543622 130350
rect 543678 130294 561250 130350
rect 561306 130294 561374 130350
rect 561430 130294 561498 130350
rect 561554 130294 561622 130350
rect 561678 130294 579250 130350
rect 579306 130294 579374 130350
rect 579430 130294 579498 130350
rect 579554 130294 579622 130350
rect 579678 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 3250 130226
rect 3306 130170 3374 130226
rect 3430 130170 3498 130226
rect 3554 130170 3622 130226
rect 3678 130170 21250 130226
rect 21306 130170 21374 130226
rect 21430 130170 21498 130226
rect 21554 130170 21622 130226
rect 21678 130170 39250 130226
rect 39306 130170 39374 130226
rect 39430 130170 39498 130226
rect 39554 130170 39622 130226
rect 39678 130170 57250 130226
rect 57306 130170 57374 130226
rect 57430 130170 57498 130226
rect 57554 130170 57622 130226
rect 57678 130170 75250 130226
rect 75306 130170 75374 130226
rect 75430 130170 75498 130226
rect 75554 130170 75622 130226
rect 75678 130170 93250 130226
rect 93306 130170 93374 130226
rect 93430 130170 93498 130226
rect 93554 130170 93622 130226
rect 93678 130170 111250 130226
rect 111306 130170 111374 130226
rect 111430 130170 111498 130226
rect 111554 130170 111622 130226
rect 111678 130170 129250 130226
rect 129306 130170 129374 130226
rect 129430 130170 129498 130226
rect 129554 130170 129622 130226
rect 129678 130170 147250 130226
rect 147306 130170 147374 130226
rect 147430 130170 147498 130226
rect 147554 130170 147622 130226
rect 147678 130170 165250 130226
rect 165306 130170 165374 130226
rect 165430 130170 165498 130226
rect 165554 130170 165622 130226
rect 165678 130170 183250 130226
rect 183306 130170 183374 130226
rect 183430 130170 183498 130226
rect 183554 130170 183622 130226
rect 183678 130170 201250 130226
rect 201306 130170 201374 130226
rect 201430 130170 201498 130226
rect 201554 130170 201622 130226
rect 201678 130170 219250 130226
rect 219306 130170 219374 130226
rect 219430 130170 219498 130226
rect 219554 130170 219622 130226
rect 219678 130170 237250 130226
rect 237306 130170 237374 130226
rect 237430 130170 237498 130226
rect 237554 130170 237622 130226
rect 237678 130170 255250 130226
rect 255306 130170 255374 130226
rect 255430 130170 255498 130226
rect 255554 130170 255622 130226
rect 255678 130170 273250 130226
rect 273306 130170 273374 130226
rect 273430 130170 273498 130226
rect 273554 130170 273622 130226
rect 273678 130170 291250 130226
rect 291306 130170 291374 130226
rect 291430 130170 291498 130226
rect 291554 130170 291622 130226
rect 291678 130170 309250 130226
rect 309306 130170 309374 130226
rect 309430 130170 309498 130226
rect 309554 130170 309622 130226
rect 309678 130170 327250 130226
rect 327306 130170 327374 130226
rect 327430 130170 327498 130226
rect 327554 130170 327622 130226
rect 327678 130170 345250 130226
rect 345306 130170 345374 130226
rect 345430 130170 345498 130226
rect 345554 130170 345622 130226
rect 345678 130170 363250 130226
rect 363306 130170 363374 130226
rect 363430 130170 363498 130226
rect 363554 130170 363622 130226
rect 363678 130170 381250 130226
rect 381306 130170 381374 130226
rect 381430 130170 381498 130226
rect 381554 130170 381622 130226
rect 381678 130170 399250 130226
rect 399306 130170 399374 130226
rect 399430 130170 399498 130226
rect 399554 130170 399622 130226
rect 399678 130170 417250 130226
rect 417306 130170 417374 130226
rect 417430 130170 417498 130226
rect 417554 130170 417622 130226
rect 417678 130170 435250 130226
rect 435306 130170 435374 130226
rect 435430 130170 435498 130226
rect 435554 130170 435622 130226
rect 435678 130170 453250 130226
rect 453306 130170 453374 130226
rect 453430 130170 453498 130226
rect 453554 130170 453622 130226
rect 453678 130170 471250 130226
rect 471306 130170 471374 130226
rect 471430 130170 471498 130226
rect 471554 130170 471622 130226
rect 471678 130170 489250 130226
rect 489306 130170 489374 130226
rect 489430 130170 489498 130226
rect 489554 130170 489622 130226
rect 489678 130170 507250 130226
rect 507306 130170 507374 130226
rect 507430 130170 507498 130226
rect 507554 130170 507622 130226
rect 507678 130170 525250 130226
rect 525306 130170 525374 130226
rect 525430 130170 525498 130226
rect 525554 130170 525622 130226
rect 525678 130170 543250 130226
rect 543306 130170 543374 130226
rect 543430 130170 543498 130226
rect 543554 130170 543622 130226
rect 543678 130170 561250 130226
rect 561306 130170 561374 130226
rect 561430 130170 561498 130226
rect 561554 130170 561622 130226
rect 561678 130170 579250 130226
rect 579306 130170 579374 130226
rect 579430 130170 579498 130226
rect 579554 130170 579622 130226
rect 579678 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 3250 130102
rect 3306 130046 3374 130102
rect 3430 130046 3498 130102
rect 3554 130046 3622 130102
rect 3678 130046 21250 130102
rect 21306 130046 21374 130102
rect 21430 130046 21498 130102
rect 21554 130046 21622 130102
rect 21678 130046 39250 130102
rect 39306 130046 39374 130102
rect 39430 130046 39498 130102
rect 39554 130046 39622 130102
rect 39678 130046 57250 130102
rect 57306 130046 57374 130102
rect 57430 130046 57498 130102
rect 57554 130046 57622 130102
rect 57678 130046 75250 130102
rect 75306 130046 75374 130102
rect 75430 130046 75498 130102
rect 75554 130046 75622 130102
rect 75678 130046 93250 130102
rect 93306 130046 93374 130102
rect 93430 130046 93498 130102
rect 93554 130046 93622 130102
rect 93678 130046 111250 130102
rect 111306 130046 111374 130102
rect 111430 130046 111498 130102
rect 111554 130046 111622 130102
rect 111678 130046 129250 130102
rect 129306 130046 129374 130102
rect 129430 130046 129498 130102
rect 129554 130046 129622 130102
rect 129678 130046 147250 130102
rect 147306 130046 147374 130102
rect 147430 130046 147498 130102
rect 147554 130046 147622 130102
rect 147678 130046 165250 130102
rect 165306 130046 165374 130102
rect 165430 130046 165498 130102
rect 165554 130046 165622 130102
rect 165678 130046 183250 130102
rect 183306 130046 183374 130102
rect 183430 130046 183498 130102
rect 183554 130046 183622 130102
rect 183678 130046 201250 130102
rect 201306 130046 201374 130102
rect 201430 130046 201498 130102
rect 201554 130046 201622 130102
rect 201678 130046 219250 130102
rect 219306 130046 219374 130102
rect 219430 130046 219498 130102
rect 219554 130046 219622 130102
rect 219678 130046 237250 130102
rect 237306 130046 237374 130102
rect 237430 130046 237498 130102
rect 237554 130046 237622 130102
rect 237678 130046 255250 130102
rect 255306 130046 255374 130102
rect 255430 130046 255498 130102
rect 255554 130046 255622 130102
rect 255678 130046 273250 130102
rect 273306 130046 273374 130102
rect 273430 130046 273498 130102
rect 273554 130046 273622 130102
rect 273678 130046 291250 130102
rect 291306 130046 291374 130102
rect 291430 130046 291498 130102
rect 291554 130046 291622 130102
rect 291678 130046 309250 130102
rect 309306 130046 309374 130102
rect 309430 130046 309498 130102
rect 309554 130046 309622 130102
rect 309678 130046 327250 130102
rect 327306 130046 327374 130102
rect 327430 130046 327498 130102
rect 327554 130046 327622 130102
rect 327678 130046 345250 130102
rect 345306 130046 345374 130102
rect 345430 130046 345498 130102
rect 345554 130046 345622 130102
rect 345678 130046 363250 130102
rect 363306 130046 363374 130102
rect 363430 130046 363498 130102
rect 363554 130046 363622 130102
rect 363678 130046 381250 130102
rect 381306 130046 381374 130102
rect 381430 130046 381498 130102
rect 381554 130046 381622 130102
rect 381678 130046 399250 130102
rect 399306 130046 399374 130102
rect 399430 130046 399498 130102
rect 399554 130046 399622 130102
rect 399678 130046 417250 130102
rect 417306 130046 417374 130102
rect 417430 130046 417498 130102
rect 417554 130046 417622 130102
rect 417678 130046 435250 130102
rect 435306 130046 435374 130102
rect 435430 130046 435498 130102
rect 435554 130046 435622 130102
rect 435678 130046 453250 130102
rect 453306 130046 453374 130102
rect 453430 130046 453498 130102
rect 453554 130046 453622 130102
rect 453678 130046 471250 130102
rect 471306 130046 471374 130102
rect 471430 130046 471498 130102
rect 471554 130046 471622 130102
rect 471678 130046 489250 130102
rect 489306 130046 489374 130102
rect 489430 130046 489498 130102
rect 489554 130046 489622 130102
rect 489678 130046 507250 130102
rect 507306 130046 507374 130102
rect 507430 130046 507498 130102
rect 507554 130046 507622 130102
rect 507678 130046 525250 130102
rect 525306 130046 525374 130102
rect 525430 130046 525498 130102
rect 525554 130046 525622 130102
rect 525678 130046 543250 130102
rect 543306 130046 543374 130102
rect 543430 130046 543498 130102
rect 543554 130046 543622 130102
rect 543678 130046 561250 130102
rect 561306 130046 561374 130102
rect 561430 130046 561498 130102
rect 561554 130046 561622 130102
rect 561678 130046 579250 130102
rect 579306 130046 579374 130102
rect 579430 130046 579498 130102
rect 579554 130046 579622 130102
rect 579678 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 3250 129978
rect 3306 129922 3374 129978
rect 3430 129922 3498 129978
rect 3554 129922 3622 129978
rect 3678 129922 21250 129978
rect 21306 129922 21374 129978
rect 21430 129922 21498 129978
rect 21554 129922 21622 129978
rect 21678 129922 39250 129978
rect 39306 129922 39374 129978
rect 39430 129922 39498 129978
rect 39554 129922 39622 129978
rect 39678 129922 57250 129978
rect 57306 129922 57374 129978
rect 57430 129922 57498 129978
rect 57554 129922 57622 129978
rect 57678 129922 75250 129978
rect 75306 129922 75374 129978
rect 75430 129922 75498 129978
rect 75554 129922 75622 129978
rect 75678 129922 93250 129978
rect 93306 129922 93374 129978
rect 93430 129922 93498 129978
rect 93554 129922 93622 129978
rect 93678 129922 111250 129978
rect 111306 129922 111374 129978
rect 111430 129922 111498 129978
rect 111554 129922 111622 129978
rect 111678 129922 129250 129978
rect 129306 129922 129374 129978
rect 129430 129922 129498 129978
rect 129554 129922 129622 129978
rect 129678 129922 147250 129978
rect 147306 129922 147374 129978
rect 147430 129922 147498 129978
rect 147554 129922 147622 129978
rect 147678 129922 165250 129978
rect 165306 129922 165374 129978
rect 165430 129922 165498 129978
rect 165554 129922 165622 129978
rect 165678 129922 183250 129978
rect 183306 129922 183374 129978
rect 183430 129922 183498 129978
rect 183554 129922 183622 129978
rect 183678 129922 201250 129978
rect 201306 129922 201374 129978
rect 201430 129922 201498 129978
rect 201554 129922 201622 129978
rect 201678 129922 219250 129978
rect 219306 129922 219374 129978
rect 219430 129922 219498 129978
rect 219554 129922 219622 129978
rect 219678 129922 237250 129978
rect 237306 129922 237374 129978
rect 237430 129922 237498 129978
rect 237554 129922 237622 129978
rect 237678 129922 255250 129978
rect 255306 129922 255374 129978
rect 255430 129922 255498 129978
rect 255554 129922 255622 129978
rect 255678 129922 273250 129978
rect 273306 129922 273374 129978
rect 273430 129922 273498 129978
rect 273554 129922 273622 129978
rect 273678 129922 291250 129978
rect 291306 129922 291374 129978
rect 291430 129922 291498 129978
rect 291554 129922 291622 129978
rect 291678 129922 309250 129978
rect 309306 129922 309374 129978
rect 309430 129922 309498 129978
rect 309554 129922 309622 129978
rect 309678 129922 327250 129978
rect 327306 129922 327374 129978
rect 327430 129922 327498 129978
rect 327554 129922 327622 129978
rect 327678 129922 345250 129978
rect 345306 129922 345374 129978
rect 345430 129922 345498 129978
rect 345554 129922 345622 129978
rect 345678 129922 363250 129978
rect 363306 129922 363374 129978
rect 363430 129922 363498 129978
rect 363554 129922 363622 129978
rect 363678 129922 381250 129978
rect 381306 129922 381374 129978
rect 381430 129922 381498 129978
rect 381554 129922 381622 129978
rect 381678 129922 399250 129978
rect 399306 129922 399374 129978
rect 399430 129922 399498 129978
rect 399554 129922 399622 129978
rect 399678 129922 417250 129978
rect 417306 129922 417374 129978
rect 417430 129922 417498 129978
rect 417554 129922 417622 129978
rect 417678 129922 435250 129978
rect 435306 129922 435374 129978
rect 435430 129922 435498 129978
rect 435554 129922 435622 129978
rect 435678 129922 453250 129978
rect 453306 129922 453374 129978
rect 453430 129922 453498 129978
rect 453554 129922 453622 129978
rect 453678 129922 471250 129978
rect 471306 129922 471374 129978
rect 471430 129922 471498 129978
rect 471554 129922 471622 129978
rect 471678 129922 489250 129978
rect 489306 129922 489374 129978
rect 489430 129922 489498 129978
rect 489554 129922 489622 129978
rect 489678 129922 507250 129978
rect 507306 129922 507374 129978
rect 507430 129922 507498 129978
rect 507554 129922 507622 129978
rect 507678 129922 525250 129978
rect 525306 129922 525374 129978
rect 525430 129922 525498 129978
rect 525554 129922 525622 129978
rect 525678 129922 543250 129978
rect 543306 129922 543374 129978
rect 543430 129922 543498 129978
rect 543554 129922 543622 129978
rect 543678 129922 561250 129978
rect 561306 129922 561374 129978
rect 561430 129922 561498 129978
rect 561554 129922 561622 129978
rect 561678 129922 579250 129978
rect 579306 129922 579374 129978
rect 579430 129922 579498 129978
rect 579554 129922 579622 129978
rect 579678 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 6970 118350
rect 7026 118294 7094 118350
rect 7150 118294 7218 118350
rect 7274 118294 7342 118350
rect 7398 118294 24970 118350
rect 25026 118294 25094 118350
rect 25150 118294 25218 118350
rect 25274 118294 25342 118350
rect 25398 118294 42970 118350
rect 43026 118294 43094 118350
rect 43150 118294 43218 118350
rect 43274 118294 43342 118350
rect 43398 118294 60970 118350
rect 61026 118294 61094 118350
rect 61150 118294 61218 118350
rect 61274 118294 61342 118350
rect 61398 118294 78970 118350
rect 79026 118294 79094 118350
rect 79150 118294 79218 118350
rect 79274 118294 79342 118350
rect 79398 118294 96970 118350
rect 97026 118294 97094 118350
rect 97150 118294 97218 118350
rect 97274 118294 97342 118350
rect 97398 118294 114970 118350
rect 115026 118294 115094 118350
rect 115150 118294 115218 118350
rect 115274 118294 115342 118350
rect 115398 118294 132970 118350
rect 133026 118294 133094 118350
rect 133150 118294 133218 118350
rect 133274 118294 133342 118350
rect 133398 118294 150970 118350
rect 151026 118294 151094 118350
rect 151150 118294 151218 118350
rect 151274 118294 151342 118350
rect 151398 118294 168970 118350
rect 169026 118294 169094 118350
rect 169150 118294 169218 118350
rect 169274 118294 169342 118350
rect 169398 118294 186970 118350
rect 187026 118294 187094 118350
rect 187150 118294 187218 118350
rect 187274 118294 187342 118350
rect 187398 118294 204970 118350
rect 205026 118294 205094 118350
rect 205150 118294 205218 118350
rect 205274 118294 205342 118350
rect 205398 118294 222970 118350
rect 223026 118294 223094 118350
rect 223150 118294 223218 118350
rect 223274 118294 223342 118350
rect 223398 118294 240970 118350
rect 241026 118294 241094 118350
rect 241150 118294 241218 118350
rect 241274 118294 241342 118350
rect 241398 118294 258970 118350
rect 259026 118294 259094 118350
rect 259150 118294 259218 118350
rect 259274 118294 259342 118350
rect 259398 118294 276970 118350
rect 277026 118294 277094 118350
rect 277150 118294 277218 118350
rect 277274 118294 277342 118350
rect 277398 118294 294970 118350
rect 295026 118294 295094 118350
rect 295150 118294 295218 118350
rect 295274 118294 295342 118350
rect 295398 118294 312970 118350
rect 313026 118294 313094 118350
rect 313150 118294 313218 118350
rect 313274 118294 313342 118350
rect 313398 118294 330970 118350
rect 331026 118294 331094 118350
rect 331150 118294 331218 118350
rect 331274 118294 331342 118350
rect 331398 118294 348970 118350
rect 349026 118294 349094 118350
rect 349150 118294 349218 118350
rect 349274 118294 349342 118350
rect 349398 118294 366970 118350
rect 367026 118294 367094 118350
rect 367150 118294 367218 118350
rect 367274 118294 367342 118350
rect 367398 118294 384970 118350
rect 385026 118294 385094 118350
rect 385150 118294 385218 118350
rect 385274 118294 385342 118350
rect 385398 118294 402970 118350
rect 403026 118294 403094 118350
rect 403150 118294 403218 118350
rect 403274 118294 403342 118350
rect 403398 118294 420970 118350
rect 421026 118294 421094 118350
rect 421150 118294 421218 118350
rect 421274 118294 421342 118350
rect 421398 118294 438970 118350
rect 439026 118294 439094 118350
rect 439150 118294 439218 118350
rect 439274 118294 439342 118350
rect 439398 118294 456970 118350
rect 457026 118294 457094 118350
rect 457150 118294 457218 118350
rect 457274 118294 457342 118350
rect 457398 118294 474970 118350
rect 475026 118294 475094 118350
rect 475150 118294 475218 118350
rect 475274 118294 475342 118350
rect 475398 118294 492970 118350
rect 493026 118294 493094 118350
rect 493150 118294 493218 118350
rect 493274 118294 493342 118350
rect 493398 118294 510970 118350
rect 511026 118294 511094 118350
rect 511150 118294 511218 118350
rect 511274 118294 511342 118350
rect 511398 118294 528970 118350
rect 529026 118294 529094 118350
rect 529150 118294 529218 118350
rect 529274 118294 529342 118350
rect 529398 118294 546970 118350
rect 547026 118294 547094 118350
rect 547150 118294 547218 118350
rect 547274 118294 547342 118350
rect 547398 118294 564970 118350
rect 565026 118294 565094 118350
rect 565150 118294 565218 118350
rect 565274 118294 565342 118350
rect 565398 118294 582970 118350
rect 583026 118294 583094 118350
rect 583150 118294 583218 118350
rect 583274 118294 583342 118350
rect 583398 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 6970 118226
rect 7026 118170 7094 118226
rect 7150 118170 7218 118226
rect 7274 118170 7342 118226
rect 7398 118170 24970 118226
rect 25026 118170 25094 118226
rect 25150 118170 25218 118226
rect 25274 118170 25342 118226
rect 25398 118170 42970 118226
rect 43026 118170 43094 118226
rect 43150 118170 43218 118226
rect 43274 118170 43342 118226
rect 43398 118170 60970 118226
rect 61026 118170 61094 118226
rect 61150 118170 61218 118226
rect 61274 118170 61342 118226
rect 61398 118170 78970 118226
rect 79026 118170 79094 118226
rect 79150 118170 79218 118226
rect 79274 118170 79342 118226
rect 79398 118170 96970 118226
rect 97026 118170 97094 118226
rect 97150 118170 97218 118226
rect 97274 118170 97342 118226
rect 97398 118170 114970 118226
rect 115026 118170 115094 118226
rect 115150 118170 115218 118226
rect 115274 118170 115342 118226
rect 115398 118170 132970 118226
rect 133026 118170 133094 118226
rect 133150 118170 133218 118226
rect 133274 118170 133342 118226
rect 133398 118170 150970 118226
rect 151026 118170 151094 118226
rect 151150 118170 151218 118226
rect 151274 118170 151342 118226
rect 151398 118170 168970 118226
rect 169026 118170 169094 118226
rect 169150 118170 169218 118226
rect 169274 118170 169342 118226
rect 169398 118170 186970 118226
rect 187026 118170 187094 118226
rect 187150 118170 187218 118226
rect 187274 118170 187342 118226
rect 187398 118170 204970 118226
rect 205026 118170 205094 118226
rect 205150 118170 205218 118226
rect 205274 118170 205342 118226
rect 205398 118170 222970 118226
rect 223026 118170 223094 118226
rect 223150 118170 223218 118226
rect 223274 118170 223342 118226
rect 223398 118170 240970 118226
rect 241026 118170 241094 118226
rect 241150 118170 241218 118226
rect 241274 118170 241342 118226
rect 241398 118170 258970 118226
rect 259026 118170 259094 118226
rect 259150 118170 259218 118226
rect 259274 118170 259342 118226
rect 259398 118170 276970 118226
rect 277026 118170 277094 118226
rect 277150 118170 277218 118226
rect 277274 118170 277342 118226
rect 277398 118170 294970 118226
rect 295026 118170 295094 118226
rect 295150 118170 295218 118226
rect 295274 118170 295342 118226
rect 295398 118170 312970 118226
rect 313026 118170 313094 118226
rect 313150 118170 313218 118226
rect 313274 118170 313342 118226
rect 313398 118170 330970 118226
rect 331026 118170 331094 118226
rect 331150 118170 331218 118226
rect 331274 118170 331342 118226
rect 331398 118170 348970 118226
rect 349026 118170 349094 118226
rect 349150 118170 349218 118226
rect 349274 118170 349342 118226
rect 349398 118170 366970 118226
rect 367026 118170 367094 118226
rect 367150 118170 367218 118226
rect 367274 118170 367342 118226
rect 367398 118170 384970 118226
rect 385026 118170 385094 118226
rect 385150 118170 385218 118226
rect 385274 118170 385342 118226
rect 385398 118170 402970 118226
rect 403026 118170 403094 118226
rect 403150 118170 403218 118226
rect 403274 118170 403342 118226
rect 403398 118170 420970 118226
rect 421026 118170 421094 118226
rect 421150 118170 421218 118226
rect 421274 118170 421342 118226
rect 421398 118170 438970 118226
rect 439026 118170 439094 118226
rect 439150 118170 439218 118226
rect 439274 118170 439342 118226
rect 439398 118170 456970 118226
rect 457026 118170 457094 118226
rect 457150 118170 457218 118226
rect 457274 118170 457342 118226
rect 457398 118170 474970 118226
rect 475026 118170 475094 118226
rect 475150 118170 475218 118226
rect 475274 118170 475342 118226
rect 475398 118170 492970 118226
rect 493026 118170 493094 118226
rect 493150 118170 493218 118226
rect 493274 118170 493342 118226
rect 493398 118170 510970 118226
rect 511026 118170 511094 118226
rect 511150 118170 511218 118226
rect 511274 118170 511342 118226
rect 511398 118170 528970 118226
rect 529026 118170 529094 118226
rect 529150 118170 529218 118226
rect 529274 118170 529342 118226
rect 529398 118170 546970 118226
rect 547026 118170 547094 118226
rect 547150 118170 547218 118226
rect 547274 118170 547342 118226
rect 547398 118170 564970 118226
rect 565026 118170 565094 118226
rect 565150 118170 565218 118226
rect 565274 118170 565342 118226
rect 565398 118170 582970 118226
rect 583026 118170 583094 118226
rect 583150 118170 583218 118226
rect 583274 118170 583342 118226
rect 583398 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 6970 118102
rect 7026 118046 7094 118102
rect 7150 118046 7218 118102
rect 7274 118046 7342 118102
rect 7398 118046 24970 118102
rect 25026 118046 25094 118102
rect 25150 118046 25218 118102
rect 25274 118046 25342 118102
rect 25398 118046 42970 118102
rect 43026 118046 43094 118102
rect 43150 118046 43218 118102
rect 43274 118046 43342 118102
rect 43398 118046 60970 118102
rect 61026 118046 61094 118102
rect 61150 118046 61218 118102
rect 61274 118046 61342 118102
rect 61398 118046 78970 118102
rect 79026 118046 79094 118102
rect 79150 118046 79218 118102
rect 79274 118046 79342 118102
rect 79398 118046 96970 118102
rect 97026 118046 97094 118102
rect 97150 118046 97218 118102
rect 97274 118046 97342 118102
rect 97398 118046 114970 118102
rect 115026 118046 115094 118102
rect 115150 118046 115218 118102
rect 115274 118046 115342 118102
rect 115398 118046 132970 118102
rect 133026 118046 133094 118102
rect 133150 118046 133218 118102
rect 133274 118046 133342 118102
rect 133398 118046 150970 118102
rect 151026 118046 151094 118102
rect 151150 118046 151218 118102
rect 151274 118046 151342 118102
rect 151398 118046 168970 118102
rect 169026 118046 169094 118102
rect 169150 118046 169218 118102
rect 169274 118046 169342 118102
rect 169398 118046 186970 118102
rect 187026 118046 187094 118102
rect 187150 118046 187218 118102
rect 187274 118046 187342 118102
rect 187398 118046 204970 118102
rect 205026 118046 205094 118102
rect 205150 118046 205218 118102
rect 205274 118046 205342 118102
rect 205398 118046 222970 118102
rect 223026 118046 223094 118102
rect 223150 118046 223218 118102
rect 223274 118046 223342 118102
rect 223398 118046 240970 118102
rect 241026 118046 241094 118102
rect 241150 118046 241218 118102
rect 241274 118046 241342 118102
rect 241398 118046 258970 118102
rect 259026 118046 259094 118102
rect 259150 118046 259218 118102
rect 259274 118046 259342 118102
rect 259398 118046 276970 118102
rect 277026 118046 277094 118102
rect 277150 118046 277218 118102
rect 277274 118046 277342 118102
rect 277398 118046 294970 118102
rect 295026 118046 295094 118102
rect 295150 118046 295218 118102
rect 295274 118046 295342 118102
rect 295398 118046 312970 118102
rect 313026 118046 313094 118102
rect 313150 118046 313218 118102
rect 313274 118046 313342 118102
rect 313398 118046 330970 118102
rect 331026 118046 331094 118102
rect 331150 118046 331218 118102
rect 331274 118046 331342 118102
rect 331398 118046 348970 118102
rect 349026 118046 349094 118102
rect 349150 118046 349218 118102
rect 349274 118046 349342 118102
rect 349398 118046 366970 118102
rect 367026 118046 367094 118102
rect 367150 118046 367218 118102
rect 367274 118046 367342 118102
rect 367398 118046 384970 118102
rect 385026 118046 385094 118102
rect 385150 118046 385218 118102
rect 385274 118046 385342 118102
rect 385398 118046 402970 118102
rect 403026 118046 403094 118102
rect 403150 118046 403218 118102
rect 403274 118046 403342 118102
rect 403398 118046 420970 118102
rect 421026 118046 421094 118102
rect 421150 118046 421218 118102
rect 421274 118046 421342 118102
rect 421398 118046 438970 118102
rect 439026 118046 439094 118102
rect 439150 118046 439218 118102
rect 439274 118046 439342 118102
rect 439398 118046 456970 118102
rect 457026 118046 457094 118102
rect 457150 118046 457218 118102
rect 457274 118046 457342 118102
rect 457398 118046 474970 118102
rect 475026 118046 475094 118102
rect 475150 118046 475218 118102
rect 475274 118046 475342 118102
rect 475398 118046 492970 118102
rect 493026 118046 493094 118102
rect 493150 118046 493218 118102
rect 493274 118046 493342 118102
rect 493398 118046 510970 118102
rect 511026 118046 511094 118102
rect 511150 118046 511218 118102
rect 511274 118046 511342 118102
rect 511398 118046 528970 118102
rect 529026 118046 529094 118102
rect 529150 118046 529218 118102
rect 529274 118046 529342 118102
rect 529398 118046 546970 118102
rect 547026 118046 547094 118102
rect 547150 118046 547218 118102
rect 547274 118046 547342 118102
rect 547398 118046 564970 118102
rect 565026 118046 565094 118102
rect 565150 118046 565218 118102
rect 565274 118046 565342 118102
rect 565398 118046 582970 118102
rect 583026 118046 583094 118102
rect 583150 118046 583218 118102
rect 583274 118046 583342 118102
rect 583398 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 6970 117978
rect 7026 117922 7094 117978
rect 7150 117922 7218 117978
rect 7274 117922 7342 117978
rect 7398 117922 24970 117978
rect 25026 117922 25094 117978
rect 25150 117922 25218 117978
rect 25274 117922 25342 117978
rect 25398 117922 42970 117978
rect 43026 117922 43094 117978
rect 43150 117922 43218 117978
rect 43274 117922 43342 117978
rect 43398 117922 60970 117978
rect 61026 117922 61094 117978
rect 61150 117922 61218 117978
rect 61274 117922 61342 117978
rect 61398 117922 78970 117978
rect 79026 117922 79094 117978
rect 79150 117922 79218 117978
rect 79274 117922 79342 117978
rect 79398 117922 96970 117978
rect 97026 117922 97094 117978
rect 97150 117922 97218 117978
rect 97274 117922 97342 117978
rect 97398 117922 114970 117978
rect 115026 117922 115094 117978
rect 115150 117922 115218 117978
rect 115274 117922 115342 117978
rect 115398 117922 132970 117978
rect 133026 117922 133094 117978
rect 133150 117922 133218 117978
rect 133274 117922 133342 117978
rect 133398 117922 150970 117978
rect 151026 117922 151094 117978
rect 151150 117922 151218 117978
rect 151274 117922 151342 117978
rect 151398 117922 168970 117978
rect 169026 117922 169094 117978
rect 169150 117922 169218 117978
rect 169274 117922 169342 117978
rect 169398 117922 186970 117978
rect 187026 117922 187094 117978
rect 187150 117922 187218 117978
rect 187274 117922 187342 117978
rect 187398 117922 204970 117978
rect 205026 117922 205094 117978
rect 205150 117922 205218 117978
rect 205274 117922 205342 117978
rect 205398 117922 222970 117978
rect 223026 117922 223094 117978
rect 223150 117922 223218 117978
rect 223274 117922 223342 117978
rect 223398 117922 240970 117978
rect 241026 117922 241094 117978
rect 241150 117922 241218 117978
rect 241274 117922 241342 117978
rect 241398 117922 258970 117978
rect 259026 117922 259094 117978
rect 259150 117922 259218 117978
rect 259274 117922 259342 117978
rect 259398 117922 276970 117978
rect 277026 117922 277094 117978
rect 277150 117922 277218 117978
rect 277274 117922 277342 117978
rect 277398 117922 294970 117978
rect 295026 117922 295094 117978
rect 295150 117922 295218 117978
rect 295274 117922 295342 117978
rect 295398 117922 312970 117978
rect 313026 117922 313094 117978
rect 313150 117922 313218 117978
rect 313274 117922 313342 117978
rect 313398 117922 330970 117978
rect 331026 117922 331094 117978
rect 331150 117922 331218 117978
rect 331274 117922 331342 117978
rect 331398 117922 348970 117978
rect 349026 117922 349094 117978
rect 349150 117922 349218 117978
rect 349274 117922 349342 117978
rect 349398 117922 366970 117978
rect 367026 117922 367094 117978
rect 367150 117922 367218 117978
rect 367274 117922 367342 117978
rect 367398 117922 384970 117978
rect 385026 117922 385094 117978
rect 385150 117922 385218 117978
rect 385274 117922 385342 117978
rect 385398 117922 402970 117978
rect 403026 117922 403094 117978
rect 403150 117922 403218 117978
rect 403274 117922 403342 117978
rect 403398 117922 420970 117978
rect 421026 117922 421094 117978
rect 421150 117922 421218 117978
rect 421274 117922 421342 117978
rect 421398 117922 438970 117978
rect 439026 117922 439094 117978
rect 439150 117922 439218 117978
rect 439274 117922 439342 117978
rect 439398 117922 456970 117978
rect 457026 117922 457094 117978
rect 457150 117922 457218 117978
rect 457274 117922 457342 117978
rect 457398 117922 474970 117978
rect 475026 117922 475094 117978
rect 475150 117922 475218 117978
rect 475274 117922 475342 117978
rect 475398 117922 492970 117978
rect 493026 117922 493094 117978
rect 493150 117922 493218 117978
rect 493274 117922 493342 117978
rect 493398 117922 510970 117978
rect 511026 117922 511094 117978
rect 511150 117922 511218 117978
rect 511274 117922 511342 117978
rect 511398 117922 528970 117978
rect 529026 117922 529094 117978
rect 529150 117922 529218 117978
rect 529274 117922 529342 117978
rect 529398 117922 546970 117978
rect 547026 117922 547094 117978
rect 547150 117922 547218 117978
rect 547274 117922 547342 117978
rect 547398 117922 564970 117978
rect 565026 117922 565094 117978
rect 565150 117922 565218 117978
rect 565274 117922 565342 117978
rect 565398 117922 582970 117978
rect 583026 117922 583094 117978
rect 583150 117922 583218 117978
rect 583274 117922 583342 117978
rect 583398 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 3250 112350
rect 3306 112294 3374 112350
rect 3430 112294 3498 112350
rect 3554 112294 3622 112350
rect 3678 112294 21250 112350
rect 21306 112294 21374 112350
rect 21430 112294 21498 112350
rect 21554 112294 21622 112350
rect 21678 112294 39250 112350
rect 39306 112294 39374 112350
rect 39430 112294 39498 112350
rect 39554 112294 39622 112350
rect 39678 112294 57250 112350
rect 57306 112294 57374 112350
rect 57430 112294 57498 112350
rect 57554 112294 57622 112350
rect 57678 112294 75250 112350
rect 75306 112294 75374 112350
rect 75430 112294 75498 112350
rect 75554 112294 75622 112350
rect 75678 112294 93250 112350
rect 93306 112294 93374 112350
rect 93430 112294 93498 112350
rect 93554 112294 93622 112350
rect 93678 112294 111250 112350
rect 111306 112294 111374 112350
rect 111430 112294 111498 112350
rect 111554 112294 111622 112350
rect 111678 112294 129250 112350
rect 129306 112294 129374 112350
rect 129430 112294 129498 112350
rect 129554 112294 129622 112350
rect 129678 112294 147250 112350
rect 147306 112294 147374 112350
rect 147430 112294 147498 112350
rect 147554 112294 147622 112350
rect 147678 112294 165250 112350
rect 165306 112294 165374 112350
rect 165430 112294 165498 112350
rect 165554 112294 165622 112350
rect 165678 112294 183250 112350
rect 183306 112294 183374 112350
rect 183430 112294 183498 112350
rect 183554 112294 183622 112350
rect 183678 112294 201250 112350
rect 201306 112294 201374 112350
rect 201430 112294 201498 112350
rect 201554 112294 201622 112350
rect 201678 112294 219250 112350
rect 219306 112294 219374 112350
rect 219430 112294 219498 112350
rect 219554 112294 219622 112350
rect 219678 112294 237250 112350
rect 237306 112294 237374 112350
rect 237430 112294 237498 112350
rect 237554 112294 237622 112350
rect 237678 112294 255250 112350
rect 255306 112294 255374 112350
rect 255430 112294 255498 112350
rect 255554 112294 255622 112350
rect 255678 112294 273250 112350
rect 273306 112294 273374 112350
rect 273430 112294 273498 112350
rect 273554 112294 273622 112350
rect 273678 112294 291250 112350
rect 291306 112294 291374 112350
rect 291430 112294 291498 112350
rect 291554 112294 291622 112350
rect 291678 112294 309250 112350
rect 309306 112294 309374 112350
rect 309430 112294 309498 112350
rect 309554 112294 309622 112350
rect 309678 112294 327250 112350
rect 327306 112294 327374 112350
rect 327430 112294 327498 112350
rect 327554 112294 327622 112350
rect 327678 112294 345250 112350
rect 345306 112294 345374 112350
rect 345430 112294 345498 112350
rect 345554 112294 345622 112350
rect 345678 112294 363250 112350
rect 363306 112294 363374 112350
rect 363430 112294 363498 112350
rect 363554 112294 363622 112350
rect 363678 112294 381250 112350
rect 381306 112294 381374 112350
rect 381430 112294 381498 112350
rect 381554 112294 381622 112350
rect 381678 112294 399250 112350
rect 399306 112294 399374 112350
rect 399430 112294 399498 112350
rect 399554 112294 399622 112350
rect 399678 112294 417250 112350
rect 417306 112294 417374 112350
rect 417430 112294 417498 112350
rect 417554 112294 417622 112350
rect 417678 112294 435250 112350
rect 435306 112294 435374 112350
rect 435430 112294 435498 112350
rect 435554 112294 435622 112350
rect 435678 112294 453250 112350
rect 453306 112294 453374 112350
rect 453430 112294 453498 112350
rect 453554 112294 453622 112350
rect 453678 112294 471250 112350
rect 471306 112294 471374 112350
rect 471430 112294 471498 112350
rect 471554 112294 471622 112350
rect 471678 112294 489250 112350
rect 489306 112294 489374 112350
rect 489430 112294 489498 112350
rect 489554 112294 489622 112350
rect 489678 112294 507250 112350
rect 507306 112294 507374 112350
rect 507430 112294 507498 112350
rect 507554 112294 507622 112350
rect 507678 112294 525250 112350
rect 525306 112294 525374 112350
rect 525430 112294 525498 112350
rect 525554 112294 525622 112350
rect 525678 112294 543250 112350
rect 543306 112294 543374 112350
rect 543430 112294 543498 112350
rect 543554 112294 543622 112350
rect 543678 112294 561250 112350
rect 561306 112294 561374 112350
rect 561430 112294 561498 112350
rect 561554 112294 561622 112350
rect 561678 112294 579250 112350
rect 579306 112294 579374 112350
rect 579430 112294 579498 112350
rect 579554 112294 579622 112350
rect 579678 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 3250 112226
rect 3306 112170 3374 112226
rect 3430 112170 3498 112226
rect 3554 112170 3622 112226
rect 3678 112170 21250 112226
rect 21306 112170 21374 112226
rect 21430 112170 21498 112226
rect 21554 112170 21622 112226
rect 21678 112170 39250 112226
rect 39306 112170 39374 112226
rect 39430 112170 39498 112226
rect 39554 112170 39622 112226
rect 39678 112170 57250 112226
rect 57306 112170 57374 112226
rect 57430 112170 57498 112226
rect 57554 112170 57622 112226
rect 57678 112170 75250 112226
rect 75306 112170 75374 112226
rect 75430 112170 75498 112226
rect 75554 112170 75622 112226
rect 75678 112170 93250 112226
rect 93306 112170 93374 112226
rect 93430 112170 93498 112226
rect 93554 112170 93622 112226
rect 93678 112170 111250 112226
rect 111306 112170 111374 112226
rect 111430 112170 111498 112226
rect 111554 112170 111622 112226
rect 111678 112170 129250 112226
rect 129306 112170 129374 112226
rect 129430 112170 129498 112226
rect 129554 112170 129622 112226
rect 129678 112170 147250 112226
rect 147306 112170 147374 112226
rect 147430 112170 147498 112226
rect 147554 112170 147622 112226
rect 147678 112170 165250 112226
rect 165306 112170 165374 112226
rect 165430 112170 165498 112226
rect 165554 112170 165622 112226
rect 165678 112170 183250 112226
rect 183306 112170 183374 112226
rect 183430 112170 183498 112226
rect 183554 112170 183622 112226
rect 183678 112170 201250 112226
rect 201306 112170 201374 112226
rect 201430 112170 201498 112226
rect 201554 112170 201622 112226
rect 201678 112170 219250 112226
rect 219306 112170 219374 112226
rect 219430 112170 219498 112226
rect 219554 112170 219622 112226
rect 219678 112170 237250 112226
rect 237306 112170 237374 112226
rect 237430 112170 237498 112226
rect 237554 112170 237622 112226
rect 237678 112170 255250 112226
rect 255306 112170 255374 112226
rect 255430 112170 255498 112226
rect 255554 112170 255622 112226
rect 255678 112170 273250 112226
rect 273306 112170 273374 112226
rect 273430 112170 273498 112226
rect 273554 112170 273622 112226
rect 273678 112170 291250 112226
rect 291306 112170 291374 112226
rect 291430 112170 291498 112226
rect 291554 112170 291622 112226
rect 291678 112170 309250 112226
rect 309306 112170 309374 112226
rect 309430 112170 309498 112226
rect 309554 112170 309622 112226
rect 309678 112170 327250 112226
rect 327306 112170 327374 112226
rect 327430 112170 327498 112226
rect 327554 112170 327622 112226
rect 327678 112170 345250 112226
rect 345306 112170 345374 112226
rect 345430 112170 345498 112226
rect 345554 112170 345622 112226
rect 345678 112170 363250 112226
rect 363306 112170 363374 112226
rect 363430 112170 363498 112226
rect 363554 112170 363622 112226
rect 363678 112170 381250 112226
rect 381306 112170 381374 112226
rect 381430 112170 381498 112226
rect 381554 112170 381622 112226
rect 381678 112170 399250 112226
rect 399306 112170 399374 112226
rect 399430 112170 399498 112226
rect 399554 112170 399622 112226
rect 399678 112170 417250 112226
rect 417306 112170 417374 112226
rect 417430 112170 417498 112226
rect 417554 112170 417622 112226
rect 417678 112170 435250 112226
rect 435306 112170 435374 112226
rect 435430 112170 435498 112226
rect 435554 112170 435622 112226
rect 435678 112170 453250 112226
rect 453306 112170 453374 112226
rect 453430 112170 453498 112226
rect 453554 112170 453622 112226
rect 453678 112170 471250 112226
rect 471306 112170 471374 112226
rect 471430 112170 471498 112226
rect 471554 112170 471622 112226
rect 471678 112170 489250 112226
rect 489306 112170 489374 112226
rect 489430 112170 489498 112226
rect 489554 112170 489622 112226
rect 489678 112170 507250 112226
rect 507306 112170 507374 112226
rect 507430 112170 507498 112226
rect 507554 112170 507622 112226
rect 507678 112170 525250 112226
rect 525306 112170 525374 112226
rect 525430 112170 525498 112226
rect 525554 112170 525622 112226
rect 525678 112170 543250 112226
rect 543306 112170 543374 112226
rect 543430 112170 543498 112226
rect 543554 112170 543622 112226
rect 543678 112170 561250 112226
rect 561306 112170 561374 112226
rect 561430 112170 561498 112226
rect 561554 112170 561622 112226
rect 561678 112170 579250 112226
rect 579306 112170 579374 112226
rect 579430 112170 579498 112226
rect 579554 112170 579622 112226
rect 579678 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 3250 112102
rect 3306 112046 3374 112102
rect 3430 112046 3498 112102
rect 3554 112046 3622 112102
rect 3678 112046 21250 112102
rect 21306 112046 21374 112102
rect 21430 112046 21498 112102
rect 21554 112046 21622 112102
rect 21678 112046 39250 112102
rect 39306 112046 39374 112102
rect 39430 112046 39498 112102
rect 39554 112046 39622 112102
rect 39678 112046 57250 112102
rect 57306 112046 57374 112102
rect 57430 112046 57498 112102
rect 57554 112046 57622 112102
rect 57678 112046 75250 112102
rect 75306 112046 75374 112102
rect 75430 112046 75498 112102
rect 75554 112046 75622 112102
rect 75678 112046 93250 112102
rect 93306 112046 93374 112102
rect 93430 112046 93498 112102
rect 93554 112046 93622 112102
rect 93678 112046 111250 112102
rect 111306 112046 111374 112102
rect 111430 112046 111498 112102
rect 111554 112046 111622 112102
rect 111678 112046 129250 112102
rect 129306 112046 129374 112102
rect 129430 112046 129498 112102
rect 129554 112046 129622 112102
rect 129678 112046 147250 112102
rect 147306 112046 147374 112102
rect 147430 112046 147498 112102
rect 147554 112046 147622 112102
rect 147678 112046 165250 112102
rect 165306 112046 165374 112102
rect 165430 112046 165498 112102
rect 165554 112046 165622 112102
rect 165678 112046 183250 112102
rect 183306 112046 183374 112102
rect 183430 112046 183498 112102
rect 183554 112046 183622 112102
rect 183678 112046 201250 112102
rect 201306 112046 201374 112102
rect 201430 112046 201498 112102
rect 201554 112046 201622 112102
rect 201678 112046 219250 112102
rect 219306 112046 219374 112102
rect 219430 112046 219498 112102
rect 219554 112046 219622 112102
rect 219678 112046 237250 112102
rect 237306 112046 237374 112102
rect 237430 112046 237498 112102
rect 237554 112046 237622 112102
rect 237678 112046 255250 112102
rect 255306 112046 255374 112102
rect 255430 112046 255498 112102
rect 255554 112046 255622 112102
rect 255678 112046 273250 112102
rect 273306 112046 273374 112102
rect 273430 112046 273498 112102
rect 273554 112046 273622 112102
rect 273678 112046 291250 112102
rect 291306 112046 291374 112102
rect 291430 112046 291498 112102
rect 291554 112046 291622 112102
rect 291678 112046 309250 112102
rect 309306 112046 309374 112102
rect 309430 112046 309498 112102
rect 309554 112046 309622 112102
rect 309678 112046 327250 112102
rect 327306 112046 327374 112102
rect 327430 112046 327498 112102
rect 327554 112046 327622 112102
rect 327678 112046 345250 112102
rect 345306 112046 345374 112102
rect 345430 112046 345498 112102
rect 345554 112046 345622 112102
rect 345678 112046 363250 112102
rect 363306 112046 363374 112102
rect 363430 112046 363498 112102
rect 363554 112046 363622 112102
rect 363678 112046 381250 112102
rect 381306 112046 381374 112102
rect 381430 112046 381498 112102
rect 381554 112046 381622 112102
rect 381678 112046 399250 112102
rect 399306 112046 399374 112102
rect 399430 112046 399498 112102
rect 399554 112046 399622 112102
rect 399678 112046 417250 112102
rect 417306 112046 417374 112102
rect 417430 112046 417498 112102
rect 417554 112046 417622 112102
rect 417678 112046 435250 112102
rect 435306 112046 435374 112102
rect 435430 112046 435498 112102
rect 435554 112046 435622 112102
rect 435678 112046 453250 112102
rect 453306 112046 453374 112102
rect 453430 112046 453498 112102
rect 453554 112046 453622 112102
rect 453678 112046 471250 112102
rect 471306 112046 471374 112102
rect 471430 112046 471498 112102
rect 471554 112046 471622 112102
rect 471678 112046 489250 112102
rect 489306 112046 489374 112102
rect 489430 112046 489498 112102
rect 489554 112046 489622 112102
rect 489678 112046 507250 112102
rect 507306 112046 507374 112102
rect 507430 112046 507498 112102
rect 507554 112046 507622 112102
rect 507678 112046 525250 112102
rect 525306 112046 525374 112102
rect 525430 112046 525498 112102
rect 525554 112046 525622 112102
rect 525678 112046 543250 112102
rect 543306 112046 543374 112102
rect 543430 112046 543498 112102
rect 543554 112046 543622 112102
rect 543678 112046 561250 112102
rect 561306 112046 561374 112102
rect 561430 112046 561498 112102
rect 561554 112046 561622 112102
rect 561678 112046 579250 112102
rect 579306 112046 579374 112102
rect 579430 112046 579498 112102
rect 579554 112046 579622 112102
rect 579678 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 3250 111978
rect 3306 111922 3374 111978
rect 3430 111922 3498 111978
rect 3554 111922 3622 111978
rect 3678 111922 21250 111978
rect 21306 111922 21374 111978
rect 21430 111922 21498 111978
rect 21554 111922 21622 111978
rect 21678 111922 39250 111978
rect 39306 111922 39374 111978
rect 39430 111922 39498 111978
rect 39554 111922 39622 111978
rect 39678 111922 57250 111978
rect 57306 111922 57374 111978
rect 57430 111922 57498 111978
rect 57554 111922 57622 111978
rect 57678 111922 75250 111978
rect 75306 111922 75374 111978
rect 75430 111922 75498 111978
rect 75554 111922 75622 111978
rect 75678 111922 93250 111978
rect 93306 111922 93374 111978
rect 93430 111922 93498 111978
rect 93554 111922 93622 111978
rect 93678 111922 111250 111978
rect 111306 111922 111374 111978
rect 111430 111922 111498 111978
rect 111554 111922 111622 111978
rect 111678 111922 129250 111978
rect 129306 111922 129374 111978
rect 129430 111922 129498 111978
rect 129554 111922 129622 111978
rect 129678 111922 147250 111978
rect 147306 111922 147374 111978
rect 147430 111922 147498 111978
rect 147554 111922 147622 111978
rect 147678 111922 165250 111978
rect 165306 111922 165374 111978
rect 165430 111922 165498 111978
rect 165554 111922 165622 111978
rect 165678 111922 183250 111978
rect 183306 111922 183374 111978
rect 183430 111922 183498 111978
rect 183554 111922 183622 111978
rect 183678 111922 201250 111978
rect 201306 111922 201374 111978
rect 201430 111922 201498 111978
rect 201554 111922 201622 111978
rect 201678 111922 219250 111978
rect 219306 111922 219374 111978
rect 219430 111922 219498 111978
rect 219554 111922 219622 111978
rect 219678 111922 237250 111978
rect 237306 111922 237374 111978
rect 237430 111922 237498 111978
rect 237554 111922 237622 111978
rect 237678 111922 255250 111978
rect 255306 111922 255374 111978
rect 255430 111922 255498 111978
rect 255554 111922 255622 111978
rect 255678 111922 273250 111978
rect 273306 111922 273374 111978
rect 273430 111922 273498 111978
rect 273554 111922 273622 111978
rect 273678 111922 291250 111978
rect 291306 111922 291374 111978
rect 291430 111922 291498 111978
rect 291554 111922 291622 111978
rect 291678 111922 309250 111978
rect 309306 111922 309374 111978
rect 309430 111922 309498 111978
rect 309554 111922 309622 111978
rect 309678 111922 327250 111978
rect 327306 111922 327374 111978
rect 327430 111922 327498 111978
rect 327554 111922 327622 111978
rect 327678 111922 345250 111978
rect 345306 111922 345374 111978
rect 345430 111922 345498 111978
rect 345554 111922 345622 111978
rect 345678 111922 363250 111978
rect 363306 111922 363374 111978
rect 363430 111922 363498 111978
rect 363554 111922 363622 111978
rect 363678 111922 381250 111978
rect 381306 111922 381374 111978
rect 381430 111922 381498 111978
rect 381554 111922 381622 111978
rect 381678 111922 399250 111978
rect 399306 111922 399374 111978
rect 399430 111922 399498 111978
rect 399554 111922 399622 111978
rect 399678 111922 417250 111978
rect 417306 111922 417374 111978
rect 417430 111922 417498 111978
rect 417554 111922 417622 111978
rect 417678 111922 435250 111978
rect 435306 111922 435374 111978
rect 435430 111922 435498 111978
rect 435554 111922 435622 111978
rect 435678 111922 453250 111978
rect 453306 111922 453374 111978
rect 453430 111922 453498 111978
rect 453554 111922 453622 111978
rect 453678 111922 471250 111978
rect 471306 111922 471374 111978
rect 471430 111922 471498 111978
rect 471554 111922 471622 111978
rect 471678 111922 489250 111978
rect 489306 111922 489374 111978
rect 489430 111922 489498 111978
rect 489554 111922 489622 111978
rect 489678 111922 507250 111978
rect 507306 111922 507374 111978
rect 507430 111922 507498 111978
rect 507554 111922 507622 111978
rect 507678 111922 525250 111978
rect 525306 111922 525374 111978
rect 525430 111922 525498 111978
rect 525554 111922 525622 111978
rect 525678 111922 543250 111978
rect 543306 111922 543374 111978
rect 543430 111922 543498 111978
rect 543554 111922 543622 111978
rect 543678 111922 561250 111978
rect 561306 111922 561374 111978
rect 561430 111922 561498 111978
rect 561554 111922 561622 111978
rect 561678 111922 579250 111978
rect 579306 111922 579374 111978
rect 579430 111922 579498 111978
rect 579554 111922 579622 111978
rect 579678 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 6970 100350
rect 7026 100294 7094 100350
rect 7150 100294 7218 100350
rect 7274 100294 7342 100350
rect 7398 100294 24970 100350
rect 25026 100294 25094 100350
rect 25150 100294 25218 100350
rect 25274 100294 25342 100350
rect 25398 100294 42970 100350
rect 43026 100294 43094 100350
rect 43150 100294 43218 100350
rect 43274 100294 43342 100350
rect 43398 100294 60970 100350
rect 61026 100294 61094 100350
rect 61150 100294 61218 100350
rect 61274 100294 61342 100350
rect 61398 100294 78970 100350
rect 79026 100294 79094 100350
rect 79150 100294 79218 100350
rect 79274 100294 79342 100350
rect 79398 100294 96970 100350
rect 97026 100294 97094 100350
rect 97150 100294 97218 100350
rect 97274 100294 97342 100350
rect 97398 100294 114970 100350
rect 115026 100294 115094 100350
rect 115150 100294 115218 100350
rect 115274 100294 115342 100350
rect 115398 100294 132970 100350
rect 133026 100294 133094 100350
rect 133150 100294 133218 100350
rect 133274 100294 133342 100350
rect 133398 100294 150970 100350
rect 151026 100294 151094 100350
rect 151150 100294 151218 100350
rect 151274 100294 151342 100350
rect 151398 100294 168970 100350
rect 169026 100294 169094 100350
rect 169150 100294 169218 100350
rect 169274 100294 169342 100350
rect 169398 100294 186970 100350
rect 187026 100294 187094 100350
rect 187150 100294 187218 100350
rect 187274 100294 187342 100350
rect 187398 100294 204970 100350
rect 205026 100294 205094 100350
rect 205150 100294 205218 100350
rect 205274 100294 205342 100350
rect 205398 100294 222970 100350
rect 223026 100294 223094 100350
rect 223150 100294 223218 100350
rect 223274 100294 223342 100350
rect 223398 100294 240970 100350
rect 241026 100294 241094 100350
rect 241150 100294 241218 100350
rect 241274 100294 241342 100350
rect 241398 100294 258970 100350
rect 259026 100294 259094 100350
rect 259150 100294 259218 100350
rect 259274 100294 259342 100350
rect 259398 100294 276970 100350
rect 277026 100294 277094 100350
rect 277150 100294 277218 100350
rect 277274 100294 277342 100350
rect 277398 100294 294970 100350
rect 295026 100294 295094 100350
rect 295150 100294 295218 100350
rect 295274 100294 295342 100350
rect 295398 100294 312970 100350
rect 313026 100294 313094 100350
rect 313150 100294 313218 100350
rect 313274 100294 313342 100350
rect 313398 100294 330970 100350
rect 331026 100294 331094 100350
rect 331150 100294 331218 100350
rect 331274 100294 331342 100350
rect 331398 100294 348970 100350
rect 349026 100294 349094 100350
rect 349150 100294 349218 100350
rect 349274 100294 349342 100350
rect 349398 100294 366970 100350
rect 367026 100294 367094 100350
rect 367150 100294 367218 100350
rect 367274 100294 367342 100350
rect 367398 100294 384970 100350
rect 385026 100294 385094 100350
rect 385150 100294 385218 100350
rect 385274 100294 385342 100350
rect 385398 100294 402970 100350
rect 403026 100294 403094 100350
rect 403150 100294 403218 100350
rect 403274 100294 403342 100350
rect 403398 100294 420970 100350
rect 421026 100294 421094 100350
rect 421150 100294 421218 100350
rect 421274 100294 421342 100350
rect 421398 100294 438970 100350
rect 439026 100294 439094 100350
rect 439150 100294 439218 100350
rect 439274 100294 439342 100350
rect 439398 100294 456970 100350
rect 457026 100294 457094 100350
rect 457150 100294 457218 100350
rect 457274 100294 457342 100350
rect 457398 100294 474970 100350
rect 475026 100294 475094 100350
rect 475150 100294 475218 100350
rect 475274 100294 475342 100350
rect 475398 100294 492970 100350
rect 493026 100294 493094 100350
rect 493150 100294 493218 100350
rect 493274 100294 493342 100350
rect 493398 100294 510970 100350
rect 511026 100294 511094 100350
rect 511150 100294 511218 100350
rect 511274 100294 511342 100350
rect 511398 100294 528970 100350
rect 529026 100294 529094 100350
rect 529150 100294 529218 100350
rect 529274 100294 529342 100350
rect 529398 100294 546970 100350
rect 547026 100294 547094 100350
rect 547150 100294 547218 100350
rect 547274 100294 547342 100350
rect 547398 100294 564970 100350
rect 565026 100294 565094 100350
rect 565150 100294 565218 100350
rect 565274 100294 565342 100350
rect 565398 100294 582970 100350
rect 583026 100294 583094 100350
rect 583150 100294 583218 100350
rect 583274 100294 583342 100350
rect 583398 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 6970 100226
rect 7026 100170 7094 100226
rect 7150 100170 7218 100226
rect 7274 100170 7342 100226
rect 7398 100170 24970 100226
rect 25026 100170 25094 100226
rect 25150 100170 25218 100226
rect 25274 100170 25342 100226
rect 25398 100170 42970 100226
rect 43026 100170 43094 100226
rect 43150 100170 43218 100226
rect 43274 100170 43342 100226
rect 43398 100170 60970 100226
rect 61026 100170 61094 100226
rect 61150 100170 61218 100226
rect 61274 100170 61342 100226
rect 61398 100170 78970 100226
rect 79026 100170 79094 100226
rect 79150 100170 79218 100226
rect 79274 100170 79342 100226
rect 79398 100170 96970 100226
rect 97026 100170 97094 100226
rect 97150 100170 97218 100226
rect 97274 100170 97342 100226
rect 97398 100170 114970 100226
rect 115026 100170 115094 100226
rect 115150 100170 115218 100226
rect 115274 100170 115342 100226
rect 115398 100170 132970 100226
rect 133026 100170 133094 100226
rect 133150 100170 133218 100226
rect 133274 100170 133342 100226
rect 133398 100170 150970 100226
rect 151026 100170 151094 100226
rect 151150 100170 151218 100226
rect 151274 100170 151342 100226
rect 151398 100170 168970 100226
rect 169026 100170 169094 100226
rect 169150 100170 169218 100226
rect 169274 100170 169342 100226
rect 169398 100170 186970 100226
rect 187026 100170 187094 100226
rect 187150 100170 187218 100226
rect 187274 100170 187342 100226
rect 187398 100170 204970 100226
rect 205026 100170 205094 100226
rect 205150 100170 205218 100226
rect 205274 100170 205342 100226
rect 205398 100170 222970 100226
rect 223026 100170 223094 100226
rect 223150 100170 223218 100226
rect 223274 100170 223342 100226
rect 223398 100170 240970 100226
rect 241026 100170 241094 100226
rect 241150 100170 241218 100226
rect 241274 100170 241342 100226
rect 241398 100170 258970 100226
rect 259026 100170 259094 100226
rect 259150 100170 259218 100226
rect 259274 100170 259342 100226
rect 259398 100170 276970 100226
rect 277026 100170 277094 100226
rect 277150 100170 277218 100226
rect 277274 100170 277342 100226
rect 277398 100170 294970 100226
rect 295026 100170 295094 100226
rect 295150 100170 295218 100226
rect 295274 100170 295342 100226
rect 295398 100170 312970 100226
rect 313026 100170 313094 100226
rect 313150 100170 313218 100226
rect 313274 100170 313342 100226
rect 313398 100170 330970 100226
rect 331026 100170 331094 100226
rect 331150 100170 331218 100226
rect 331274 100170 331342 100226
rect 331398 100170 348970 100226
rect 349026 100170 349094 100226
rect 349150 100170 349218 100226
rect 349274 100170 349342 100226
rect 349398 100170 366970 100226
rect 367026 100170 367094 100226
rect 367150 100170 367218 100226
rect 367274 100170 367342 100226
rect 367398 100170 384970 100226
rect 385026 100170 385094 100226
rect 385150 100170 385218 100226
rect 385274 100170 385342 100226
rect 385398 100170 402970 100226
rect 403026 100170 403094 100226
rect 403150 100170 403218 100226
rect 403274 100170 403342 100226
rect 403398 100170 420970 100226
rect 421026 100170 421094 100226
rect 421150 100170 421218 100226
rect 421274 100170 421342 100226
rect 421398 100170 438970 100226
rect 439026 100170 439094 100226
rect 439150 100170 439218 100226
rect 439274 100170 439342 100226
rect 439398 100170 456970 100226
rect 457026 100170 457094 100226
rect 457150 100170 457218 100226
rect 457274 100170 457342 100226
rect 457398 100170 474970 100226
rect 475026 100170 475094 100226
rect 475150 100170 475218 100226
rect 475274 100170 475342 100226
rect 475398 100170 492970 100226
rect 493026 100170 493094 100226
rect 493150 100170 493218 100226
rect 493274 100170 493342 100226
rect 493398 100170 510970 100226
rect 511026 100170 511094 100226
rect 511150 100170 511218 100226
rect 511274 100170 511342 100226
rect 511398 100170 528970 100226
rect 529026 100170 529094 100226
rect 529150 100170 529218 100226
rect 529274 100170 529342 100226
rect 529398 100170 546970 100226
rect 547026 100170 547094 100226
rect 547150 100170 547218 100226
rect 547274 100170 547342 100226
rect 547398 100170 564970 100226
rect 565026 100170 565094 100226
rect 565150 100170 565218 100226
rect 565274 100170 565342 100226
rect 565398 100170 582970 100226
rect 583026 100170 583094 100226
rect 583150 100170 583218 100226
rect 583274 100170 583342 100226
rect 583398 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 6970 100102
rect 7026 100046 7094 100102
rect 7150 100046 7218 100102
rect 7274 100046 7342 100102
rect 7398 100046 24970 100102
rect 25026 100046 25094 100102
rect 25150 100046 25218 100102
rect 25274 100046 25342 100102
rect 25398 100046 42970 100102
rect 43026 100046 43094 100102
rect 43150 100046 43218 100102
rect 43274 100046 43342 100102
rect 43398 100046 60970 100102
rect 61026 100046 61094 100102
rect 61150 100046 61218 100102
rect 61274 100046 61342 100102
rect 61398 100046 78970 100102
rect 79026 100046 79094 100102
rect 79150 100046 79218 100102
rect 79274 100046 79342 100102
rect 79398 100046 96970 100102
rect 97026 100046 97094 100102
rect 97150 100046 97218 100102
rect 97274 100046 97342 100102
rect 97398 100046 114970 100102
rect 115026 100046 115094 100102
rect 115150 100046 115218 100102
rect 115274 100046 115342 100102
rect 115398 100046 132970 100102
rect 133026 100046 133094 100102
rect 133150 100046 133218 100102
rect 133274 100046 133342 100102
rect 133398 100046 150970 100102
rect 151026 100046 151094 100102
rect 151150 100046 151218 100102
rect 151274 100046 151342 100102
rect 151398 100046 168970 100102
rect 169026 100046 169094 100102
rect 169150 100046 169218 100102
rect 169274 100046 169342 100102
rect 169398 100046 186970 100102
rect 187026 100046 187094 100102
rect 187150 100046 187218 100102
rect 187274 100046 187342 100102
rect 187398 100046 204970 100102
rect 205026 100046 205094 100102
rect 205150 100046 205218 100102
rect 205274 100046 205342 100102
rect 205398 100046 222970 100102
rect 223026 100046 223094 100102
rect 223150 100046 223218 100102
rect 223274 100046 223342 100102
rect 223398 100046 240970 100102
rect 241026 100046 241094 100102
rect 241150 100046 241218 100102
rect 241274 100046 241342 100102
rect 241398 100046 258970 100102
rect 259026 100046 259094 100102
rect 259150 100046 259218 100102
rect 259274 100046 259342 100102
rect 259398 100046 276970 100102
rect 277026 100046 277094 100102
rect 277150 100046 277218 100102
rect 277274 100046 277342 100102
rect 277398 100046 294970 100102
rect 295026 100046 295094 100102
rect 295150 100046 295218 100102
rect 295274 100046 295342 100102
rect 295398 100046 312970 100102
rect 313026 100046 313094 100102
rect 313150 100046 313218 100102
rect 313274 100046 313342 100102
rect 313398 100046 330970 100102
rect 331026 100046 331094 100102
rect 331150 100046 331218 100102
rect 331274 100046 331342 100102
rect 331398 100046 348970 100102
rect 349026 100046 349094 100102
rect 349150 100046 349218 100102
rect 349274 100046 349342 100102
rect 349398 100046 366970 100102
rect 367026 100046 367094 100102
rect 367150 100046 367218 100102
rect 367274 100046 367342 100102
rect 367398 100046 384970 100102
rect 385026 100046 385094 100102
rect 385150 100046 385218 100102
rect 385274 100046 385342 100102
rect 385398 100046 402970 100102
rect 403026 100046 403094 100102
rect 403150 100046 403218 100102
rect 403274 100046 403342 100102
rect 403398 100046 420970 100102
rect 421026 100046 421094 100102
rect 421150 100046 421218 100102
rect 421274 100046 421342 100102
rect 421398 100046 438970 100102
rect 439026 100046 439094 100102
rect 439150 100046 439218 100102
rect 439274 100046 439342 100102
rect 439398 100046 456970 100102
rect 457026 100046 457094 100102
rect 457150 100046 457218 100102
rect 457274 100046 457342 100102
rect 457398 100046 474970 100102
rect 475026 100046 475094 100102
rect 475150 100046 475218 100102
rect 475274 100046 475342 100102
rect 475398 100046 492970 100102
rect 493026 100046 493094 100102
rect 493150 100046 493218 100102
rect 493274 100046 493342 100102
rect 493398 100046 510970 100102
rect 511026 100046 511094 100102
rect 511150 100046 511218 100102
rect 511274 100046 511342 100102
rect 511398 100046 528970 100102
rect 529026 100046 529094 100102
rect 529150 100046 529218 100102
rect 529274 100046 529342 100102
rect 529398 100046 546970 100102
rect 547026 100046 547094 100102
rect 547150 100046 547218 100102
rect 547274 100046 547342 100102
rect 547398 100046 564970 100102
rect 565026 100046 565094 100102
rect 565150 100046 565218 100102
rect 565274 100046 565342 100102
rect 565398 100046 582970 100102
rect 583026 100046 583094 100102
rect 583150 100046 583218 100102
rect 583274 100046 583342 100102
rect 583398 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 6970 99978
rect 7026 99922 7094 99978
rect 7150 99922 7218 99978
rect 7274 99922 7342 99978
rect 7398 99922 24970 99978
rect 25026 99922 25094 99978
rect 25150 99922 25218 99978
rect 25274 99922 25342 99978
rect 25398 99922 42970 99978
rect 43026 99922 43094 99978
rect 43150 99922 43218 99978
rect 43274 99922 43342 99978
rect 43398 99922 60970 99978
rect 61026 99922 61094 99978
rect 61150 99922 61218 99978
rect 61274 99922 61342 99978
rect 61398 99922 78970 99978
rect 79026 99922 79094 99978
rect 79150 99922 79218 99978
rect 79274 99922 79342 99978
rect 79398 99922 96970 99978
rect 97026 99922 97094 99978
rect 97150 99922 97218 99978
rect 97274 99922 97342 99978
rect 97398 99922 114970 99978
rect 115026 99922 115094 99978
rect 115150 99922 115218 99978
rect 115274 99922 115342 99978
rect 115398 99922 132970 99978
rect 133026 99922 133094 99978
rect 133150 99922 133218 99978
rect 133274 99922 133342 99978
rect 133398 99922 150970 99978
rect 151026 99922 151094 99978
rect 151150 99922 151218 99978
rect 151274 99922 151342 99978
rect 151398 99922 168970 99978
rect 169026 99922 169094 99978
rect 169150 99922 169218 99978
rect 169274 99922 169342 99978
rect 169398 99922 186970 99978
rect 187026 99922 187094 99978
rect 187150 99922 187218 99978
rect 187274 99922 187342 99978
rect 187398 99922 204970 99978
rect 205026 99922 205094 99978
rect 205150 99922 205218 99978
rect 205274 99922 205342 99978
rect 205398 99922 222970 99978
rect 223026 99922 223094 99978
rect 223150 99922 223218 99978
rect 223274 99922 223342 99978
rect 223398 99922 240970 99978
rect 241026 99922 241094 99978
rect 241150 99922 241218 99978
rect 241274 99922 241342 99978
rect 241398 99922 258970 99978
rect 259026 99922 259094 99978
rect 259150 99922 259218 99978
rect 259274 99922 259342 99978
rect 259398 99922 276970 99978
rect 277026 99922 277094 99978
rect 277150 99922 277218 99978
rect 277274 99922 277342 99978
rect 277398 99922 294970 99978
rect 295026 99922 295094 99978
rect 295150 99922 295218 99978
rect 295274 99922 295342 99978
rect 295398 99922 312970 99978
rect 313026 99922 313094 99978
rect 313150 99922 313218 99978
rect 313274 99922 313342 99978
rect 313398 99922 330970 99978
rect 331026 99922 331094 99978
rect 331150 99922 331218 99978
rect 331274 99922 331342 99978
rect 331398 99922 348970 99978
rect 349026 99922 349094 99978
rect 349150 99922 349218 99978
rect 349274 99922 349342 99978
rect 349398 99922 366970 99978
rect 367026 99922 367094 99978
rect 367150 99922 367218 99978
rect 367274 99922 367342 99978
rect 367398 99922 384970 99978
rect 385026 99922 385094 99978
rect 385150 99922 385218 99978
rect 385274 99922 385342 99978
rect 385398 99922 402970 99978
rect 403026 99922 403094 99978
rect 403150 99922 403218 99978
rect 403274 99922 403342 99978
rect 403398 99922 420970 99978
rect 421026 99922 421094 99978
rect 421150 99922 421218 99978
rect 421274 99922 421342 99978
rect 421398 99922 438970 99978
rect 439026 99922 439094 99978
rect 439150 99922 439218 99978
rect 439274 99922 439342 99978
rect 439398 99922 456970 99978
rect 457026 99922 457094 99978
rect 457150 99922 457218 99978
rect 457274 99922 457342 99978
rect 457398 99922 474970 99978
rect 475026 99922 475094 99978
rect 475150 99922 475218 99978
rect 475274 99922 475342 99978
rect 475398 99922 492970 99978
rect 493026 99922 493094 99978
rect 493150 99922 493218 99978
rect 493274 99922 493342 99978
rect 493398 99922 510970 99978
rect 511026 99922 511094 99978
rect 511150 99922 511218 99978
rect 511274 99922 511342 99978
rect 511398 99922 528970 99978
rect 529026 99922 529094 99978
rect 529150 99922 529218 99978
rect 529274 99922 529342 99978
rect 529398 99922 546970 99978
rect 547026 99922 547094 99978
rect 547150 99922 547218 99978
rect 547274 99922 547342 99978
rect 547398 99922 564970 99978
rect 565026 99922 565094 99978
rect 565150 99922 565218 99978
rect 565274 99922 565342 99978
rect 565398 99922 582970 99978
rect 583026 99922 583094 99978
rect 583150 99922 583218 99978
rect 583274 99922 583342 99978
rect 583398 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 3250 94350
rect 3306 94294 3374 94350
rect 3430 94294 3498 94350
rect 3554 94294 3622 94350
rect 3678 94294 21250 94350
rect 21306 94294 21374 94350
rect 21430 94294 21498 94350
rect 21554 94294 21622 94350
rect 21678 94294 39250 94350
rect 39306 94294 39374 94350
rect 39430 94294 39498 94350
rect 39554 94294 39622 94350
rect 39678 94294 57250 94350
rect 57306 94294 57374 94350
rect 57430 94294 57498 94350
rect 57554 94294 57622 94350
rect 57678 94294 75250 94350
rect 75306 94294 75374 94350
rect 75430 94294 75498 94350
rect 75554 94294 75622 94350
rect 75678 94294 93250 94350
rect 93306 94294 93374 94350
rect 93430 94294 93498 94350
rect 93554 94294 93622 94350
rect 93678 94294 111250 94350
rect 111306 94294 111374 94350
rect 111430 94294 111498 94350
rect 111554 94294 111622 94350
rect 111678 94294 129250 94350
rect 129306 94294 129374 94350
rect 129430 94294 129498 94350
rect 129554 94294 129622 94350
rect 129678 94294 147250 94350
rect 147306 94294 147374 94350
rect 147430 94294 147498 94350
rect 147554 94294 147622 94350
rect 147678 94294 165250 94350
rect 165306 94294 165374 94350
rect 165430 94294 165498 94350
rect 165554 94294 165622 94350
rect 165678 94294 183250 94350
rect 183306 94294 183374 94350
rect 183430 94294 183498 94350
rect 183554 94294 183622 94350
rect 183678 94294 201250 94350
rect 201306 94294 201374 94350
rect 201430 94294 201498 94350
rect 201554 94294 201622 94350
rect 201678 94294 219250 94350
rect 219306 94294 219374 94350
rect 219430 94294 219498 94350
rect 219554 94294 219622 94350
rect 219678 94294 237250 94350
rect 237306 94294 237374 94350
rect 237430 94294 237498 94350
rect 237554 94294 237622 94350
rect 237678 94294 255250 94350
rect 255306 94294 255374 94350
rect 255430 94294 255498 94350
rect 255554 94294 255622 94350
rect 255678 94294 273250 94350
rect 273306 94294 273374 94350
rect 273430 94294 273498 94350
rect 273554 94294 273622 94350
rect 273678 94294 291250 94350
rect 291306 94294 291374 94350
rect 291430 94294 291498 94350
rect 291554 94294 291622 94350
rect 291678 94294 309250 94350
rect 309306 94294 309374 94350
rect 309430 94294 309498 94350
rect 309554 94294 309622 94350
rect 309678 94294 327250 94350
rect 327306 94294 327374 94350
rect 327430 94294 327498 94350
rect 327554 94294 327622 94350
rect 327678 94294 345250 94350
rect 345306 94294 345374 94350
rect 345430 94294 345498 94350
rect 345554 94294 345622 94350
rect 345678 94294 363250 94350
rect 363306 94294 363374 94350
rect 363430 94294 363498 94350
rect 363554 94294 363622 94350
rect 363678 94294 381250 94350
rect 381306 94294 381374 94350
rect 381430 94294 381498 94350
rect 381554 94294 381622 94350
rect 381678 94294 399250 94350
rect 399306 94294 399374 94350
rect 399430 94294 399498 94350
rect 399554 94294 399622 94350
rect 399678 94294 417250 94350
rect 417306 94294 417374 94350
rect 417430 94294 417498 94350
rect 417554 94294 417622 94350
rect 417678 94294 435250 94350
rect 435306 94294 435374 94350
rect 435430 94294 435498 94350
rect 435554 94294 435622 94350
rect 435678 94294 453250 94350
rect 453306 94294 453374 94350
rect 453430 94294 453498 94350
rect 453554 94294 453622 94350
rect 453678 94294 471250 94350
rect 471306 94294 471374 94350
rect 471430 94294 471498 94350
rect 471554 94294 471622 94350
rect 471678 94294 489250 94350
rect 489306 94294 489374 94350
rect 489430 94294 489498 94350
rect 489554 94294 489622 94350
rect 489678 94294 507250 94350
rect 507306 94294 507374 94350
rect 507430 94294 507498 94350
rect 507554 94294 507622 94350
rect 507678 94294 525250 94350
rect 525306 94294 525374 94350
rect 525430 94294 525498 94350
rect 525554 94294 525622 94350
rect 525678 94294 543250 94350
rect 543306 94294 543374 94350
rect 543430 94294 543498 94350
rect 543554 94294 543622 94350
rect 543678 94294 561250 94350
rect 561306 94294 561374 94350
rect 561430 94294 561498 94350
rect 561554 94294 561622 94350
rect 561678 94294 579250 94350
rect 579306 94294 579374 94350
rect 579430 94294 579498 94350
rect 579554 94294 579622 94350
rect 579678 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 3250 94226
rect 3306 94170 3374 94226
rect 3430 94170 3498 94226
rect 3554 94170 3622 94226
rect 3678 94170 21250 94226
rect 21306 94170 21374 94226
rect 21430 94170 21498 94226
rect 21554 94170 21622 94226
rect 21678 94170 39250 94226
rect 39306 94170 39374 94226
rect 39430 94170 39498 94226
rect 39554 94170 39622 94226
rect 39678 94170 57250 94226
rect 57306 94170 57374 94226
rect 57430 94170 57498 94226
rect 57554 94170 57622 94226
rect 57678 94170 75250 94226
rect 75306 94170 75374 94226
rect 75430 94170 75498 94226
rect 75554 94170 75622 94226
rect 75678 94170 93250 94226
rect 93306 94170 93374 94226
rect 93430 94170 93498 94226
rect 93554 94170 93622 94226
rect 93678 94170 111250 94226
rect 111306 94170 111374 94226
rect 111430 94170 111498 94226
rect 111554 94170 111622 94226
rect 111678 94170 129250 94226
rect 129306 94170 129374 94226
rect 129430 94170 129498 94226
rect 129554 94170 129622 94226
rect 129678 94170 147250 94226
rect 147306 94170 147374 94226
rect 147430 94170 147498 94226
rect 147554 94170 147622 94226
rect 147678 94170 165250 94226
rect 165306 94170 165374 94226
rect 165430 94170 165498 94226
rect 165554 94170 165622 94226
rect 165678 94170 183250 94226
rect 183306 94170 183374 94226
rect 183430 94170 183498 94226
rect 183554 94170 183622 94226
rect 183678 94170 201250 94226
rect 201306 94170 201374 94226
rect 201430 94170 201498 94226
rect 201554 94170 201622 94226
rect 201678 94170 219250 94226
rect 219306 94170 219374 94226
rect 219430 94170 219498 94226
rect 219554 94170 219622 94226
rect 219678 94170 237250 94226
rect 237306 94170 237374 94226
rect 237430 94170 237498 94226
rect 237554 94170 237622 94226
rect 237678 94170 255250 94226
rect 255306 94170 255374 94226
rect 255430 94170 255498 94226
rect 255554 94170 255622 94226
rect 255678 94170 273250 94226
rect 273306 94170 273374 94226
rect 273430 94170 273498 94226
rect 273554 94170 273622 94226
rect 273678 94170 291250 94226
rect 291306 94170 291374 94226
rect 291430 94170 291498 94226
rect 291554 94170 291622 94226
rect 291678 94170 309250 94226
rect 309306 94170 309374 94226
rect 309430 94170 309498 94226
rect 309554 94170 309622 94226
rect 309678 94170 327250 94226
rect 327306 94170 327374 94226
rect 327430 94170 327498 94226
rect 327554 94170 327622 94226
rect 327678 94170 345250 94226
rect 345306 94170 345374 94226
rect 345430 94170 345498 94226
rect 345554 94170 345622 94226
rect 345678 94170 363250 94226
rect 363306 94170 363374 94226
rect 363430 94170 363498 94226
rect 363554 94170 363622 94226
rect 363678 94170 381250 94226
rect 381306 94170 381374 94226
rect 381430 94170 381498 94226
rect 381554 94170 381622 94226
rect 381678 94170 399250 94226
rect 399306 94170 399374 94226
rect 399430 94170 399498 94226
rect 399554 94170 399622 94226
rect 399678 94170 417250 94226
rect 417306 94170 417374 94226
rect 417430 94170 417498 94226
rect 417554 94170 417622 94226
rect 417678 94170 435250 94226
rect 435306 94170 435374 94226
rect 435430 94170 435498 94226
rect 435554 94170 435622 94226
rect 435678 94170 453250 94226
rect 453306 94170 453374 94226
rect 453430 94170 453498 94226
rect 453554 94170 453622 94226
rect 453678 94170 471250 94226
rect 471306 94170 471374 94226
rect 471430 94170 471498 94226
rect 471554 94170 471622 94226
rect 471678 94170 489250 94226
rect 489306 94170 489374 94226
rect 489430 94170 489498 94226
rect 489554 94170 489622 94226
rect 489678 94170 507250 94226
rect 507306 94170 507374 94226
rect 507430 94170 507498 94226
rect 507554 94170 507622 94226
rect 507678 94170 525250 94226
rect 525306 94170 525374 94226
rect 525430 94170 525498 94226
rect 525554 94170 525622 94226
rect 525678 94170 543250 94226
rect 543306 94170 543374 94226
rect 543430 94170 543498 94226
rect 543554 94170 543622 94226
rect 543678 94170 561250 94226
rect 561306 94170 561374 94226
rect 561430 94170 561498 94226
rect 561554 94170 561622 94226
rect 561678 94170 579250 94226
rect 579306 94170 579374 94226
rect 579430 94170 579498 94226
rect 579554 94170 579622 94226
rect 579678 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 3250 94102
rect 3306 94046 3374 94102
rect 3430 94046 3498 94102
rect 3554 94046 3622 94102
rect 3678 94046 21250 94102
rect 21306 94046 21374 94102
rect 21430 94046 21498 94102
rect 21554 94046 21622 94102
rect 21678 94046 39250 94102
rect 39306 94046 39374 94102
rect 39430 94046 39498 94102
rect 39554 94046 39622 94102
rect 39678 94046 57250 94102
rect 57306 94046 57374 94102
rect 57430 94046 57498 94102
rect 57554 94046 57622 94102
rect 57678 94046 75250 94102
rect 75306 94046 75374 94102
rect 75430 94046 75498 94102
rect 75554 94046 75622 94102
rect 75678 94046 93250 94102
rect 93306 94046 93374 94102
rect 93430 94046 93498 94102
rect 93554 94046 93622 94102
rect 93678 94046 111250 94102
rect 111306 94046 111374 94102
rect 111430 94046 111498 94102
rect 111554 94046 111622 94102
rect 111678 94046 129250 94102
rect 129306 94046 129374 94102
rect 129430 94046 129498 94102
rect 129554 94046 129622 94102
rect 129678 94046 147250 94102
rect 147306 94046 147374 94102
rect 147430 94046 147498 94102
rect 147554 94046 147622 94102
rect 147678 94046 165250 94102
rect 165306 94046 165374 94102
rect 165430 94046 165498 94102
rect 165554 94046 165622 94102
rect 165678 94046 183250 94102
rect 183306 94046 183374 94102
rect 183430 94046 183498 94102
rect 183554 94046 183622 94102
rect 183678 94046 201250 94102
rect 201306 94046 201374 94102
rect 201430 94046 201498 94102
rect 201554 94046 201622 94102
rect 201678 94046 219250 94102
rect 219306 94046 219374 94102
rect 219430 94046 219498 94102
rect 219554 94046 219622 94102
rect 219678 94046 237250 94102
rect 237306 94046 237374 94102
rect 237430 94046 237498 94102
rect 237554 94046 237622 94102
rect 237678 94046 255250 94102
rect 255306 94046 255374 94102
rect 255430 94046 255498 94102
rect 255554 94046 255622 94102
rect 255678 94046 273250 94102
rect 273306 94046 273374 94102
rect 273430 94046 273498 94102
rect 273554 94046 273622 94102
rect 273678 94046 291250 94102
rect 291306 94046 291374 94102
rect 291430 94046 291498 94102
rect 291554 94046 291622 94102
rect 291678 94046 309250 94102
rect 309306 94046 309374 94102
rect 309430 94046 309498 94102
rect 309554 94046 309622 94102
rect 309678 94046 327250 94102
rect 327306 94046 327374 94102
rect 327430 94046 327498 94102
rect 327554 94046 327622 94102
rect 327678 94046 345250 94102
rect 345306 94046 345374 94102
rect 345430 94046 345498 94102
rect 345554 94046 345622 94102
rect 345678 94046 363250 94102
rect 363306 94046 363374 94102
rect 363430 94046 363498 94102
rect 363554 94046 363622 94102
rect 363678 94046 381250 94102
rect 381306 94046 381374 94102
rect 381430 94046 381498 94102
rect 381554 94046 381622 94102
rect 381678 94046 399250 94102
rect 399306 94046 399374 94102
rect 399430 94046 399498 94102
rect 399554 94046 399622 94102
rect 399678 94046 417250 94102
rect 417306 94046 417374 94102
rect 417430 94046 417498 94102
rect 417554 94046 417622 94102
rect 417678 94046 435250 94102
rect 435306 94046 435374 94102
rect 435430 94046 435498 94102
rect 435554 94046 435622 94102
rect 435678 94046 453250 94102
rect 453306 94046 453374 94102
rect 453430 94046 453498 94102
rect 453554 94046 453622 94102
rect 453678 94046 471250 94102
rect 471306 94046 471374 94102
rect 471430 94046 471498 94102
rect 471554 94046 471622 94102
rect 471678 94046 489250 94102
rect 489306 94046 489374 94102
rect 489430 94046 489498 94102
rect 489554 94046 489622 94102
rect 489678 94046 507250 94102
rect 507306 94046 507374 94102
rect 507430 94046 507498 94102
rect 507554 94046 507622 94102
rect 507678 94046 525250 94102
rect 525306 94046 525374 94102
rect 525430 94046 525498 94102
rect 525554 94046 525622 94102
rect 525678 94046 543250 94102
rect 543306 94046 543374 94102
rect 543430 94046 543498 94102
rect 543554 94046 543622 94102
rect 543678 94046 561250 94102
rect 561306 94046 561374 94102
rect 561430 94046 561498 94102
rect 561554 94046 561622 94102
rect 561678 94046 579250 94102
rect 579306 94046 579374 94102
rect 579430 94046 579498 94102
rect 579554 94046 579622 94102
rect 579678 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 3250 93978
rect 3306 93922 3374 93978
rect 3430 93922 3498 93978
rect 3554 93922 3622 93978
rect 3678 93922 21250 93978
rect 21306 93922 21374 93978
rect 21430 93922 21498 93978
rect 21554 93922 21622 93978
rect 21678 93922 39250 93978
rect 39306 93922 39374 93978
rect 39430 93922 39498 93978
rect 39554 93922 39622 93978
rect 39678 93922 57250 93978
rect 57306 93922 57374 93978
rect 57430 93922 57498 93978
rect 57554 93922 57622 93978
rect 57678 93922 75250 93978
rect 75306 93922 75374 93978
rect 75430 93922 75498 93978
rect 75554 93922 75622 93978
rect 75678 93922 93250 93978
rect 93306 93922 93374 93978
rect 93430 93922 93498 93978
rect 93554 93922 93622 93978
rect 93678 93922 111250 93978
rect 111306 93922 111374 93978
rect 111430 93922 111498 93978
rect 111554 93922 111622 93978
rect 111678 93922 129250 93978
rect 129306 93922 129374 93978
rect 129430 93922 129498 93978
rect 129554 93922 129622 93978
rect 129678 93922 147250 93978
rect 147306 93922 147374 93978
rect 147430 93922 147498 93978
rect 147554 93922 147622 93978
rect 147678 93922 165250 93978
rect 165306 93922 165374 93978
rect 165430 93922 165498 93978
rect 165554 93922 165622 93978
rect 165678 93922 183250 93978
rect 183306 93922 183374 93978
rect 183430 93922 183498 93978
rect 183554 93922 183622 93978
rect 183678 93922 201250 93978
rect 201306 93922 201374 93978
rect 201430 93922 201498 93978
rect 201554 93922 201622 93978
rect 201678 93922 219250 93978
rect 219306 93922 219374 93978
rect 219430 93922 219498 93978
rect 219554 93922 219622 93978
rect 219678 93922 237250 93978
rect 237306 93922 237374 93978
rect 237430 93922 237498 93978
rect 237554 93922 237622 93978
rect 237678 93922 255250 93978
rect 255306 93922 255374 93978
rect 255430 93922 255498 93978
rect 255554 93922 255622 93978
rect 255678 93922 273250 93978
rect 273306 93922 273374 93978
rect 273430 93922 273498 93978
rect 273554 93922 273622 93978
rect 273678 93922 291250 93978
rect 291306 93922 291374 93978
rect 291430 93922 291498 93978
rect 291554 93922 291622 93978
rect 291678 93922 309250 93978
rect 309306 93922 309374 93978
rect 309430 93922 309498 93978
rect 309554 93922 309622 93978
rect 309678 93922 327250 93978
rect 327306 93922 327374 93978
rect 327430 93922 327498 93978
rect 327554 93922 327622 93978
rect 327678 93922 345250 93978
rect 345306 93922 345374 93978
rect 345430 93922 345498 93978
rect 345554 93922 345622 93978
rect 345678 93922 363250 93978
rect 363306 93922 363374 93978
rect 363430 93922 363498 93978
rect 363554 93922 363622 93978
rect 363678 93922 381250 93978
rect 381306 93922 381374 93978
rect 381430 93922 381498 93978
rect 381554 93922 381622 93978
rect 381678 93922 399250 93978
rect 399306 93922 399374 93978
rect 399430 93922 399498 93978
rect 399554 93922 399622 93978
rect 399678 93922 417250 93978
rect 417306 93922 417374 93978
rect 417430 93922 417498 93978
rect 417554 93922 417622 93978
rect 417678 93922 435250 93978
rect 435306 93922 435374 93978
rect 435430 93922 435498 93978
rect 435554 93922 435622 93978
rect 435678 93922 453250 93978
rect 453306 93922 453374 93978
rect 453430 93922 453498 93978
rect 453554 93922 453622 93978
rect 453678 93922 471250 93978
rect 471306 93922 471374 93978
rect 471430 93922 471498 93978
rect 471554 93922 471622 93978
rect 471678 93922 489250 93978
rect 489306 93922 489374 93978
rect 489430 93922 489498 93978
rect 489554 93922 489622 93978
rect 489678 93922 507250 93978
rect 507306 93922 507374 93978
rect 507430 93922 507498 93978
rect 507554 93922 507622 93978
rect 507678 93922 525250 93978
rect 525306 93922 525374 93978
rect 525430 93922 525498 93978
rect 525554 93922 525622 93978
rect 525678 93922 543250 93978
rect 543306 93922 543374 93978
rect 543430 93922 543498 93978
rect 543554 93922 543622 93978
rect 543678 93922 561250 93978
rect 561306 93922 561374 93978
rect 561430 93922 561498 93978
rect 561554 93922 561622 93978
rect 561678 93922 579250 93978
rect 579306 93922 579374 93978
rect 579430 93922 579498 93978
rect 579554 93922 579622 93978
rect 579678 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 6970 82350
rect 7026 82294 7094 82350
rect 7150 82294 7218 82350
rect 7274 82294 7342 82350
rect 7398 82294 24970 82350
rect 25026 82294 25094 82350
rect 25150 82294 25218 82350
rect 25274 82294 25342 82350
rect 25398 82294 42970 82350
rect 43026 82294 43094 82350
rect 43150 82294 43218 82350
rect 43274 82294 43342 82350
rect 43398 82294 60970 82350
rect 61026 82294 61094 82350
rect 61150 82294 61218 82350
rect 61274 82294 61342 82350
rect 61398 82294 78970 82350
rect 79026 82294 79094 82350
rect 79150 82294 79218 82350
rect 79274 82294 79342 82350
rect 79398 82294 96970 82350
rect 97026 82294 97094 82350
rect 97150 82294 97218 82350
rect 97274 82294 97342 82350
rect 97398 82294 114970 82350
rect 115026 82294 115094 82350
rect 115150 82294 115218 82350
rect 115274 82294 115342 82350
rect 115398 82294 132970 82350
rect 133026 82294 133094 82350
rect 133150 82294 133218 82350
rect 133274 82294 133342 82350
rect 133398 82294 150970 82350
rect 151026 82294 151094 82350
rect 151150 82294 151218 82350
rect 151274 82294 151342 82350
rect 151398 82294 168970 82350
rect 169026 82294 169094 82350
rect 169150 82294 169218 82350
rect 169274 82294 169342 82350
rect 169398 82294 186970 82350
rect 187026 82294 187094 82350
rect 187150 82294 187218 82350
rect 187274 82294 187342 82350
rect 187398 82294 204970 82350
rect 205026 82294 205094 82350
rect 205150 82294 205218 82350
rect 205274 82294 205342 82350
rect 205398 82294 222970 82350
rect 223026 82294 223094 82350
rect 223150 82294 223218 82350
rect 223274 82294 223342 82350
rect 223398 82294 240970 82350
rect 241026 82294 241094 82350
rect 241150 82294 241218 82350
rect 241274 82294 241342 82350
rect 241398 82294 258970 82350
rect 259026 82294 259094 82350
rect 259150 82294 259218 82350
rect 259274 82294 259342 82350
rect 259398 82294 276970 82350
rect 277026 82294 277094 82350
rect 277150 82294 277218 82350
rect 277274 82294 277342 82350
rect 277398 82294 294970 82350
rect 295026 82294 295094 82350
rect 295150 82294 295218 82350
rect 295274 82294 295342 82350
rect 295398 82294 312970 82350
rect 313026 82294 313094 82350
rect 313150 82294 313218 82350
rect 313274 82294 313342 82350
rect 313398 82294 330970 82350
rect 331026 82294 331094 82350
rect 331150 82294 331218 82350
rect 331274 82294 331342 82350
rect 331398 82294 348970 82350
rect 349026 82294 349094 82350
rect 349150 82294 349218 82350
rect 349274 82294 349342 82350
rect 349398 82294 366970 82350
rect 367026 82294 367094 82350
rect 367150 82294 367218 82350
rect 367274 82294 367342 82350
rect 367398 82294 384970 82350
rect 385026 82294 385094 82350
rect 385150 82294 385218 82350
rect 385274 82294 385342 82350
rect 385398 82294 402970 82350
rect 403026 82294 403094 82350
rect 403150 82294 403218 82350
rect 403274 82294 403342 82350
rect 403398 82294 420970 82350
rect 421026 82294 421094 82350
rect 421150 82294 421218 82350
rect 421274 82294 421342 82350
rect 421398 82294 438970 82350
rect 439026 82294 439094 82350
rect 439150 82294 439218 82350
rect 439274 82294 439342 82350
rect 439398 82294 456970 82350
rect 457026 82294 457094 82350
rect 457150 82294 457218 82350
rect 457274 82294 457342 82350
rect 457398 82294 474970 82350
rect 475026 82294 475094 82350
rect 475150 82294 475218 82350
rect 475274 82294 475342 82350
rect 475398 82294 492970 82350
rect 493026 82294 493094 82350
rect 493150 82294 493218 82350
rect 493274 82294 493342 82350
rect 493398 82294 510970 82350
rect 511026 82294 511094 82350
rect 511150 82294 511218 82350
rect 511274 82294 511342 82350
rect 511398 82294 528970 82350
rect 529026 82294 529094 82350
rect 529150 82294 529218 82350
rect 529274 82294 529342 82350
rect 529398 82294 546970 82350
rect 547026 82294 547094 82350
rect 547150 82294 547218 82350
rect 547274 82294 547342 82350
rect 547398 82294 564970 82350
rect 565026 82294 565094 82350
rect 565150 82294 565218 82350
rect 565274 82294 565342 82350
rect 565398 82294 582970 82350
rect 583026 82294 583094 82350
rect 583150 82294 583218 82350
rect 583274 82294 583342 82350
rect 583398 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 6970 82226
rect 7026 82170 7094 82226
rect 7150 82170 7218 82226
rect 7274 82170 7342 82226
rect 7398 82170 24970 82226
rect 25026 82170 25094 82226
rect 25150 82170 25218 82226
rect 25274 82170 25342 82226
rect 25398 82170 42970 82226
rect 43026 82170 43094 82226
rect 43150 82170 43218 82226
rect 43274 82170 43342 82226
rect 43398 82170 60970 82226
rect 61026 82170 61094 82226
rect 61150 82170 61218 82226
rect 61274 82170 61342 82226
rect 61398 82170 78970 82226
rect 79026 82170 79094 82226
rect 79150 82170 79218 82226
rect 79274 82170 79342 82226
rect 79398 82170 96970 82226
rect 97026 82170 97094 82226
rect 97150 82170 97218 82226
rect 97274 82170 97342 82226
rect 97398 82170 114970 82226
rect 115026 82170 115094 82226
rect 115150 82170 115218 82226
rect 115274 82170 115342 82226
rect 115398 82170 132970 82226
rect 133026 82170 133094 82226
rect 133150 82170 133218 82226
rect 133274 82170 133342 82226
rect 133398 82170 150970 82226
rect 151026 82170 151094 82226
rect 151150 82170 151218 82226
rect 151274 82170 151342 82226
rect 151398 82170 168970 82226
rect 169026 82170 169094 82226
rect 169150 82170 169218 82226
rect 169274 82170 169342 82226
rect 169398 82170 186970 82226
rect 187026 82170 187094 82226
rect 187150 82170 187218 82226
rect 187274 82170 187342 82226
rect 187398 82170 204970 82226
rect 205026 82170 205094 82226
rect 205150 82170 205218 82226
rect 205274 82170 205342 82226
rect 205398 82170 222970 82226
rect 223026 82170 223094 82226
rect 223150 82170 223218 82226
rect 223274 82170 223342 82226
rect 223398 82170 240970 82226
rect 241026 82170 241094 82226
rect 241150 82170 241218 82226
rect 241274 82170 241342 82226
rect 241398 82170 258970 82226
rect 259026 82170 259094 82226
rect 259150 82170 259218 82226
rect 259274 82170 259342 82226
rect 259398 82170 276970 82226
rect 277026 82170 277094 82226
rect 277150 82170 277218 82226
rect 277274 82170 277342 82226
rect 277398 82170 294970 82226
rect 295026 82170 295094 82226
rect 295150 82170 295218 82226
rect 295274 82170 295342 82226
rect 295398 82170 312970 82226
rect 313026 82170 313094 82226
rect 313150 82170 313218 82226
rect 313274 82170 313342 82226
rect 313398 82170 330970 82226
rect 331026 82170 331094 82226
rect 331150 82170 331218 82226
rect 331274 82170 331342 82226
rect 331398 82170 348970 82226
rect 349026 82170 349094 82226
rect 349150 82170 349218 82226
rect 349274 82170 349342 82226
rect 349398 82170 366970 82226
rect 367026 82170 367094 82226
rect 367150 82170 367218 82226
rect 367274 82170 367342 82226
rect 367398 82170 384970 82226
rect 385026 82170 385094 82226
rect 385150 82170 385218 82226
rect 385274 82170 385342 82226
rect 385398 82170 402970 82226
rect 403026 82170 403094 82226
rect 403150 82170 403218 82226
rect 403274 82170 403342 82226
rect 403398 82170 420970 82226
rect 421026 82170 421094 82226
rect 421150 82170 421218 82226
rect 421274 82170 421342 82226
rect 421398 82170 438970 82226
rect 439026 82170 439094 82226
rect 439150 82170 439218 82226
rect 439274 82170 439342 82226
rect 439398 82170 456970 82226
rect 457026 82170 457094 82226
rect 457150 82170 457218 82226
rect 457274 82170 457342 82226
rect 457398 82170 474970 82226
rect 475026 82170 475094 82226
rect 475150 82170 475218 82226
rect 475274 82170 475342 82226
rect 475398 82170 492970 82226
rect 493026 82170 493094 82226
rect 493150 82170 493218 82226
rect 493274 82170 493342 82226
rect 493398 82170 510970 82226
rect 511026 82170 511094 82226
rect 511150 82170 511218 82226
rect 511274 82170 511342 82226
rect 511398 82170 528970 82226
rect 529026 82170 529094 82226
rect 529150 82170 529218 82226
rect 529274 82170 529342 82226
rect 529398 82170 546970 82226
rect 547026 82170 547094 82226
rect 547150 82170 547218 82226
rect 547274 82170 547342 82226
rect 547398 82170 564970 82226
rect 565026 82170 565094 82226
rect 565150 82170 565218 82226
rect 565274 82170 565342 82226
rect 565398 82170 582970 82226
rect 583026 82170 583094 82226
rect 583150 82170 583218 82226
rect 583274 82170 583342 82226
rect 583398 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 6970 82102
rect 7026 82046 7094 82102
rect 7150 82046 7218 82102
rect 7274 82046 7342 82102
rect 7398 82046 24970 82102
rect 25026 82046 25094 82102
rect 25150 82046 25218 82102
rect 25274 82046 25342 82102
rect 25398 82046 42970 82102
rect 43026 82046 43094 82102
rect 43150 82046 43218 82102
rect 43274 82046 43342 82102
rect 43398 82046 60970 82102
rect 61026 82046 61094 82102
rect 61150 82046 61218 82102
rect 61274 82046 61342 82102
rect 61398 82046 78970 82102
rect 79026 82046 79094 82102
rect 79150 82046 79218 82102
rect 79274 82046 79342 82102
rect 79398 82046 96970 82102
rect 97026 82046 97094 82102
rect 97150 82046 97218 82102
rect 97274 82046 97342 82102
rect 97398 82046 114970 82102
rect 115026 82046 115094 82102
rect 115150 82046 115218 82102
rect 115274 82046 115342 82102
rect 115398 82046 132970 82102
rect 133026 82046 133094 82102
rect 133150 82046 133218 82102
rect 133274 82046 133342 82102
rect 133398 82046 150970 82102
rect 151026 82046 151094 82102
rect 151150 82046 151218 82102
rect 151274 82046 151342 82102
rect 151398 82046 168970 82102
rect 169026 82046 169094 82102
rect 169150 82046 169218 82102
rect 169274 82046 169342 82102
rect 169398 82046 186970 82102
rect 187026 82046 187094 82102
rect 187150 82046 187218 82102
rect 187274 82046 187342 82102
rect 187398 82046 204970 82102
rect 205026 82046 205094 82102
rect 205150 82046 205218 82102
rect 205274 82046 205342 82102
rect 205398 82046 222970 82102
rect 223026 82046 223094 82102
rect 223150 82046 223218 82102
rect 223274 82046 223342 82102
rect 223398 82046 240970 82102
rect 241026 82046 241094 82102
rect 241150 82046 241218 82102
rect 241274 82046 241342 82102
rect 241398 82046 258970 82102
rect 259026 82046 259094 82102
rect 259150 82046 259218 82102
rect 259274 82046 259342 82102
rect 259398 82046 276970 82102
rect 277026 82046 277094 82102
rect 277150 82046 277218 82102
rect 277274 82046 277342 82102
rect 277398 82046 294970 82102
rect 295026 82046 295094 82102
rect 295150 82046 295218 82102
rect 295274 82046 295342 82102
rect 295398 82046 312970 82102
rect 313026 82046 313094 82102
rect 313150 82046 313218 82102
rect 313274 82046 313342 82102
rect 313398 82046 330970 82102
rect 331026 82046 331094 82102
rect 331150 82046 331218 82102
rect 331274 82046 331342 82102
rect 331398 82046 348970 82102
rect 349026 82046 349094 82102
rect 349150 82046 349218 82102
rect 349274 82046 349342 82102
rect 349398 82046 366970 82102
rect 367026 82046 367094 82102
rect 367150 82046 367218 82102
rect 367274 82046 367342 82102
rect 367398 82046 384970 82102
rect 385026 82046 385094 82102
rect 385150 82046 385218 82102
rect 385274 82046 385342 82102
rect 385398 82046 402970 82102
rect 403026 82046 403094 82102
rect 403150 82046 403218 82102
rect 403274 82046 403342 82102
rect 403398 82046 420970 82102
rect 421026 82046 421094 82102
rect 421150 82046 421218 82102
rect 421274 82046 421342 82102
rect 421398 82046 438970 82102
rect 439026 82046 439094 82102
rect 439150 82046 439218 82102
rect 439274 82046 439342 82102
rect 439398 82046 456970 82102
rect 457026 82046 457094 82102
rect 457150 82046 457218 82102
rect 457274 82046 457342 82102
rect 457398 82046 474970 82102
rect 475026 82046 475094 82102
rect 475150 82046 475218 82102
rect 475274 82046 475342 82102
rect 475398 82046 492970 82102
rect 493026 82046 493094 82102
rect 493150 82046 493218 82102
rect 493274 82046 493342 82102
rect 493398 82046 510970 82102
rect 511026 82046 511094 82102
rect 511150 82046 511218 82102
rect 511274 82046 511342 82102
rect 511398 82046 528970 82102
rect 529026 82046 529094 82102
rect 529150 82046 529218 82102
rect 529274 82046 529342 82102
rect 529398 82046 546970 82102
rect 547026 82046 547094 82102
rect 547150 82046 547218 82102
rect 547274 82046 547342 82102
rect 547398 82046 564970 82102
rect 565026 82046 565094 82102
rect 565150 82046 565218 82102
rect 565274 82046 565342 82102
rect 565398 82046 582970 82102
rect 583026 82046 583094 82102
rect 583150 82046 583218 82102
rect 583274 82046 583342 82102
rect 583398 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 6970 81978
rect 7026 81922 7094 81978
rect 7150 81922 7218 81978
rect 7274 81922 7342 81978
rect 7398 81922 24970 81978
rect 25026 81922 25094 81978
rect 25150 81922 25218 81978
rect 25274 81922 25342 81978
rect 25398 81922 42970 81978
rect 43026 81922 43094 81978
rect 43150 81922 43218 81978
rect 43274 81922 43342 81978
rect 43398 81922 60970 81978
rect 61026 81922 61094 81978
rect 61150 81922 61218 81978
rect 61274 81922 61342 81978
rect 61398 81922 78970 81978
rect 79026 81922 79094 81978
rect 79150 81922 79218 81978
rect 79274 81922 79342 81978
rect 79398 81922 96970 81978
rect 97026 81922 97094 81978
rect 97150 81922 97218 81978
rect 97274 81922 97342 81978
rect 97398 81922 114970 81978
rect 115026 81922 115094 81978
rect 115150 81922 115218 81978
rect 115274 81922 115342 81978
rect 115398 81922 132970 81978
rect 133026 81922 133094 81978
rect 133150 81922 133218 81978
rect 133274 81922 133342 81978
rect 133398 81922 150970 81978
rect 151026 81922 151094 81978
rect 151150 81922 151218 81978
rect 151274 81922 151342 81978
rect 151398 81922 168970 81978
rect 169026 81922 169094 81978
rect 169150 81922 169218 81978
rect 169274 81922 169342 81978
rect 169398 81922 186970 81978
rect 187026 81922 187094 81978
rect 187150 81922 187218 81978
rect 187274 81922 187342 81978
rect 187398 81922 204970 81978
rect 205026 81922 205094 81978
rect 205150 81922 205218 81978
rect 205274 81922 205342 81978
rect 205398 81922 222970 81978
rect 223026 81922 223094 81978
rect 223150 81922 223218 81978
rect 223274 81922 223342 81978
rect 223398 81922 240970 81978
rect 241026 81922 241094 81978
rect 241150 81922 241218 81978
rect 241274 81922 241342 81978
rect 241398 81922 258970 81978
rect 259026 81922 259094 81978
rect 259150 81922 259218 81978
rect 259274 81922 259342 81978
rect 259398 81922 276970 81978
rect 277026 81922 277094 81978
rect 277150 81922 277218 81978
rect 277274 81922 277342 81978
rect 277398 81922 294970 81978
rect 295026 81922 295094 81978
rect 295150 81922 295218 81978
rect 295274 81922 295342 81978
rect 295398 81922 312970 81978
rect 313026 81922 313094 81978
rect 313150 81922 313218 81978
rect 313274 81922 313342 81978
rect 313398 81922 330970 81978
rect 331026 81922 331094 81978
rect 331150 81922 331218 81978
rect 331274 81922 331342 81978
rect 331398 81922 348970 81978
rect 349026 81922 349094 81978
rect 349150 81922 349218 81978
rect 349274 81922 349342 81978
rect 349398 81922 366970 81978
rect 367026 81922 367094 81978
rect 367150 81922 367218 81978
rect 367274 81922 367342 81978
rect 367398 81922 384970 81978
rect 385026 81922 385094 81978
rect 385150 81922 385218 81978
rect 385274 81922 385342 81978
rect 385398 81922 402970 81978
rect 403026 81922 403094 81978
rect 403150 81922 403218 81978
rect 403274 81922 403342 81978
rect 403398 81922 420970 81978
rect 421026 81922 421094 81978
rect 421150 81922 421218 81978
rect 421274 81922 421342 81978
rect 421398 81922 438970 81978
rect 439026 81922 439094 81978
rect 439150 81922 439218 81978
rect 439274 81922 439342 81978
rect 439398 81922 456970 81978
rect 457026 81922 457094 81978
rect 457150 81922 457218 81978
rect 457274 81922 457342 81978
rect 457398 81922 474970 81978
rect 475026 81922 475094 81978
rect 475150 81922 475218 81978
rect 475274 81922 475342 81978
rect 475398 81922 492970 81978
rect 493026 81922 493094 81978
rect 493150 81922 493218 81978
rect 493274 81922 493342 81978
rect 493398 81922 510970 81978
rect 511026 81922 511094 81978
rect 511150 81922 511218 81978
rect 511274 81922 511342 81978
rect 511398 81922 528970 81978
rect 529026 81922 529094 81978
rect 529150 81922 529218 81978
rect 529274 81922 529342 81978
rect 529398 81922 546970 81978
rect 547026 81922 547094 81978
rect 547150 81922 547218 81978
rect 547274 81922 547342 81978
rect 547398 81922 564970 81978
rect 565026 81922 565094 81978
rect 565150 81922 565218 81978
rect 565274 81922 565342 81978
rect 565398 81922 582970 81978
rect 583026 81922 583094 81978
rect 583150 81922 583218 81978
rect 583274 81922 583342 81978
rect 583398 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 3250 76350
rect 3306 76294 3374 76350
rect 3430 76294 3498 76350
rect 3554 76294 3622 76350
rect 3678 76294 21250 76350
rect 21306 76294 21374 76350
rect 21430 76294 21498 76350
rect 21554 76294 21622 76350
rect 21678 76294 39250 76350
rect 39306 76294 39374 76350
rect 39430 76294 39498 76350
rect 39554 76294 39622 76350
rect 39678 76294 57250 76350
rect 57306 76294 57374 76350
rect 57430 76294 57498 76350
rect 57554 76294 57622 76350
rect 57678 76294 75250 76350
rect 75306 76294 75374 76350
rect 75430 76294 75498 76350
rect 75554 76294 75622 76350
rect 75678 76294 93250 76350
rect 93306 76294 93374 76350
rect 93430 76294 93498 76350
rect 93554 76294 93622 76350
rect 93678 76294 111250 76350
rect 111306 76294 111374 76350
rect 111430 76294 111498 76350
rect 111554 76294 111622 76350
rect 111678 76294 129250 76350
rect 129306 76294 129374 76350
rect 129430 76294 129498 76350
rect 129554 76294 129622 76350
rect 129678 76294 147250 76350
rect 147306 76294 147374 76350
rect 147430 76294 147498 76350
rect 147554 76294 147622 76350
rect 147678 76294 165250 76350
rect 165306 76294 165374 76350
rect 165430 76294 165498 76350
rect 165554 76294 165622 76350
rect 165678 76294 183250 76350
rect 183306 76294 183374 76350
rect 183430 76294 183498 76350
rect 183554 76294 183622 76350
rect 183678 76294 201250 76350
rect 201306 76294 201374 76350
rect 201430 76294 201498 76350
rect 201554 76294 201622 76350
rect 201678 76294 219250 76350
rect 219306 76294 219374 76350
rect 219430 76294 219498 76350
rect 219554 76294 219622 76350
rect 219678 76294 237250 76350
rect 237306 76294 237374 76350
rect 237430 76294 237498 76350
rect 237554 76294 237622 76350
rect 237678 76294 255250 76350
rect 255306 76294 255374 76350
rect 255430 76294 255498 76350
rect 255554 76294 255622 76350
rect 255678 76294 273250 76350
rect 273306 76294 273374 76350
rect 273430 76294 273498 76350
rect 273554 76294 273622 76350
rect 273678 76294 291250 76350
rect 291306 76294 291374 76350
rect 291430 76294 291498 76350
rect 291554 76294 291622 76350
rect 291678 76294 309250 76350
rect 309306 76294 309374 76350
rect 309430 76294 309498 76350
rect 309554 76294 309622 76350
rect 309678 76294 327250 76350
rect 327306 76294 327374 76350
rect 327430 76294 327498 76350
rect 327554 76294 327622 76350
rect 327678 76294 345250 76350
rect 345306 76294 345374 76350
rect 345430 76294 345498 76350
rect 345554 76294 345622 76350
rect 345678 76294 363250 76350
rect 363306 76294 363374 76350
rect 363430 76294 363498 76350
rect 363554 76294 363622 76350
rect 363678 76294 381250 76350
rect 381306 76294 381374 76350
rect 381430 76294 381498 76350
rect 381554 76294 381622 76350
rect 381678 76294 399250 76350
rect 399306 76294 399374 76350
rect 399430 76294 399498 76350
rect 399554 76294 399622 76350
rect 399678 76294 417250 76350
rect 417306 76294 417374 76350
rect 417430 76294 417498 76350
rect 417554 76294 417622 76350
rect 417678 76294 435250 76350
rect 435306 76294 435374 76350
rect 435430 76294 435498 76350
rect 435554 76294 435622 76350
rect 435678 76294 453250 76350
rect 453306 76294 453374 76350
rect 453430 76294 453498 76350
rect 453554 76294 453622 76350
rect 453678 76294 471250 76350
rect 471306 76294 471374 76350
rect 471430 76294 471498 76350
rect 471554 76294 471622 76350
rect 471678 76294 489250 76350
rect 489306 76294 489374 76350
rect 489430 76294 489498 76350
rect 489554 76294 489622 76350
rect 489678 76294 507250 76350
rect 507306 76294 507374 76350
rect 507430 76294 507498 76350
rect 507554 76294 507622 76350
rect 507678 76294 525250 76350
rect 525306 76294 525374 76350
rect 525430 76294 525498 76350
rect 525554 76294 525622 76350
rect 525678 76294 543250 76350
rect 543306 76294 543374 76350
rect 543430 76294 543498 76350
rect 543554 76294 543622 76350
rect 543678 76294 561250 76350
rect 561306 76294 561374 76350
rect 561430 76294 561498 76350
rect 561554 76294 561622 76350
rect 561678 76294 579250 76350
rect 579306 76294 579374 76350
rect 579430 76294 579498 76350
rect 579554 76294 579622 76350
rect 579678 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 3250 76226
rect 3306 76170 3374 76226
rect 3430 76170 3498 76226
rect 3554 76170 3622 76226
rect 3678 76170 21250 76226
rect 21306 76170 21374 76226
rect 21430 76170 21498 76226
rect 21554 76170 21622 76226
rect 21678 76170 39250 76226
rect 39306 76170 39374 76226
rect 39430 76170 39498 76226
rect 39554 76170 39622 76226
rect 39678 76170 57250 76226
rect 57306 76170 57374 76226
rect 57430 76170 57498 76226
rect 57554 76170 57622 76226
rect 57678 76170 75250 76226
rect 75306 76170 75374 76226
rect 75430 76170 75498 76226
rect 75554 76170 75622 76226
rect 75678 76170 93250 76226
rect 93306 76170 93374 76226
rect 93430 76170 93498 76226
rect 93554 76170 93622 76226
rect 93678 76170 111250 76226
rect 111306 76170 111374 76226
rect 111430 76170 111498 76226
rect 111554 76170 111622 76226
rect 111678 76170 129250 76226
rect 129306 76170 129374 76226
rect 129430 76170 129498 76226
rect 129554 76170 129622 76226
rect 129678 76170 147250 76226
rect 147306 76170 147374 76226
rect 147430 76170 147498 76226
rect 147554 76170 147622 76226
rect 147678 76170 165250 76226
rect 165306 76170 165374 76226
rect 165430 76170 165498 76226
rect 165554 76170 165622 76226
rect 165678 76170 183250 76226
rect 183306 76170 183374 76226
rect 183430 76170 183498 76226
rect 183554 76170 183622 76226
rect 183678 76170 201250 76226
rect 201306 76170 201374 76226
rect 201430 76170 201498 76226
rect 201554 76170 201622 76226
rect 201678 76170 219250 76226
rect 219306 76170 219374 76226
rect 219430 76170 219498 76226
rect 219554 76170 219622 76226
rect 219678 76170 237250 76226
rect 237306 76170 237374 76226
rect 237430 76170 237498 76226
rect 237554 76170 237622 76226
rect 237678 76170 255250 76226
rect 255306 76170 255374 76226
rect 255430 76170 255498 76226
rect 255554 76170 255622 76226
rect 255678 76170 273250 76226
rect 273306 76170 273374 76226
rect 273430 76170 273498 76226
rect 273554 76170 273622 76226
rect 273678 76170 291250 76226
rect 291306 76170 291374 76226
rect 291430 76170 291498 76226
rect 291554 76170 291622 76226
rect 291678 76170 309250 76226
rect 309306 76170 309374 76226
rect 309430 76170 309498 76226
rect 309554 76170 309622 76226
rect 309678 76170 327250 76226
rect 327306 76170 327374 76226
rect 327430 76170 327498 76226
rect 327554 76170 327622 76226
rect 327678 76170 345250 76226
rect 345306 76170 345374 76226
rect 345430 76170 345498 76226
rect 345554 76170 345622 76226
rect 345678 76170 363250 76226
rect 363306 76170 363374 76226
rect 363430 76170 363498 76226
rect 363554 76170 363622 76226
rect 363678 76170 381250 76226
rect 381306 76170 381374 76226
rect 381430 76170 381498 76226
rect 381554 76170 381622 76226
rect 381678 76170 399250 76226
rect 399306 76170 399374 76226
rect 399430 76170 399498 76226
rect 399554 76170 399622 76226
rect 399678 76170 417250 76226
rect 417306 76170 417374 76226
rect 417430 76170 417498 76226
rect 417554 76170 417622 76226
rect 417678 76170 435250 76226
rect 435306 76170 435374 76226
rect 435430 76170 435498 76226
rect 435554 76170 435622 76226
rect 435678 76170 453250 76226
rect 453306 76170 453374 76226
rect 453430 76170 453498 76226
rect 453554 76170 453622 76226
rect 453678 76170 471250 76226
rect 471306 76170 471374 76226
rect 471430 76170 471498 76226
rect 471554 76170 471622 76226
rect 471678 76170 489250 76226
rect 489306 76170 489374 76226
rect 489430 76170 489498 76226
rect 489554 76170 489622 76226
rect 489678 76170 507250 76226
rect 507306 76170 507374 76226
rect 507430 76170 507498 76226
rect 507554 76170 507622 76226
rect 507678 76170 525250 76226
rect 525306 76170 525374 76226
rect 525430 76170 525498 76226
rect 525554 76170 525622 76226
rect 525678 76170 543250 76226
rect 543306 76170 543374 76226
rect 543430 76170 543498 76226
rect 543554 76170 543622 76226
rect 543678 76170 561250 76226
rect 561306 76170 561374 76226
rect 561430 76170 561498 76226
rect 561554 76170 561622 76226
rect 561678 76170 579250 76226
rect 579306 76170 579374 76226
rect 579430 76170 579498 76226
rect 579554 76170 579622 76226
rect 579678 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 3250 76102
rect 3306 76046 3374 76102
rect 3430 76046 3498 76102
rect 3554 76046 3622 76102
rect 3678 76046 21250 76102
rect 21306 76046 21374 76102
rect 21430 76046 21498 76102
rect 21554 76046 21622 76102
rect 21678 76046 39250 76102
rect 39306 76046 39374 76102
rect 39430 76046 39498 76102
rect 39554 76046 39622 76102
rect 39678 76046 57250 76102
rect 57306 76046 57374 76102
rect 57430 76046 57498 76102
rect 57554 76046 57622 76102
rect 57678 76046 75250 76102
rect 75306 76046 75374 76102
rect 75430 76046 75498 76102
rect 75554 76046 75622 76102
rect 75678 76046 93250 76102
rect 93306 76046 93374 76102
rect 93430 76046 93498 76102
rect 93554 76046 93622 76102
rect 93678 76046 111250 76102
rect 111306 76046 111374 76102
rect 111430 76046 111498 76102
rect 111554 76046 111622 76102
rect 111678 76046 129250 76102
rect 129306 76046 129374 76102
rect 129430 76046 129498 76102
rect 129554 76046 129622 76102
rect 129678 76046 147250 76102
rect 147306 76046 147374 76102
rect 147430 76046 147498 76102
rect 147554 76046 147622 76102
rect 147678 76046 165250 76102
rect 165306 76046 165374 76102
rect 165430 76046 165498 76102
rect 165554 76046 165622 76102
rect 165678 76046 183250 76102
rect 183306 76046 183374 76102
rect 183430 76046 183498 76102
rect 183554 76046 183622 76102
rect 183678 76046 201250 76102
rect 201306 76046 201374 76102
rect 201430 76046 201498 76102
rect 201554 76046 201622 76102
rect 201678 76046 219250 76102
rect 219306 76046 219374 76102
rect 219430 76046 219498 76102
rect 219554 76046 219622 76102
rect 219678 76046 237250 76102
rect 237306 76046 237374 76102
rect 237430 76046 237498 76102
rect 237554 76046 237622 76102
rect 237678 76046 255250 76102
rect 255306 76046 255374 76102
rect 255430 76046 255498 76102
rect 255554 76046 255622 76102
rect 255678 76046 273250 76102
rect 273306 76046 273374 76102
rect 273430 76046 273498 76102
rect 273554 76046 273622 76102
rect 273678 76046 291250 76102
rect 291306 76046 291374 76102
rect 291430 76046 291498 76102
rect 291554 76046 291622 76102
rect 291678 76046 309250 76102
rect 309306 76046 309374 76102
rect 309430 76046 309498 76102
rect 309554 76046 309622 76102
rect 309678 76046 327250 76102
rect 327306 76046 327374 76102
rect 327430 76046 327498 76102
rect 327554 76046 327622 76102
rect 327678 76046 345250 76102
rect 345306 76046 345374 76102
rect 345430 76046 345498 76102
rect 345554 76046 345622 76102
rect 345678 76046 363250 76102
rect 363306 76046 363374 76102
rect 363430 76046 363498 76102
rect 363554 76046 363622 76102
rect 363678 76046 381250 76102
rect 381306 76046 381374 76102
rect 381430 76046 381498 76102
rect 381554 76046 381622 76102
rect 381678 76046 399250 76102
rect 399306 76046 399374 76102
rect 399430 76046 399498 76102
rect 399554 76046 399622 76102
rect 399678 76046 417250 76102
rect 417306 76046 417374 76102
rect 417430 76046 417498 76102
rect 417554 76046 417622 76102
rect 417678 76046 435250 76102
rect 435306 76046 435374 76102
rect 435430 76046 435498 76102
rect 435554 76046 435622 76102
rect 435678 76046 453250 76102
rect 453306 76046 453374 76102
rect 453430 76046 453498 76102
rect 453554 76046 453622 76102
rect 453678 76046 471250 76102
rect 471306 76046 471374 76102
rect 471430 76046 471498 76102
rect 471554 76046 471622 76102
rect 471678 76046 489250 76102
rect 489306 76046 489374 76102
rect 489430 76046 489498 76102
rect 489554 76046 489622 76102
rect 489678 76046 507250 76102
rect 507306 76046 507374 76102
rect 507430 76046 507498 76102
rect 507554 76046 507622 76102
rect 507678 76046 525250 76102
rect 525306 76046 525374 76102
rect 525430 76046 525498 76102
rect 525554 76046 525622 76102
rect 525678 76046 543250 76102
rect 543306 76046 543374 76102
rect 543430 76046 543498 76102
rect 543554 76046 543622 76102
rect 543678 76046 561250 76102
rect 561306 76046 561374 76102
rect 561430 76046 561498 76102
rect 561554 76046 561622 76102
rect 561678 76046 579250 76102
rect 579306 76046 579374 76102
rect 579430 76046 579498 76102
rect 579554 76046 579622 76102
rect 579678 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 3250 75978
rect 3306 75922 3374 75978
rect 3430 75922 3498 75978
rect 3554 75922 3622 75978
rect 3678 75922 21250 75978
rect 21306 75922 21374 75978
rect 21430 75922 21498 75978
rect 21554 75922 21622 75978
rect 21678 75922 39250 75978
rect 39306 75922 39374 75978
rect 39430 75922 39498 75978
rect 39554 75922 39622 75978
rect 39678 75922 57250 75978
rect 57306 75922 57374 75978
rect 57430 75922 57498 75978
rect 57554 75922 57622 75978
rect 57678 75922 75250 75978
rect 75306 75922 75374 75978
rect 75430 75922 75498 75978
rect 75554 75922 75622 75978
rect 75678 75922 93250 75978
rect 93306 75922 93374 75978
rect 93430 75922 93498 75978
rect 93554 75922 93622 75978
rect 93678 75922 111250 75978
rect 111306 75922 111374 75978
rect 111430 75922 111498 75978
rect 111554 75922 111622 75978
rect 111678 75922 129250 75978
rect 129306 75922 129374 75978
rect 129430 75922 129498 75978
rect 129554 75922 129622 75978
rect 129678 75922 147250 75978
rect 147306 75922 147374 75978
rect 147430 75922 147498 75978
rect 147554 75922 147622 75978
rect 147678 75922 165250 75978
rect 165306 75922 165374 75978
rect 165430 75922 165498 75978
rect 165554 75922 165622 75978
rect 165678 75922 183250 75978
rect 183306 75922 183374 75978
rect 183430 75922 183498 75978
rect 183554 75922 183622 75978
rect 183678 75922 201250 75978
rect 201306 75922 201374 75978
rect 201430 75922 201498 75978
rect 201554 75922 201622 75978
rect 201678 75922 219250 75978
rect 219306 75922 219374 75978
rect 219430 75922 219498 75978
rect 219554 75922 219622 75978
rect 219678 75922 237250 75978
rect 237306 75922 237374 75978
rect 237430 75922 237498 75978
rect 237554 75922 237622 75978
rect 237678 75922 255250 75978
rect 255306 75922 255374 75978
rect 255430 75922 255498 75978
rect 255554 75922 255622 75978
rect 255678 75922 273250 75978
rect 273306 75922 273374 75978
rect 273430 75922 273498 75978
rect 273554 75922 273622 75978
rect 273678 75922 291250 75978
rect 291306 75922 291374 75978
rect 291430 75922 291498 75978
rect 291554 75922 291622 75978
rect 291678 75922 309250 75978
rect 309306 75922 309374 75978
rect 309430 75922 309498 75978
rect 309554 75922 309622 75978
rect 309678 75922 327250 75978
rect 327306 75922 327374 75978
rect 327430 75922 327498 75978
rect 327554 75922 327622 75978
rect 327678 75922 345250 75978
rect 345306 75922 345374 75978
rect 345430 75922 345498 75978
rect 345554 75922 345622 75978
rect 345678 75922 363250 75978
rect 363306 75922 363374 75978
rect 363430 75922 363498 75978
rect 363554 75922 363622 75978
rect 363678 75922 381250 75978
rect 381306 75922 381374 75978
rect 381430 75922 381498 75978
rect 381554 75922 381622 75978
rect 381678 75922 399250 75978
rect 399306 75922 399374 75978
rect 399430 75922 399498 75978
rect 399554 75922 399622 75978
rect 399678 75922 417250 75978
rect 417306 75922 417374 75978
rect 417430 75922 417498 75978
rect 417554 75922 417622 75978
rect 417678 75922 435250 75978
rect 435306 75922 435374 75978
rect 435430 75922 435498 75978
rect 435554 75922 435622 75978
rect 435678 75922 453250 75978
rect 453306 75922 453374 75978
rect 453430 75922 453498 75978
rect 453554 75922 453622 75978
rect 453678 75922 471250 75978
rect 471306 75922 471374 75978
rect 471430 75922 471498 75978
rect 471554 75922 471622 75978
rect 471678 75922 489250 75978
rect 489306 75922 489374 75978
rect 489430 75922 489498 75978
rect 489554 75922 489622 75978
rect 489678 75922 507250 75978
rect 507306 75922 507374 75978
rect 507430 75922 507498 75978
rect 507554 75922 507622 75978
rect 507678 75922 525250 75978
rect 525306 75922 525374 75978
rect 525430 75922 525498 75978
rect 525554 75922 525622 75978
rect 525678 75922 543250 75978
rect 543306 75922 543374 75978
rect 543430 75922 543498 75978
rect 543554 75922 543622 75978
rect 543678 75922 561250 75978
rect 561306 75922 561374 75978
rect 561430 75922 561498 75978
rect 561554 75922 561622 75978
rect 561678 75922 579250 75978
rect 579306 75922 579374 75978
rect 579430 75922 579498 75978
rect 579554 75922 579622 75978
rect 579678 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 6970 64350
rect 7026 64294 7094 64350
rect 7150 64294 7218 64350
rect 7274 64294 7342 64350
rect 7398 64294 24970 64350
rect 25026 64294 25094 64350
rect 25150 64294 25218 64350
rect 25274 64294 25342 64350
rect 25398 64294 42970 64350
rect 43026 64294 43094 64350
rect 43150 64294 43218 64350
rect 43274 64294 43342 64350
rect 43398 64294 60970 64350
rect 61026 64294 61094 64350
rect 61150 64294 61218 64350
rect 61274 64294 61342 64350
rect 61398 64294 78970 64350
rect 79026 64294 79094 64350
rect 79150 64294 79218 64350
rect 79274 64294 79342 64350
rect 79398 64294 96970 64350
rect 97026 64294 97094 64350
rect 97150 64294 97218 64350
rect 97274 64294 97342 64350
rect 97398 64294 114970 64350
rect 115026 64294 115094 64350
rect 115150 64294 115218 64350
rect 115274 64294 115342 64350
rect 115398 64294 132970 64350
rect 133026 64294 133094 64350
rect 133150 64294 133218 64350
rect 133274 64294 133342 64350
rect 133398 64294 150970 64350
rect 151026 64294 151094 64350
rect 151150 64294 151218 64350
rect 151274 64294 151342 64350
rect 151398 64294 168970 64350
rect 169026 64294 169094 64350
rect 169150 64294 169218 64350
rect 169274 64294 169342 64350
rect 169398 64294 186970 64350
rect 187026 64294 187094 64350
rect 187150 64294 187218 64350
rect 187274 64294 187342 64350
rect 187398 64294 204970 64350
rect 205026 64294 205094 64350
rect 205150 64294 205218 64350
rect 205274 64294 205342 64350
rect 205398 64294 222970 64350
rect 223026 64294 223094 64350
rect 223150 64294 223218 64350
rect 223274 64294 223342 64350
rect 223398 64294 240970 64350
rect 241026 64294 241094 64350
rect 241150 64294 241218 64350
rect 241274 64294 241342 64350
rect 241398 64294 258970 64350
rect 259026 64294 259094 64350
rect 259150 64294 259218 64350
rect 259274 64294 259342 64350
rect 259398 64294 276970 64350
rect 277026 64294 277094 64350
rect 277150 64294 277218 64350
rect 277274 64294 277342 64350
rect 277398 64294 294970 64350
rect 295026 64294 295094 64350
rect 295150 64294 295218 64350
rect 295274 64294 295342 64350
rect 295398 64294 312970 64350
rect 313026 64294 313094 64350
rect 313150 64294 313218 64350
rect 313274 64294 313342 64350
rect 313398 64294 330970 64350
rect 331026 64294 331094 64350
rect 331150 64294 331218 64350
rect 331274 64294 331342 64350
rect 331398 64294 348970 64350
rect 349026 64294 349094 64350
rect 349150 64294 349218 64350
rect 349274 64294 349342 64350
rect 349398 64294 366970 64350
rect 367026 64294 367094 64350
rect 367150 64294 367218 64350
rect 367274 64294 367342 64350
rect 367398 64294 384970 64350
rect 385026 64294 385094 64350
rect 385150 64294 385218 64350
rect 385274 64294 385342 64350
rect 385398 64294 402970 64350
rect 403026 64294 403094 64350
rect 403150 64294 403218 64350
rect 403274 64294 403342 64350
rect 403398 64294 420970 64350
rect 421026 64294 421094 64350
rect 421150 64294 421218 64350
rect 421274 64294 421342 64350
rect 421398 64294 438970 64350
rect 439026 64294 439094 64350
rect 439150 64294 439218 64350
rect 439274 64294 439342 64350
rect 439398 64294 456970 64350
rect 457026 64294 457094 64350
rect 457150 64294 457218 64350
rect 457274 64294 457342 64350
rect 457398 64294 474970 64350
rect 475026 64294 475094 64350
rect 475150 64294 475218 64350
rect 475274 64294 475342 64350
rect 475398 64294 492970 64350
rect 493026 64294 493094 64350
rect 493150 64294 493218 64350
rect 493274 64294 493342 64350
rect 493398 64294 510970 64350
rect 511026 64294 511094 64350
rect 511150 64294 511218 64350
rect 511274 64294 511342 64350
rect 511398 64294 528970 64350
rect 529026 64294 529094 64350
rect 529150 64294 529218 64350
rect 529274 64294 529342 64350
rect 529398 64294 546970 64350
rect 547026 64294 547094 64350
rect 547150 64294 547218 64350
rect 547274 64294 547342 64350
rect 547398 64294 564970 64350
rect 565026 64294 565094 64350
rect 565150 64294 565218 64350
rect 565274 64294 565342 64350
rect 565398 64294 582970 64350
rect 583026 64294 583094 64350
rect 583150 64294 583218 64350
rect 583274 64294 583342 64350
rect 583398 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 6970 64226
rect 7026 64170 7094 64226
rect 7150 64170 7218 64226
rect 7274 64170 7342 64226
rect 7398 64170 24970 64226
rect 25026 64170 25094 64226
rect 25150 64170 25218 64226
rect 25274 64170 25342 64226
rect 25398 64170 42970 64226
rect 43026 64170 43094 64226
rect 43150 64170 43218 64226
rect 43274 64170 43342 64226
rect 43398 64170 60970 64226
rect 61026 64170 61094 64226
rect 61150 64170 61218 64226
rect 61274 64170 61342 64226
rect 61398 64170 78970 64226
rect 79026 64170 79094 64226
rect 79150 64170 79218 64226
rect 79274 64170 79342 64226
rect 79398 64170 96970 64226
rect 97026 64170 97094 64226
rect 97150 64170 97218 64226
rect 97274 64170 97342 64226
rect 97398 64170 114970 64226
rect 115026 64170 115094 64226
rect 115150 64170 115218 64226
rect 115274 64170 115342 64226
rect 115398 64170 132970 64226
rect 133026 64170 133094 64226
rect 133150 64170 133218 64226
rect 133274 64170 133342 64226
rect 133398 64170 150970 64226
rect 151026 64170 151094 64226
rect 151150 64170 151218 64226
rect 151274 64170 151342 64226
rect 151398 64170 168970 64226
rect 169026 64170 169094 64226
rect 169150 64170 169218 64226
rect 169274 64170 169342 64226
rect 169398 64170 186970 64226
rect 187026 64170 187094 64226
rect 187150 64170 187218 64226
rect 187274 64170 187342 64226
rect 187398 64170 204970 64226
rect 205026 64170 205094 64226
rect 205150 64170 205218 64226
rect 205274 64170 205342 64226
rect 205398 64170 222970 64226
rect 223026 64170 223094 64226
rect 223150 64170 223218 64226
rect 223274 64170 223342 64226
rect 223398 64170 240970 64226
rect 241026 64170 241094 64226
rect 241150 64170 241218 64226
rect 241274 64170 241342 64226
rect 241398 64170 258970 64226
rect 259026 64170 259094 64226
rect 259150 64170 259218 64226
rect 259274 64170 259342 64226
rect 259398 64170 276970 64226
rect 277026 64170 277094 64226
rect 277150 64170 277218 64226
rect 277274 64170 277342 64226
rect 277398 64170 294970 64226
rect 295026 64170 295094 64226
rect 295150 64170 295218 64226
rect 295274 64170 295342 64226
rect 295398 64170 312970 64226
rect 313026 64170 313094 64226
rect 313150 64170 313218 64226
rect 313274 64170 313342 64226
rect 313398 64170 330970 64226
rect 331026 64170 331094 64226
rect 331150 64170 331218 64226
rect 331274 64170 331342 64226
rect 331398 64170 348970 64226
rect 349026 64170 349094 64226
rect 349150 64170 349218 64226
rect 349274 64170 349342 64226
rect 349398 64170 366970 64226
rect 367026 64170 367094 64226
rect 367150 64170 367218 64226
rect 367274 64170 367342 64226
rect 367398 64170 384970 64226
rect 385026 64170 385094 64226
rect 385150 64170 385218 64226
rect 385274 64170 385342 64226
rect 385398 64170 402970 64226
rect 403026 64170 403094 64226
rect 403150 64170 403218 64226
rect 403274 64170 403342 64226
rect 403398 64170 420970 64226
rect 421026 64170 421094 64226
rect 421150 64170 421218 64226
rect 421274 64170 421342 64226
rect 421398 64170 438970 64226
rect 439026 64170 439094 64226
rect 439150 64170 439218 64226
rect 439274 64170 439342 64226
rect 439398 64170 456970 64226
rect 457026 64170 457094 64226
rect 457150 64170 457218 64226
rect 457274 64170 457342 64226
rect 457398 64170 474970 64226
rect 475026 64170 475094 64226
rect 475150 64170 475218 64226
rect 475274 64170 475342 64226
rect 475398 64170 492970 64226
rect 493026 64170 493094 64226
rect 493150 64170 493218 64226
rect 493274 64170 493342 64226
rect 493398 64170 510970 64226
rect 511026 64170 511094 64226
rect 511150 64170 511218 64226
rect 511274 64170 511342 64226
rect 511398 64170 528970 64226
rect 529026 64170 529094 64226
rect 529150 64170 529218 64226
rect 529274 64170 529342 64226
rect 529398 64170 546970 64226
rect 547026 64170 547094 64226
rect 547150 64170 547218 64226
rect 547274 64170 547342 64226
rect 547398 64170 564970 64226
rect 565026 64170 565094 64226
rect 565150 64170 565218 64226
rect 565274 64170 565342 64226
rect 565398 64170 582970 64226
rect 583026 64170 583094 64226
rect 583150 64170 583218 64226
rect 583274 64170 583342 64226
rect 583398 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 6970 64102
rect 7026 64046 7094 64102
rect 7150 64046 7218 64102
rect 7274 64046 7342 64102
rect 7398 64046 24970 64102
rect 25026 64046 25094 64102
rect 25150 64046 25218 64102
rect 25274 64046 25342 64102
rect 25398 64046 42970 64102
rect 43026 64046 43094 64102
rect 43150 64046 43218 64102
rect 43274 64046 43342 64102
rect 43398 64046 60970 64102
rect 61026 64046 61094 64102
rect 61150 64046 61218 64102
rect 61274 64046 61342 64102
rect 61398 64046 78970 64102
rect 79026 64046 79094 64102
rect 79150 64046 79218 64102
rect 79274 64046 79342 64102
rect 79398 64046 96970 64102
rect 97026 64046 97094 64102
rect 97150 64046 97218 64102
rect 97274 64046 97342 64102
rect 97398 64046 114970 64102
rect 115026 64046 115094 64102
rect 115150 64046 115218 64102
rect 115274 64046 115342 64102
rect 115398 64046 132970 64102
rect 133026 64046 133094 64102
rect 133150 64046 133218 64102
rect 133274 64046 133342 64102
rect 133398 64046 150970 64102
rect 151026 64046 151094 64102
rect 151150 64046 151218 64102
rect 151274 64046 151342 64102
rect 151398 64046 168970 64102
rect 169026 64046 169094 64102
rect 169150 64046 169218 64102
rect 169274 64046 169342 64102
rect 169398 64046 186970 64102
rect 187026 64046 187094 64102
rect 187150 64046 187218 64102
rect 187274 64046 187342 64102
rect 187398 64046 204970 64102
rect 205026 64046 205094 64102
rect 205150 64046 205218 64102
rect 205274 64046 205342 64102
rect 205398 64046 222970 64102
rect 223026 64046 223094 64102
rect 223150 64046 223218 64102
rect 223274 64046 223342 64102
rect 223398 64046 240970 64102
rect 241026 64046 241094 64102
rect 241150 64046 241218 64102
rect 241274 64046 241342 64102
rect 241398 64046 258970 64102
rect 259026 64046 259094 64102
rect 259150 64046 259218 64102
rect 259274 64046 259342 64102
rect 259398 64046 276970 64102
rect 277026 64046 277094 64102
rect 277150 64046 277218 64102
rect 277274 64046 277342 64102
rect 277398 64046 294970 64102
rect 295026 64046 295094 64102
rect 295150 64046 295218 64102
rect 295274 64046 295342 64102
rect 295398 64046 312970 64102
rect 313026 64046 313094 64102
rect 313150 64046 313218 64102
rect 313274 64046 313342 64102
rect 313398 64046 330970 64102
rect 331026 64046 331094 64102
rect 331150 64046 331218 64102
rect 331274 64046 331342 64102
rect 331398 64046 348970 64102
rect 349026 64046 349094 64102
rect 349150 64046 349218 64102
rect 349274 64046 349342 64102
rect 349398 64046 366970 64102
rect 367026 64046 367094 64102
rect 367150 64046 367218 64102
rect 367274 64046 367342 64102
rect 367398 64046 384970 64102
rect 385026 64046 385094 64102
rect 385150 64046 385218 64102
rect 385274 64046 385342 64102
rect 385398 64046 402970 64102
rect 403026 64046 403094 64102
rect 403150 64046 403218 64102
rect 403274 64046 403342 64102
rect 403398 64046 420970 64102
rect 421026 64046 421094 64102
rect 421150 64046 421218 64102
rect 421274 64046 421342 64102
rect 421398 64046 438970 64102
rect 439026 64046 439094 64102
rect 439150 64046 439218 64102
rect 439274 64046 439342 64102
rect 439398 64046 456970 64102
rect 457026 64046 457094 64102
rect 457150 64046 457218 64102
rect 457274 64046 457342 64102
rect 457398 64046 474970 64102
rect 475026 64046 475094 64102
rect 475150 64046 475218 64102
rect 475274 64046 475342 64102
rect 475398 64046 492970 64102
rect 493026 64046 493094 64102
rect 493150 64046 493218 64102
rect 493274 64046 493342 64102
rect 493398 64046 510970 64102
rect 511026 64046 511094 64102
rect 511150 64046 511218 64102
rect 511274 64046 511342 64102
rect 511398 64046 528970 64102
rect 529026 64046 529094 64102
rect 529150 64046 529218 64102
rect 529274 64046 529342 64102
rect 529398 64046 546970 64102
rect 547026 64046 547094 64102
rect 547150 64046 547218 64102
rect 547274 64046 547342 64102
rect 547398 64046 564970 64102
rect 565026 64046 565094 64102
rect 565150 64046 565218 64102
rect 565274 64046 565342 64102
rect 565398 64046 582970 64102
rect 583026 64046 583094 64102
rect 583150 64046 583218 64102
rect 583274 64046 583342 64102
rect 583398 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 6970 63978
rect 7026 63922 7094 63978
rect 7150 63922 7218 63978
rect 7274 63922 7342 63978
rect 7398 63922 24970 63978
rect 25026 63922 25094 63978
rect 25150 63922 25218 63978
rect 25274 63922 25342 63978
rect 25398 63922 42970 63978
rect 43026 63922 43094 63978
rect 43150 63922 43218 63978
rect 43274 63922 43342 63978
rect 43398 63922 60970 63978
rect 61026 63922 61094 63978
rect 61150 63922 61218 63978
rect 61274 63922 61342 63978
rect 61398 63922 78970 63978
rect 79026 63922 79094 63978
rect 79150 63922 79218 63978
rect 79274 63922 79342 63978
rect 79398 63922 96970 63978
rect 97026 63922 97094 63978
rect 97150 63922 97218 63978
rect 97274 63922 97342 63978
rect 97398 63922 114970 63978
rect 115026 63922 115094 63978
rect 115150 63922 115218 63978
rect 115274 63922 115342 63978
rect 115398 63922 132970 63978
rect 133026 63922 133094 63978
rect 133150 63922 133218 63978
rect 133274 63922 133342 63978
rect 133398 63922 150970 63978
rect 151026 63922 151094 63978
rect 151150 63922 151218 63978
rect 151274 63922 151342 63978
rect 151398 63922 168970 63978
rect 169026 63922 169094 63978
rect 169150 63922 169218 63978
rect 169274 63922 169342 63978
rect 169398 63922 186970 63978
rect 187026 63922 187094 63978
rect 187150 63922 187218 63978
rect 187274 63922 187342 63978
rect 187398 63922 204970 63978
rect 205026 63922 205094 63978
rect 205150 63922 205218 63978
rect 205274 63922 205342 63978
rect 205398 63922 222970 63978
rect 223026 63922 223094 63978
rect 223150 63922 223218 63978
rect 223274 63922 223342 63978
rect 223398 63922 240970 63978
rect 241026 63922 241094 63978
rect 241150 63922 241218 63978
rect 241274 63922 241342 63978
rect 241398 63922 258970 63978
rect 259026 63922 259094 63978
rect 259150 63922 259218 63978
rect 259274 63922 259342 63978
rect 259398 63922 276970 63978
rect 277026 63922 277094 63978
rect 277150 63922 277218 63978
rect 277274 63922 277342 63978
rect 277398 63922 294970 63978
rect 295026 63922 295094 63978
rect 295150 63922 295218 63978
rect 295274 63922 295342 63978
rect 295398 63922 312970 63978
rect 313026 63922 313094 63978
rect 313150 63922 313218 63978
rect 313274 63922 313342 63978
rect 313398 63922 330970 63978
rect 331026 63922 331094 63978
rect 331150 63922 331218 63978
rect 331274 63922 331342 63978
rect 331398 63922 348970 63978
rect 349026 63922 349094 63978
rect 349150 63922 349218 63978
rect 349274 63922 349342 63978
rect 349398 63922 366970 63978
rect 367026 63922 367094 63978
rect 367150 63922 367218 63978
rect 367274 63922 367342 63978
rect 367398 63922 384970 63978
rect 385026 63922 385094 63978
rect 385150 63922 385218 63978
rect 385274 63922 385342 63978
rect 385398 63922 402970 63978
rect 403026 63922 403094 63978
rect 403150 63922 403218 63978
rect 403274 63922 403342 63978
rect 403398 63922 420970 63978
rect 421026 63922 421094 63978
rect 421150 63922 421218 63978
rect 421274 63922 421342 63978
rect 421398 63922 438970 63978
rect 439026 63922 439094 63978
rect 439150 63922 439218 63978
rect 439274 63922 439342 63978
rect 439398 63922 456970 63978
rect 457026 63922 457094 63978
rect 457150 63922 457218 63978
rect 457274 63922 457342 63978
rect 457398 63922 474970 63978
rect 475026 63922 475094 63978
rect 475150 63922 475218 63978
rect 475274 63922 475342 63978
rect 475398 63922 492970 63978
rect 493026 63922 493094 63978
rect 493150 63922 493218 63978
rect 493274 63922 493342 63978
rect 493398 63922 510970 63978
rect 511026 63922 511094 63978
rect 511150 63922 511218 63978
rect 511274 63922 511342 63978
rect 511398 63922 528970 63978
rect 529026 63922 529094 63978
rect 529150 63922 529218 63978
rect 529274 63922 529342 63978
rect 529398 63922 546970 63978
rect 547026 63922 547094 63978
rect 547150 63922 547218 63978
rect 547274 63922 547342 63978
rect 547398 63922 564970 63978
rect 565026 63922 565094 63978
rect 565150 63922 565218 63978
rect 565274 63922 565342 63978
rect 565398 63922 582970 63978
rect 583026 63922 583094 63978
rect 583150 63922 583218 63978
rect 583274 63922 583342 63978
rect 583398 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 3250 58350
rect 3306 58294 3374 58350
rect 3430 58294 3498 58350
rect 3554 58294 3622 58350
rect 3678 58294 21250 58350
rect 21306 58294 21374 58350
rect 21430 58294 21498 58350
rect 21554 58294 21622 58350
rect 21678 58294 39250 58350
rect 39306 58294 39374 58350
rect 39430 58294 39498 58350
rect 39554 58294 39622 58350
rect 39678 58294 57250 58350
rect 57306 58294 57374 58350
rect 57430 58294 57498 58350
rect 57554 58294 57622 58350
rect 57678 58294 75250 58350
rect 75306 58294 75374 58350
rect 75430 58294 75498 58350
rect 75554 58294 75622 58350
rect 75678 58294 93250 58350
rect 93306 58294 93374 58350
rect 93430 58294 93498 58350
rect 93554 58294 93622 58350
rect 93678 58294 111250 58350
rect 111306 58294 111374 58350
rect 111430 58294 111498 58350
rect 111554 58294 111622 58350
rect 111678 58294 129250 58350
rect 129306 58294 129374 58350
rect 129430 58294 129498 58350
rect 129554 58294 129622 58350
rect 129678 58294 147250 58350
rect 147306 58294 147374 58350
rect 147430 58294 147498 58350
rect 147554 58294 147622 58350
rect 147678 58294 165250 58350
rect 165306 58294 165374 58350
rect 165430 58294 165498 58350
rect 165554 58294 165622 58350
rect 165678 58294 183250 58350
rect 183306 58294 183374 58350
rect 183430 58294 183498 58350
rect 183554 58294 183622 58350
rect 183678 58294 201250 58350
rect 201306 58294 201374 58350
rect 201430 58294 201498 58350
rect 201554 58294 201622 58350
rect 201678 58294 219250 58350
rect 219306 58294 219374 58350
rect 219430 58294 219498 58350
rect 219554 58294 219622 58350
rect 219678 58294 237250 58350
rect 237306 58294 237374 58350
rect 237430 58294 237498 58350
rect 237554 58294 237622 58350
rect 237678 58294 255250 58350
rect 255306 58294 255374 58350
rect 255430 58294 255498 58350
rect 255554 58294 255622 58350
rect 255678 58294 273250 58350
rect 273306 58294 273374 58350
rect 273430 58294 273498 58350
rect 273554 58294 273622 58350
rect 273678 58294 291250 58350
rect 291306 58294 291374 58350
rect 291430 58294 291498 58350
rect 291554 58294 291622 58350
rect 291678 58294 309250 58350
rect 309306 58294 309374 58350
rect 309430 58294 309498 58350
rect 309554 58294 309622 58350
rect 309678 58294 327250 58350
rect 327306 58294 327374 58350
rect 327430 58294 327498 58350
rect 327554 58294 327622 58350
rect 327678 58294 345250 58350
rect 345306 58294 345374 58350
rect 345430 58294 345498 58350
rect 345554 58294 345622 58350
rect 345678 58294 363250 58350
rect 363306 58294 363374 58350
rect 363430 58294 363498 58350
rect 363554 58294 363622 58350
rect 363678 58294 381250 58350
rect 381306 58294 381374 58350
rect 381430 58294 381498 58350
rect 381554 58294 381622 58350
rect 381678 58294 399250 58350
rect 399306 58294 399374 58350
rect 399430 58294 399498 58350
rect 399554 58294 399622 58350
rect 399678 58294 417250 58350
rect 417306 58294 417374 58350
rect 417430 58294 417498 58350
rect 417554 58294 417622 58350
rect 417678 58294 435250 58350
rect 435306 58294 435374 58350
rect 435430 58294 435498 58350
rect 435554 58294 435622 58350
rect 435678 58294 453250 58350
rect 453306 58294 453374 58350
rect 453430 58294 453498 58350
rect 453554 58294 453622 58350
rect 453678 58294 471250 58350
rect 471306 58294 471374 58350
rect 471430 58294 471498 58350
rect 471554 58294 471622 58350
rect 471678 58294 489250 58350
rect 489306 58294 489374 58350
rect 489430 58294 489498 58350
rect 489554 58294 489622 58350
rect 489678 58294 507250 58350
rect 507306 58294 507374 58350
rect 507430 58294 507498 58350
rect 507554 58294 507622 58350
rect 507678 58294 525250 58350
rect 525306 58294 525374 58350
rect 525430 58294 525498 58350
rect 525554 58294 525622 58350
rect 525678 58294 543250 58350
rect 543306 58294 543374 58350
rect 543430 58294 543498 58350
rect 543554 58294 543622 58350
rect 543678 58294 561250 58350
rect 561306 58294 561374 58350
rect 561430 58294 561498 58350
rect 561554 58294 561622 58350
rect 561678 58294 579250 58350
rect 579306 58294 579374 58350
rect 579430 58294 579498 58350
rect 579554 58294 579622 58350
rect 579678 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 3250 58226
rect 3306 58170 3374 58226
rect 3430 58170 3498 58226
rect 3554 58170 3622 58226
rect 3678 58170 21250 58226
rect 21306 58170 21374 58226
rect 21430 58170 21498 58226
rect 21554 58170 21622 58226
rect 21678 58170 39250 58226
rect 39306 58170 39374 58226
rect 39430 58170 39498 58226
rect 39554 58170 39622 58226
rect 39678 58170 57250 58226
rect 57306 58170 57374 58226
rect 57430 58170 57498 58226
rect 57554 58170 57622 58226
rect 57678 58170 75250 58226
rect 75306 58170 75374 58226
rect 75430 58170 75498 58226
rect 75554 58170 75622 58226
rect 75678 58170 93250 58226
rect 93306 58170 93374 58226
rect 93430 58170 93498 58226
rect 93554 58170 93622 58226
rect 93678 58170 111250 58226
rect 111306 58170 111374 58226
rect 111430 58170 111498 58226
rect 111554 58170 111622 58226
rect 111678 58170 129250 58226
rect 129306 58170 129374 58226
rect 129430 58170 129498 58226
rect 129554 58170 129622 58226
rect 129678 58170 147250 58226
rect 147306 58170 147374 58226
rect 147430 58170 147498 58226
rect 147554 58170 147622 58226
rect 147678 58170 165250 58226
rect 165306 58170 165374 58226
rect 165430 58170 165498 58226
rect 165554 58170 165622 58226
rect 165678 58170 183250 58226
rect 183306 58170 183374 58226
rect 183430 58170 183498 58226
rect 183554 58170 183622 58226
rect 183678 58170 201250 58226
rect 201306 58170 201374 58226
rect 201430 58170 201498 58226
rect 201554 58170 201622 58226
rect 201678 58170 219250 58226
rect 219306 58170 219374 58226
rect 219430 58170 219498 58226
rect 219554 58170 219622 58226
rect 219678 58170 237250 58226
rect 237306 58170 237374 58226
rect 237430 58170 237498 58226
rect 237554 58170 237622 58226
rect 237678 58170 255250 58226
rect 255306 58170 255374 58226
rect 255430 58170 255498 58226
rect 255554 58170 255622 58226
rect 255678 58170 273250 58226
rect 273306 58170 273374 58226
rect 273430 58170 273498 58226
rect 273554 58170 273622 58226
rect 273678 58170 291250 58226
rect 291306 58170 291374 58226
rect 291430 58170 291498 58226
rect 291554 58170 291622 58226
rect 291678 58170 309250 58226
rect 309306 58170 309374 58226
rect 309430 58170 309498 58226
rect 309554 58170 309622 58226
rect 309678 58170 327250 58226
rect 327306 58170 327374 58226
rect 327430 58170 327498 58226
rect 327554 58170 327622 58226
rect 327678 58170 345250 58226
rect 345306 58170 345374 58226
rect 345430 58170 345498 58226
rect 345554 58170 345622 58226
rect 345678 58170 363250 58226
rect 363306 58170 363374 58226
rect 363430 58170 363498 58226
rect 363554 58170 363622 58226
rect 363678 58170 381250 58226
rect 381306 58170 381374 58226
rect 381430 58170 381498 58226
rect 381554 58170 381622 58226
rect 381678 58170 399250 58226
rect 399306 58170 399374 58226
rect 399430 58170 399498 58226
rect 399554 58170 399622 58226
rect 399678 58170 417250 58226
rect 417306 58170 417374 58226
rect 417430 58170 417498 58226
rect 417554 58170 417622 58226
rect 417678 58170 435250 58226
rect 435306 58170 435374 58226
rect 435430 58170 435498 58226
rect 435554 58170 435622 58226
rect 435678 58170 453250 58226
rect 453306 58170 453374 58226
rect 453430 58170 453498 58226
rect 453554 58170 453622 58226
rect 453678 58170 471250 58226
rect 471306 58170 471374 58226
rect 471430 58170 471498 58226
rect 471554 58170 471622 58226
rect 471678 58170 489250 58226
rect 489306 58170 489374 58226
rect 489430 58170 489498 58226
rect 489554 58170 489622 58226
rect 489678 58170 507250 58226
rect 507306 58170 507374 58226
rect 507430 58170 507498 58226
rect 507554 58170 507622 58226
rect 507678 58170 525250 58226
rect 525306 58170 525374 58226
rect 525430 58170 525498 58226
rect 525554 58170 525622 58226
rect 525678 58170 543250 58226
rect 543306 58170 543374 58226
rect 543430 58170 543498 58226
rect 543554 58170 543622 58226
rect 543678 58170 561250 58226
rect 561306 58170 561374 58226
rect 561430 58170 561498 58226
rect 561554 58170 561622 58226
rect 561678 58170 579250 58226
rect 579306 58170 579374 58226
rect 579430 58170 579498 58226
rect 579554 58170 579622 58226
rect 579678 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 3250 58102
rect 3306 58046 3374 58102
rect 3430 58046 3498 58102
rect 3554 58046 3622 58102
rect 3678 58046 21250 58102
rect 21306 58046 21374 58102
rect 21430 58046 21498 58102
rect 21554 58046 21622 58102
rect 21678 58046 39250 58102
rect 39306 58046 39374 58102
rect 39430 58046 39498 58102
rect 39554 58046 39622 58102
rect 39678 58046 57250 58102
rect 57306 58046 57374 58102
rect 57430 58046 57498 58102
rect 57554 58046 57622 58102
rect 57678 58046 75250 58102
rect 75306 58046 75374 58102
rect 75430 58046 75498 58102
rect 75554 58046 75622 58102
rect 75678 58046 93250 58102
rect 93306 58046 93374 58102
rect 93430 58046 93498 58102
rect 93554 58046 93622 58102
rect 93678 58046 111250 58102
rect 111306 58046 111374 58102
rect 111430 58046 111498 58102
rect 111554 58046 111622 58102
rect 111678 58046 129250 58102
rect 129306 58046 129374 58102
rect 129430 58046 129498 58102
rect 129554 58046 129622 58102
rect 129678 58046 147250 58102
rect 147306 58046 147374 58102
rect 147430 58046 147498 58102
rect 147554 58046 147622 58102
rect 147678 58046 165250 58102
rect 165306 58046 165374 58102
rect 165430 58046 165498 58102
rect 165554 58046 165622 58102
rect 165678 58046 183250 58102
rect 183306 58046 183374 58102
rect 183430 58046 183498 58102
rect 183554 58046 183622 58102
rect 183678 58046 201250 58102
rect 201306 58046 201374 58102
rect 201430 58046 201498 58102
rect 201554 58046 201622 58102
rect 201678 58046 219250 58102
rect 219306 58046 219374 58102
rect 219430 58046 219498 58102
rect 219554 58046 219622 58102
rect 219678 58046 237250 58102
rect 237306 58046 237374 58102
rect 237430 58046 237498 58102
rect 237554 58046 237622 58102
rect 237678 58046 255250 58102
rect 255306 58046 255374 58102
rect 255430 58046 255498 58102
rect 255554 58046 255622 58102
rect 255678 58046 273250 58102
rect 273306 58046 273374 58102
rect 273430 58046 273498 58102
rect 273554 58046 273622 58102
rect 273678 58046 291250 58102
rect 291306 58046 291374 58102
rect 291430 58046 291498 58102
rect 291554 58046 291622 58102
rect 291678 58046 309250 58102
rect 309306 58046 309374 58102
rect 309430 58046 309498 58102
rect 309554 58046 309622 58102
rect 309678 58046 327250 58102
rect 327306 58046 327374 58102
rect 327430 58046 327498 58102
rect 327554 58046 327622 58102
rect 327678 58046 345250 58102
rect 345306 58046 345374 58102
rect 345430 58046 345498 58102
rect 345554 58046 345622 58102
rect 345678 58046 363250 58102
rect 363306 58046 363374 58102
rect 363430 58046 363498 58102
rect 363554 58046 363622 58102
rect 363678 58046 381250 58102
rect 381306 58046 381374 58102
rect 381430 58046 381498 58102
rect 381554 58046 381622 58102
rect 381678 58046 399250 58102
rect 399306 58046 399374 58102
rect 399430 58046 399498 58102
rect 399554 58046 399622 58102
rect 399678 58046 417250 58102
rect 417306 58046 417374 58102
rect 417430 58046 417498 58102
rect 417554 58046 417622 58102
rect 417678 58046 435250 58102
rect 435306 58046 435374 58102
rect 435430 58046 435498 58102
rect 435554 58046 435622 58102
rect 435678 58046 453250 58102
rect 453306 58046 453374 58102
rect 453430 58046 453498 58102
rect 453554 58046 453622 58102
rect 453678 58046 471250 58102
rect 471306 58046 471374 58102
rect 471430 58046 471498 58102
rect 471554 58046 471622 58102
rect 471678 58046 489250 58102
rect 489306 58046 489374 58102
rect 489430 58046 489498 58102
rect 489554 58046 489622 58102
rect 489678 58046 507250 58102
rect 507306 58046 507374 58102
rect 507430 58046 507498 58102
rect 507554 58046 507622 58102
rect 507678 58046 525250 58102
rect 525306 58046 525374 58102
rect 525430 58046 525498 58102
rect 525554 58046 525622 58102
rect 525678 58046 543250 58102
rect 543306 58046 543374 58102
rect 543430 58046 543498 58102
rect 543554 58046 543622 58102
rect 543678 58046 561250 58102
rect 561306 58046 561374 58102
rect 561430 58046 561498 58102
rect 561554 58046 561622 58102
rect 561678 58046 579250 58102
rect 579306 58046 579374 58102
rect 579430 58046 579498 58102
rect 579554 58046 579622 58102
rect 579678 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 3250 57978
rect 3306 57922 3374 57978
rect 3430 57922 3498 57978
rect 3554 57922 3622 57978
rect 3678 57922 21250 57978
rect 21306 57922 21374 57978
rect 21430 57922 21498 57978
rect 21554 57922 21622 57978
rect 21678 57922 39250 57978
rect 39306 57922 39374 57978
rect 39430 57922 39498 57978
rect 39554 57922 39622 57978
rect 39678 57922 57250 57978
rect 57306 57922 57374 57978
rect 57430 57922 57498 57978
rect 57554 57922 57622 57978
rect 57678 57922 75250 57978
rect 75306 57922 75374 57978
rect 75430 57922 75498 57978
rect 75554 57922 75622 57978
rect 75678 57922 93250 57978
rect 93306 57922 93374 57978
rect 93430 57922 93498 57978
rect 93554 57922 93622 57978
rect 93678 57922 111250 57978
rect 111306 57922 111374 57978
rect 111430 57922 111498 57978
rect 111554 57922 111622 57978
rect 111678 57922 129250 57978
rect 129306 57922 129374 57978
rect 129430 57922 129498 57978
rect 129554 57922 129622 57978
rect 129678 57922 147250 57978
rect 147306 57922 147374 57978
rect 147430 57922 147498 57978
rect 147554 57922 147622 57978
rect 147678 57922 165250 57978
rect 165306 57922 165374 57978
rect 165430 57922 165498 57978
rect 165554 57922 165622 57978
rect 165678 57922 183250 57978
rect 183306 57922 183374 57978
rect 183430 57922 183498 57978
rect 183554 57922 183622 57978
rect 183678 57922 201250 57978
rect 201306 57922 201374 57978
rect 201430 57922 201498 57978
rect 201554 57922 201622 57978
rect 201678 57922 219250 57978
rect 219306 57922 219374 57978
rect 219430 57922 219498 57978
rect 219554 57922 219622 57978
rect 219678 57922 237250 57978
rect 237306 57922 237374 57978
rect 237430 57922 237498 57978
rect 237554 57922 237622 57978
rect 237678 57922 255250 57978
rect 255306 57922 255374 57978
rect 255430 57922 255498 57978
rect 255554 57922 255622 57978
rect 255678 57922 273250 57978
rect 273306 57922 273374 57978
rect 273430 57922 273498 57978
rect 273554 57922 273622 57978
rect 273678 57922 291250 57978
rect 291306 57922 291374 57978
rect 291430 57922 291498 57978
rect 291554 57922 291622 57978
rect 291678 57922 309250 57978
rect 309306 57922 309374 57978
rect 309430 57922 309498 57978
rect 309554 57922 309622 57978
rect 309678 57922 327250 57978
rect 327306 57922 327374 57978
rect 327430 57922 327498 57978
rect 327554 57922 327622 57978
rect 327678 57922 345250 57978
rect 345306 57922 345374 57978
rect 345430 57922 345498 57978
rect 345554 57922 345622 57978
rect 345678 57922 363250 57978
rect 363306 57922 363374 57978
rect 363430 57922 363498 57978
rect 363554 57922 363622 57978
rect 363678 57922 381250 57978
rect 381306 57922 381374 57978
rect 381430 57922 381498 57978
rect 381554 57922 381622 57978
rect 381678 57922 399250 57978
rect 399306 57922 399374 57978
rect 399430 57922 399498 57978
rect 399554 57922 399622 57978
rect 399678 57922 417250 57978
rect 417306 57922 417374 57978
rect 417430 57922 417498 57978
rect 417554 57922 417622 57978
rect 417678 57922 435250 57978
rect 435306 57922 435374 57978
rect 435430 57922 435498 57978
rect 435554 57922 435622 57978
rect 435678 57922 453250 57978
rect 453306 57922 453374 57978
rect 453430 57922 453498 57978
rect 453554 57922 453622 57978
rect 453678 57922 471250 57978
rect 471306 57922 471374 57978
rect 471430 57922 471498 57978
rect 471554 57922 471622 57978
rect 471678 57922 489250 57978
rect 489306 57922 489374 57978
rect 489430 57922 489498 57978
rect 489554 57922 489622 57978
rect 489678 57922 507250 57978
rect 507306 57922 507374 57978
rect 507430 57922 507498 57978
rect 507554 57922 507622 57978
rect 507678 57922 525250 57978
rect 525306 57922 525374 57978
rect 525430 57922 525498 57978
rect 525554 57922 525622 57978
rect 525678 57922 543250 57978
rect 543306 57922 543374 57978
rect 543430 57922 543498 57978
rect 543554 57922 543622 57978
rect 543678 57922 561250 57978
rect 561306 57922 561374 57978
rect 561430 57922 561498 57978
rect 561554 57922 561622 57978
rect 561678 57922 579250 57978
rect 579306 57922 579374 57978
rect 579430 57922 579498 57978
rect 579554 57922 579622 57978
rect 579678 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 6970 46350
rect 7026 46294 7094 46350
rect 7150 46294 7218 46350
rect 7274 46294 7342 46350
rect 7398 46294 24970 46350
rect 25026 46294 25094 46350
rect 25150 46294 25218 46350
rect 25274 46294 25342 46350
rect 25398 46294 42970 46350
rect 43026 46294 43094 46350
rect 43150 46294 43218 46350
rect 43274 46294 43342 46350
rect 43398 46294 60970 46350
rect 61026 46294 61094 46350
rect 61150 46294 61218 46350
rect 61274 46294 61342 46350
rect 61398 46294 78970 46350
rect 79026 46294 79094 46350
rect 79150 46294 79218 46350
rect 79274 46294 79342 46350
rect 79398 46294 96970 46350
rect 97026 46294 97094 46350
rect 97150 46294 97218 46350
rect 97274 46294 97342 46350
rect 97398 46294 114970 46350
rect 115026 46294 115094 46350
rect 115150 46294 115218 46350
rect 115274 46294 115342 46350
rect 115398 46294 132970 46350
rect 133026 46294 133094 46350
rect 133150 46294 133218 46350
rect 133274 46294 133342 46350
rect 133398 46294 150970 46350
rect 151026 46294 151094 46350
rect 151150 46294 151218 46350
rect 151274 46294 151342 46350
rect 151398 46294 168970 46350
rect 169026 46294 169094 46350
rect 169150 46294 169218 46350
rect 169274 46294 169342 46350
rect 169398 46294 186970 46350
rect 187026 46294 187094 46350
rect 187150 46294 187218 46350
rect 187274 46294 187342 46350
rect 187398 46294 204970 46350
rect 205026 46294 205094 46350
rect 205150 46294 205218 46350
rect 205274 46294 205342 46350
rect 205398 46294 222970 46350
rect 223026 46294 223094 46350
rect 223150 46294 223218 46350
rect 223274 46294 223342 46350
rect 223398 46294 240970 46350
rect 241026 46294 241094 46350
rect 241150 46294 241218 46350
rect 241274 46294 241342 46350
rect 241398 46294 258970 46350
rect 259026 46294 259094 46350
rect 259150 46294 259218 46350
rect 259274 46294 259342 46350
rect 259398 46294 276970 46350
rect 277026 46294 277094 46350
rect 277150 46294 277218 46350
rect 277274 46294 277342 46350
rect 277398 46294 294970 46350
rect 295026 46294 295094 46350
rect 295150 46294 295218 46350
rect 295274 46294 295342 46350
rect 295398 46294 312970 46350
rect 313026 46294 313094 46350
rect 313150 46294 313218 46350
rect 313274 46294 313342 46350
rect 313398 46294 330970 46350
rect 331026 46294 331094 46350
rect 331150 46294 331218 46350
rect 331274 46294 331342 46350
rect 331398 46294 348970 46350
rect 349026 46294 349094 46350
rect 349150 46294 349218 46350
rect 349274 46294 349342 46350
rect 349398 46294 366970 46350
rect 367026 46294 367094 46350
rect 367150 46294 367218 46350
rect 367274 46294 367342 46350
rect 367398 46294 384970 46350
rect 385026 46294 385094 46350
rect 385150 46294 385218 46350
rect 385274 46294 385342 46350
rect 385398 46294 402970 46350
rect 403026 46294 403094 46350
rect 403150 46294 403218 46350
rect 403274 46294 403342 46350
rect 403398 46294 420970 46350
rect 421026 46294 421094 46350
rect 421150 46294 421218 46350
rect 421274 46294 421342 46350
rect 421398 46294 438970 46350
rect 439026 46294 439094 46350
rect 439150 46294 439218 46350
rect 439274 46294 439342 46350
rect 439398 46294 456970 46350
rect 457026 46294 457094 46350
rect 457150 46294 457218 46350
rect 457274 46294 457342 46350
rect 457398 46294 474970 46350
rect 475026 46294 475094 46350
rect 475150 46294 475218 46350
rect 475274 46294 475342 46350
rect 475398 46294 492970 46350
rect 493026 46294 493094 46350
rect 493150 46294 493218 46350
rect 493274 46294 493342 46350
rect 493398 46294 510970 46350
rect 511026 46294 511094 46350
rect 511150 46294 511218 46350
rect 511274 46294 511342 46350
rect 511398 46294 528970 46350
rect 529026 46294 529094 46350
rect 529150 46294 529218 46350
rect 529274 46294 529342 46350
rect 529398 46294 546970 46350
rect 547026 46294 547094 46350
rect 547150 46294 547218 46350
rect 547274 46294 547342 46350
rect 547398 46294 564970 46350
rect 565026 46294 565094 46350
rect 565150 46294 565218 46350
rect 565274 46294 565342 46350
rect 565398 46294 582970 46350
rect 583026 46294 583094 46350
rect 583150 46294 583218 46350
rect 583274 46294 583342 46350
rect 583398 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 6970 46226
rect 7026 46170 7094 46226
rect 7150 46170 7218 46226
rect 7274 46170 7342 46226
rect 7398 46170 24970 46226
rect 25026 46170 25094 46226
rect 25150 46170 25218 46226
rect 25274 46170 25342 46226
rect 25398 46170 42970 46226
rect 43026 46170 43094 46226
rect 43150 46170 43218 46226
rect 43274 46170 43342 46226
rect 43398 46170 60970 46226
rect 61026 46170 61094 46226
rect 61150 46170 61218 46226
rect 61274 46170 61342 46226
rect 61398 46170 78970 46226
rect 79026 46170 79094 46226
rect 79150 46170 79218 46226
rect 79274 46170 79342 46226
rect 79398 46170 96970 46226
rect 97026 46170 97094 46226
rect 97150 46170 97218 46226
rect 97274 46170 97342 46226
rect 97398 46170 114970 46226
rect 115026 46170 115094 46226
rect 115150 46170 115218 46226
rect 115274 46170 115342 46226
rect 115398 46170 132970 46226
rect 133026 46170 133094 46226
rect 133150 46170 133218 46226
rect 133274 46170 133342 46226
rect 133398 46170 150970 46226
rect 151026 46170 151094 46226
rect 151150 46170 151218 46226
rect 151274 46170 151342 46226
rect 151398 46170 168970 46226
rect 169026 46170 169094 46226
rect 169150 46170 169218 46226
rect 169274 46170 169342 46226
rect 169398 46170 186970 46226
rect 187026 46170 187094 46226
rect 187150 46170 187218 46226
rect 187274 46170 187342 46226
rect 187398 46170 204970 46226
rect 205026 46170 205094 46226
rect 205150 46170 205218 46226
rect 205274 46170 205342 46226
rect 205398 46170 222970 46226
rect 223026 46170 223094 46226
rect 223150 46170 223218 46226
rect 223274 46170 223342 46226
rect 223398 46170 240970 46226
rect 241026 46170 241094 46226
rect 241150 46170 241218 46226
rect 241274 46170 241342 46226
rect 241398 46170 258970 46226
rect 259026 46170 259094 46226
rect 259150 46170 259218 46226
rect 259274 46170 259342 46226
rect 259398 46170 276970 46226
rect 277026 46170 277094 46226
rect 277150 46170 277218 46226
rect 277274 46170 277342 46226
rect 277398 46170 294970 46226
rect 295026 46170 295094 46226
rect 295150 46170 295218 46226
rect 295274 46170 295342 46226
rect 295398 46170 312970 46226
rect 313026 46170 313094 46226
rect 313150 46170 313218 46226
rect 313274 46170 313342 46226
rect 313398 46170 330970 46226
rect 331026 46170 331094 46226
rect 331150 46170 331218 46226
rect 331274 46170 331342 46226
rect 331398 46170 348970 46226
rect 349026 46170 349094 46226
rect 349150 46170 349218 46226
rect 349274 46170 349342 46226
rect 349398 46170 366970 46226
rect 367026 46170 367094 46226
rect 367150 46170 367218 46226
rect 367274 46170 367342 46226
rect 367398 46170 384970 46226
rect 385026 46170 385094 46226
rect 385150 46170 385218 46226
rect 385274 46170 385342 46226
rect 385398 46170 402970 46226
rect 403026 46170 403094 46226
rect 403150 46170 403218 46226
rect 403274 46170 403342 46226
rect 403398 46170 420970 46226
rect 421026 46170 421094 46226
rect 421150 46170 421218 46226
rect 421274 46170 421342 46226
rect 421398 46170 438970 46226
rect 439026 46170 439094 46226
rect 439150 46170 439218 46226
rect 439274 46170 439342 46226
rect 439398 46170 456970 46226
rect 457026 46170 457094 46226
rect 457150 46170 457218 46226
rect 457274 46170 457342 46226
rect 457398 46170 474970 46226
rect 475026 46170 475094 46226
rect 475150 46170 475218 46226
rect 475274 46170 475342 46226
rect 475398 46170 492970 46226
rect 493026 46170 493094 46226
rect 493150 46170 493218 46226
rect 493274 46170 493342 46226
rect 493398 46170 510970 46226
rect 511026 46170 511094 46226
rect 511150 46170 511218 46226
rect 511274 46170 511342 46226
rect 511398 46170 528970 46226
rect 529026 46170 529094 46226
rect 529150 46170 529218 46226
rect 529274 46170 529342 46226
rect 529398 46170 546970 46226
rect 547026 46170 547094 46226
rect 547150 46170 547218 46226
rect 547274 46170 547342 46226
rect 547398 46170 564970 46226
rect 565026 46170 565094 46226
rect 565150 46170 565218 46226
rect 565274 46170 565342 46226
rect 565398 46170 582970 46226
rect 583026 46170 583094 46226
rect 583150 46170 583218 46226
rect 583274 46170 583342 46226
rect 583398 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 6970 46102
rect 7026 46046 7094 46102
rect 7150 46046 7218 46102
rect 7274 46046 7342 46102
rect 7398 46046 24970 46102
rect 25026 46046 25094 46102
rect 25150 46046 25218 46102
rect 25274 46046 25342 46102
rect 25398 46046 42970 46102
rect 43026 46046 43094 46102
rect 43150 46046 43218 46102
rect 43274 46046 43342 46102
rect 43398 46046 60970 46102
rect 61026 46046 61094 46102
rect 61150 46046 61218 46102
rect 61274 46046 61342 46102
rect 61398 46046 78970 46102
rect 79026 46046 79094 46102
rect 79150 46046 79218 46102
rect 79274 46046 79342 46102
rect 79398 46046 96970 46102
rect 97026 46046 97094 46102
rect 97150 46046 97218 46102
rect 97274 46046 97342 46102
rect 97398 46046 114970 46102
rect 115026 46046 115094 46102
rect 115150 46046 115218 46102
rect 115274 46046 115342 46102
rect 115398 46046 132970 46102
rect 133026 46046 133094 46102
rect 133150 46046 133218 46102
rect 133274 46046 133342 46102
rect 133398 46046 150970 46102
rect 151026 46046 151094 46102
rect 151150 46046 151218 46102
rect 151274 46046 151342 46102
rect 151398 46046 168970 46102
rect 169026 46046 169094 46102
rect 169150 46046 169218 46102
rect 169274 46046 169342 46102
rect 169398 46046 186970 46102
rect 187026 46046 187094 46102
rect 187150 46046 187218 46102
rect 187274 46046 187342 46102
rect 187398 46046 204970 46102
rect 205026 46046 205094 46102
rect 205150 46046 205218 46102
rect 205274 46046 205342 46102
rect 205398 46046 222970 46102
rect 223026 46046 223094 46102
rect 223150 46046 223218 46102
rect 223274 46046 223342 46102
rect 223398 46046 240970 46102
rect 241026 46046 241094 46102
rect 241150 46046 241218 46102
rect 241274 46046 241342 46102
rect 241398 46046 258970 46102
rect 259026 46046 259094 46102
rect 259150 46046 259218 46102
rect 259274 46046 259342 46102
rect 259398 46046 276970 46102
rect 277026 46046 277094 46102
rect 277150 46046 277218 46102
rect 277274 46046 277342 46102
rect 277398 46046 294970 46102
rect 295026 46046 295094 46102
rect 295150 46046 295218 46102
rect 295274 46046 295342 46102
rect 295398 46046 312970 46102
rect 313026 46046 313094 46102
rect 313150 46046 313218 46102
rect 313274 46046 313342 46102
rect 313398 46046 330970 46102
rect 331026 46046 331094 46102
rect 331150 46046 331218 46102
rect 331274 46046 331342 46102
rect 331398 46046 348970 46102
rect 349026 46046 349094 46102
rect 349150 46046 349218 46102
rect 349274 46046 349342 46102
rect 349398 46046 366970 46102
rect 367026 46046 367094 46102
rect 367150 46046 367218 46102
rect 367274 46046 367342 46102
rect 367398 46046 384970 46102
rect 385026 46046 385094 46102
rect 385150 46046 385218 46102
rect 385274 46046 385342 46102
rect 385398 46046 402970 46102
rect 403026 46046 403094 46102
rect 403150 46046 403218 46102
rect 403274 46046 403342 46102
rect 403398 46046 420970 46102
rect 421026 46046 421094 46102
rect 421150 46046 421218 46102
rect 421274 46046 421342 46102
rect 421398 46046 438970 46102
rect 439026 46046 439094 46102
rect 439150 46046 439218 46102
rect 439274 46046 439342 46102
rect 439398 46046 456970 46102
rect 457026 46046 457094 46102
rect 457150 46046 457218 46102
rect 457274 46046 457342 46102
rect 457398 46046 474970 46102
rect 475026 46046 475094 46102
rect 475150 46046 475218 46102
rect 475274 46046 475342 46102
rect 475398 46046 492970 46102
rect 493026 46046 493094 46102
rect 493150 46046 493218 46102
rect 493274 46046 493342 46102
rect 493398 46046 510970 46102
rect 511026 46046 511094 46102
rect 511150 46046 511218 46102
rect 511274 46046 511342 46102
rect 511398 46046 528970 46102
rect 529026 46046 529094 46102
rect 529150 46046 529218 46102
rect 529274 46046 529342 46102
rect 529398 46046 546970 46102
rect 547026 46046 547094 46102
rect 547150 46046 547218 46102
rect 547274 46046 547342 46102
rect 547398 46046 564970 46102
rect 565026 46046 565094 46102
rect 565150 46046 565218 46102
rect 565274 46046 565342 46102
rect 565398 46046 582970 46102
rect 583026 46046 583094 46102
rect 583150 46046 583218 46102
rect 583274 46046 583342 46102
rect 583398 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 6970 45978
rect 7026 45922 7094 45978
rect 7150 45922 7218 45978
rect 7274 45922 7342 45978
rect 7398 45922 24970 45978
rect 25026 45922 25094 45978
rect 25150 45922 25218 45978
rect 25274 45922 25342 45978
rect 25398 45922 42970 45978
rect 43026 45922 43094 45978
rect 43150 45922 43218 45978
rect 43274 45922 43342 45978
rect 43398 45922 60970 45978
rect 61026 45922 61094 45978
rect 61150 45922 61218 45978
rect 61274 45922 61342 45978
rect 61398 45922 78970 45978
rect 79026 45922 79094 45978
rect 79150 45922 79218 45978
rect 79274 45922 79342 45978
rect 79398 45922 96970 45978
rect 97026 45922 97094 45978
rect 97150 45922 97218 45978
rect 97274 45922 97342 45978
rect 97398 45922 114970 45978
rect 115026 45922 115094 45978
rect 115150 45922 115218 45978
rect 115274 45922 115342 45978
rect 115398 45922 132970 45978
rect 133026 45922 133094 45978
rect 133150 45922 133218 45978
rect 133274 45922 133342 45978
rect 133398 45922 150970 45978
rect 151026 45922 151094 45978
rect 151150 45922 151218 45978
rect 151274 45922 151342 45978
rect 151398 45922 168970 45978
rect 169026 45922 169094 45978
rect 169150 45922 169218 45978
rect 169274 45922 169342 45978
rect 169398 45922 186970 45978
rect 187026 45922 187094 45978
rect 187150 45922 187218 45978
rect 187274 45922 187342 45978
rect 187398 45922 204970 45978
rect 205026 45922 205094 45978
rect 205150 45922 205218 45978
rect 205274 45922 205342 45978
rect 205398 45922 222970 45978
rect 223026 45922 223094 45978
rect 223150 45922 223218 45978
rect 223274 45922 223342 45978
rect 223398 45922 240970 45978
rect 241026 45922 241094 45978
rect 241150 45922 241218 45978
rect 241274 45922 241342 45978
rect 241398 45922 258970 45978
rect 259026 45922 259094 45978
rect 259150 45922 259218 45978
rect 259274 45922 259342 45978
rect 259398 45922 276970 45978
rect 277026 45922 277094 45978
rect 277150 45922 277218 45978
rect 277274 45922 277342 45978
rect 277398 45922 294970 45978
rect 295026 45922 295094 45978
rect 295150 45922 295218 45978
rect 295274 45922 295342 45978
rect 295398 45922 312970 45978
rect 313026 45922 313094 45978
rect 313150 45922 313218 45978
rect 313274 45922 313342 45978
rect 313398 45922 330970 45978
rect 331026 45922 331094 45978
rect 331150 45922 331218 45978
rect 331274 45922 331342 45978
rect 331398 45922 348970 45978
rect 349026 45922 349094 45978
rect 349150 45922 349218 45978
rect 349274 45922 349342 45978
rect 349398 45922 366970 45978
rect 367026 45922 367094 45978
rect 367150 45922 367218 45978
rect 367274 45922 367342 45978
rect 367398 45922 384970 45978
rect 385026 45922 385094 45978
rect 385150 45922 385218 45978
rect 385274 45922 385342 45978
rect 385398 45922 402970 45978
rect 403026 45922 403094 45978
rect 403150 45922 403218 45978
rect 403274 45922 403342 45978
rect 403398 45922 420970 45978
rect 421026 45922 421094 45978
rect 421150 45922 421218 45978
rect 421274 45922 421342 45978
rect 421398 45922 438970 45978
rect 439026 45922 439094 45978
rect 439150 45922 439218 45978
rect 439274 45922 439342 45978
rect 439398 45922 456970 45978
rect 457026 45922 457094 45978
rect 457150 45922 457218 45978
rect 457274 45922 457342 45978
rect 457398 45922 474970 45978
rect 475026 45922 475094 45978
rect 475150 45922 475218 45978
rect 475274 45922 475342 45978
rect 475398 45922 492970 45978
rect 493026 45922 493094 45978
rect 493150 45922 493218 45978
rect 493274 45922 493342 45978
rect 493398 45922 510970 45978
rect 511026 45922 511094 45978
rect 511150 45922 511218 45978
rect 511274 45922 511342 45978
rect 511398 45922 528970 45978
rect 529026 45922 529094 45978
rect 529150 45922 529218 45978
rect 529274 45922 529342 45978
rect 529398 45922 546970 45978
rect 547026 45922 547094 45978
rect 547150 45922 547218 45978
rect 547274 45922 547342 45978
rect 547398 45922 564970 45978
rect 565026 45922 565094 45978
rect 565150 45922 565218 45978
rect 565274 45922 565342 45978
rect 565398 45922 582970 45978
rect 583026 45922 583094 45978
rect 583150 45922 583218 45978
rect 583274 45922 583342 45978
rect 583398 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 3250 40350
rect 3306 40294 3374 40350
rect 3430 40294 3498 40350
rect 3554 40294 3622 40350
rect 3678 40294 21250 40350
rect 21306 40294 21374 40350
rect 21430 40294 21498 40350
rect 21554 40294 21622 40350
rect 21678 40294 39250 40350
rect 39306 40294 39374 40350
rect 39430 40294 39498 40350
rect 39554 40294 39622 40350
rect 39678 40294 57250 40350
rect 57306 40294 57374 40350
rect 57430 40294 57498 40350
rect 57554 40294 57622 40350
rect 57678 40294 75250 40350
rect 75306 40294 75374 40350
rect 75430 40294 75498 40350
rect 75554 40294 75622 40350
rect 75678 40294 93250 40350
rect 93306 40294 93374 40350
rect 93430 40294 93498 40350
rect 93554 40294 93622 40350
rect 93678 40294 111250 40350
rect 111306 40294 111374 40350
rect 111430 40294 111498 40350
rect 111554 40294 111622 40350
rect 111678 40294 129250 40350
rect 129306 40294 129374 40350
rect 129430 40294 129498 40350
rect 129554 40294 129622 40350
rect 129678 40294 147250 40350
rect 147306 40294 147374 40350
rect 147430 40294 147498 40350
rect 147554 40294 147622 40350
rect 147678 40294 165250 40350
rect 165306 40294 165374 40350
rect 165430 40294 165498 40350
rect 165554 40294 165622 40350
rect 165678 40294 183250 40350
rect 183306 40294 183374 40350
rect 183430 40294 183498 40350
rect 183554 40294 183622 40350
rect 183678 40294 201250 40350
rect 201306 40294 201374 40350
rect 201430 40294 201498 40350
rect 201554 40294 201622 40350
rect 201678 40294 219250 40350
rect 219306 40294 219374 40350
rect 219430 40294 219498 40350
rect 219554 40294 219622 40350
rect 219678 40294 237250 40350
rect 237306 40294 237374 40350
rect 237430 40294 237498 40350
rect 237554 40294 237622 40350
rect 237678 40294 255250 40350
rect 255306 40294 255374 40350
rect 255430 40294 255498 40350
rect 255554 40294 255622 40350
rect 255678 40294 273250 40350
rect 273306 40294 273374 40350
rect 273430 40294 273498 40350
rect 273554 40294 273622 40350
rect 273678 40294 291250 40350
rect 291306 40294 291374 40350
rect 291430 40294 291498 40350
rect 291554 40294 291622 40350
rect 291678 40294 309250 40350
rect 309306 40294 309374 40350
rect 309430 40294 309498 40350
rect 309554 40294 309622 40350
rect 309678 40294 327250 40350
rect 327306 40294 327374 40350
rect 327430 40294 327498 40350
rect 327554 40294 327622 40350
rect 327678 40294 345250 40350
rect 345306 40294 345374 40350
rect 345430 40294 345498 40350
rect 345554 40294 345622 40350
rect 345678 40294 363250 40350
rect 363306 40294 363374 40350
rect 363430 40294 363498 40350
rect 363554 40294 363622 40350
rect 363678 40294 381250 40350
rect 381306 40294 381374 40350
rect 381430 40294 381498 40350
rect 381554 40294 381622 40350
rect 381678 40294 399250 40350
rect 399306 40294 399374 40350
rect 399430 40294 399498 40350
rect 399554 40294 399622 40350
rect 399678 40294 417250 40350
rect 417306 40294 417374 40350
rect 417430 40294 417498 40350
rect 417554 40294 417622 40350
rect 417678 40294 435250 40350
rect 435306 40294 435374 40350
rect 435430 40294 435498 40350
rect 435554 40294 435622 40350
rect 435678 40294 453250 40350
rect 453306 40294 453374 40350
rect 453430 40294 453498 40350
rect 453554 40294 453622 40350
rect 453678 40294 471250 40350
rect 471306 40294 471374 40350
rect 471430 40294 471498 40350
rect 471554 40294 471622 40350
rect 471678 40294 489250 40350
rect 489306 40294 489374 40350
rect 489430 40294 489498 40350
rect 489554 40294 489622 40350
rect 489678 40294 507250 40350
rect 507306 40294 507374 40350
rect 507430 40294 507498 40350
rect 507554 40294 507622 40350
rect 507678 40294 525250 40350
rect 525306 40294 525374 40350
rect 525430 40294 525498 40350
rect 525554 40294 525622 40350
rect 525678 40294 543250 40350
rect 543306 40294 543374 40350
rect 543430 40294 543498 40350
rect 543554 40294 543622 40350
rect 543678 40294 561250 40350
rect 561306 40294 561374 40350
rect 561430 40294 561498 40350
rect 561554 40294 561622 40350
rect 561678 40294 579250 40350
rect 579306 40294 579374 40350
rect 579430 40294 579498 40350
rect 579554 40294 579622 40350
rect 579678 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 3250 40226
rect 3306 40170 3374 40226
rect 3430 40170 3498 40226
rect 3554 40170 3622 40226
rect 3678 40170 21250 40226
rect 21306 40170 21374 40226
rect 21430 40170 21498 40226
rect 21554 40170 21622 40226
rect 21678 40170 39250 40226
rect 39306 40170 39374 40226
rect 39430 40170 39498 40226
rect 39554 40170 39622 40226
rect 39678 40170 57250 40226
rect 57306 40170 57374 40226
rect 57430 40170 57498 40226
rect 57554 40170 57622 40226
rect 57678 40170 75250 40226
rect 75306 40170 75374 40226
rect 75430 40170 75498 40226
rect 75554 40170 75622 40226
rect 75678 40170 93250 40226
rect 93306 40170 93374 40226
rect 93430 40170 93498 40226
rect 93554 40170 93622 40226
rect 93678 40170 111250 40226
rect 111306 40170 111374 40226
rect 111430 40170 111498 40226
rect 111554 40170 111622 40226
rect 111678 40170 129250 40226
rect 129306 40170 129374 40226
rect 129430 40170 129498 40226
rect 129554 40170 129622 40226
rect 129678 40170 147250 40226
rect 147306 40170 147374 40226
rect 147430 40170 147498 40226
rect 147554 40170 147622 40226
rect 147678 40170 165250 40226
rect 165306 40170 165374 40226
rect 165430 40170 165498 40226
rect 165554 40170 165622 40226
rect 165678 40170 183250 40226
rect 183306 40170 183374 40226
rect 183430 40170 183498 40226
rect 183554 40170 183622 40226
rect 183678 40170 201250 40226
rect 201306 40170 201374 40226
rect 201430 40170 201498 40226
rect 201554 40170 201622 40226
rect 201678 40170 219250 40226
rect 219306 40170 219374 40226
rect 219430 40170 219498 40226
rect 219554 40170 219622 40226
rect 219678 40170 237250 40226
rect 237306 40170 237374 40226
rect 237430 40170 237498 40226
rect 237554 40170 237622 40226
rect 237678 40170 255250 40226
rect 255306 40170 255374 40226
rect 255430 40170 255498 40226
rect 255554 40170 255622 40226
rect 255678 40170 273250 40226
rect 273306 40170 273374 40226
rect 273430 40170 273498 40226
rect 273554 40170 273622 40226
rect 273678 40170 291250 40226
rect 291306 40170 291374 40226
rect 291430 40170 291498 40226
rect 291554 40170 291622 40226
rect 291678 40170 309250 40226
rect 309306 40170 309374 40226
rect 309430 40170 309498 40226
rect 309554 40170 309622 40226
rect 309678 40170 327250 40226
rect 327306 40170 327374 40226
rect 327430 40170 327498 40226
rect 327554 40170 327622 40226
rect 327678 40170 345250 40226
rect 345306 40170 345374 40226
rect 345430 40170 345498 40226
rect 345554 40170 345622 40226
rect 345678 40170 363250 40226
rect 363306 40170 363374 40226
rect 363430 40170 363498 40226
rect 363554 40170 363622 40226
rect 363678 40170 381250 40226
rect 381306 40170 381374 40226
rect 381430 40170 381498 40226
rect 381554 40170 381622 40226
rect 381678 40170 399250 40226
rect 399306 40170 399374 40226
rect 399430 40170 399498 40226
rect 399554 40170 399622 40226
rect 399678 40170 417250 40226
rect 417306 40170 417374 40226
rect 417430 40170 417498 40226
rect 417554 40170 417622 40226
rect 417678 40170 435250 40226
rect 435306 40170 435374 40226
rect 435430 40170 435498 40226
rect 435554 40170 435622 40226
rect 435678 40170 453250 40226
rect 453306 40170 453374 40226
rect 453430 40170 453498 40226
rect 453554 40170 453622 40226
rect 453678 40170 471250 40226
rect 471306 40170 471374 40226
rect 471430 40170 471498 40226
rect 471554 40170 471622 40226
rect 471678 40170 489250 40226
rect 489306 40170 489374 40226
rect 489430 40170 489498 40226
rect 489554 40170 489622 40226
rect 489678 40170 507250 40226
rect 507306 40170 507374 40226
rect 507430 40170 507498 40226
rect 507554 40170 507622 40226
rect 507678 40170 525250 40226
rect 525306 40170 525374 40226
rect 525430 40170 525498 40226
rect 525554 40170 525622 40226
rect 525678 40170 543250 40226
rect 543306 40170 543374 40226
rect 543430 40170 543498 40226
rect 543554 40170 543622 40226
rect 543678 40170 561250 40226
rect 561306 40170 561374 40226
rect 561430 40170 561498 40226
rect 561554 40170 561622 40226
rect 561678 40170 579250 40226
rect 579306 40170 579374 40226
rect 579430 40170 579498 40226
rect 579554 40170 579622 40226
rect 579678 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 3250 40102
rect 3306 40046 3374 40102
rect 3430 40046 3498 40102
rect 3554 40046 3622 40102
rect 3678 40046 21250 40102
rect 21306 40046 21374 40102
rect 21430 40046 21498 40102
rect 21554 40046 21622 40102
rect 21678 40046 39250 40102
rect 39306 40046 39374 40102
rect 39430 40046 39498 40102
rect 39554 40046 39622 40102
rect 39678 40046 57250 40102
rect 57306 40046 57374 40102
rect 57430 40046 57498 40102
rect 57554 40046 57622 40102
rect 57678 40046 75250 40102
rect 75306 40046 75374 40102
rect 75430 40046 75498 40102
rect 75554 40046 75622 40102
rect 75678 40046 93250 40102
rect 93306 40046 93374 40102
rect 93430 40046 93498 40102
rect 93554 40046 93622 40102
rect 93678 40046 111250 40102
rect 111306 40046 111374 40102
rect 111430 40046 111498 40102
rect 111554 40046 111622 40102
rect 111678 40046 129250 40102
rect 129306 40046 129374 40102
rect 129430 40046 129498 40102
rect 129554 40046 129622 40102
rect 129678 40046 147250 40102
rect 147306 40046 147374 40102
rect 147430 40046 147498 40102
rect 147554 40046 147622 40102
rect 147678 40046 165250 40102
rect 165306 40046 165374 40102
rect 165430 40046 165498 40102
rect 165554 40046 165622 40102
rect 165678 40046 183250 40102
rect 183306 40046 183374 40102
rect 183430 40046 183498 40102
rect 183554 40046 183622 40102
rect 183678 40046 201250 40102
rect 201306 40046 201374 40102
rect 201430 40046 201498 40102
rect 201554 40046 201622 40102
rect 201678 40046 219250 40102
rect 219306 40046 219374 40102
rect 219430 40046 219498 40102
rect 219554 40046 219622 40102
rect 219678 40046 237250 40102
rect 237306 40046 237374 40102
rect 237430 40046 237498 40102
rect 237554 40046 237622 40102
rect 237678 40046 255250 40102
rect 255306 40046 255374 40102
rect 255430 40046 255498 40102
rect 255554 40046 255622 40102
rect 255678 40046 273250 40102
rect 273306 40046 273374 40102
rect 273430 40046 273498 40102
rect 273554 40046 273622 40102
rect 273678 40046 291250 40102
rect 291306 40046 291374 40102
rect 291430 40046 291498 40102
rect 291554 40046 291622 40102
rect 291678 40046 309250 40102
rect 309306 40046 309374 40102
rect 309430 40046 309498 40102
rect 309554 40046 309622 40102
rect 309678 40046 327250 40102
rect 327306 40046 327374 40102
rect 327430 40046 327498 40102
rect 327554 40046 327622 40102
rect 327678 40046 345250 40102
rect 345306 40046 345374 40102
rect 345430 40046 345498 40102
rect 345554 40046 345622 40102
rect 345678 40046 363250 40102
rect 363306 40046 363374 40102
rect 363430 40046 363498 40102
rect 363554 40046 363622 40102
rect 363678 40046 381250 40102
rect 381306 40046 381374 40102
rect 381430 40046 381498 40102
rect 381554 40046 381622 40102
rect 381678 40046 399250 40102
rect 399306 40046 399374 40102
rect 399430 40046 399498 40102
rect 399554 40046 399622 40102
rect 399678 40046 417250 40102
rect 417306 40046 417374 40102
rect 417430 40046 417498 40102
rect 417554 40046 417622 40102
rect 417678 40046 435250 40102
rect 435306 40046 435374 40102
rect 435430 40046 435498 40102
rect 435554 40046 435622 40102
rect 435678 40046 453250 40102
rect 453306 40046 453374 40102
rect 453430 40046 453498 40102
rect 453554 40046 453622 40102
rect 453678 40046 471250 40102
rect 471306 40046 471374 40102
rect 471430 40046 471498 40102
rect 471554 40046 471622 40102
rect 471678 40046 489250 40102
rect 489306 40046 489374 40102
rect 489430 40046 489498 40102
rect 489554 40046 489622 40102
rect 489678 40046 507250 40102
rect 507306 40046 507374 40102
rect 507430 40046 507498 40102
rect 507554 40046 507622 40102
rect 507678 40046 525250 40102
rect 525306 40046 525374 40102
rect 525430 40046 525498 40102
rect 525554 40046 525622 40102
rect 525678 40046 543250 40102
rect 543306 40046 543374 40102
rect 543430 40046 543498 40102
rect 543554 40046 543622 40102
rect 543678 40046 561250 40102
rect 561306 40046 561374 40102
rect 561430 40046 561498 40102
rect 561554 40046 561622 40102
rect 561678 40046 579250 40102
rect 579306 40046 579374 40102
rect 579430 40046 579498 40102
rect 579554 40046 579622 40102
rect 579678 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 3250 39978
rect 3306 39922 3374 39978
rect 3430 39922 3498 39978
rect 3554 39922 3622 39978
rect 3678 39922 21250 39978
rect 21306 39922 21374 39978
rect 21430 39922 21498 39978
rect 21554 39922 21622 39978
rect 21678 39922 39250 39978
rect 39306 39922 39374 39978
rect 39430 39922 39498 39978
rect 39554 39922 39622 39978
rect 39678 39922 57250 39978
rect 57306 39922 57374 39978
rect 57430 39922 57498 39978
rect 57554 39922 57622 39978
rect 57678 39922 75250 39978
rect 75306 39922 75374 39978
rect 75430 39922 75498 39978
rect 75554 39922 75622 39978
rect 75678 39922 93250 39978
rect 93306 39922 93374 39978
rect 93430 39922 93498 39978
rect 93554 39922 93622 39978
rect 93678 39922 111250 39978
rect 111306 39922 111374 39978
rect 111430 39922 111498 39978
rect 111554 39922 111622 39978
rect 111678 39922 129250 39978
rect 129306 39922 129374 39978
rect 129430 39922 129498 39978
rect 129554 39922 129622 39978
rect 129678 39922 147250 39978
rect 147306 39922 147374 39978
rect 147430 39922 147498 39978
rect 147554 39922 147622 39978
rect 147678 39922 165250 39978
rect 165306 39922 165374 39978
rect 165430 39922 165498 39978
rect 165554 39922 165622 39978
rect 165678 39922 183250 39978
rect 183306 39922 183374 39978
rect 183430 39922 183498 39978
rect 183554 39922 183622 39978
rect 183678 39922 201250 39978
rect 201306 39922 201374 39978
rect 201430 39922 201498 39978
rect 201554 39922 201622 39978
rect 201678 39922 219250 39978
rect 219306 39922 219374 39978
rect 219430 39922 219498 39978
rect 219554 39922 219622 39978
rect 219678 39922 237250 39978
rect 237306 39922 237374 39978
rect 237430 39922 237498 39978
rect 237554 39922 237622 39978
rect 237678 39922 255250 39978
rect 255306 39922 255374 39978
rect 255430 39922 255498 39978
rect 255554 39922 255622 39978
rect 255678 39922 273250 39978
rect 273306 39922 273374 39978
rect 273430 39922 273498 39978
rect 273554 39922 273622 39978
rect 273678 39922 291250 39978
rect 291306 39922 291374 39978
rect 291430 39922 291498 39978
rect 291554 39922 291622 39978
rect 291678 39922 309250 39978
rect 309306 39922 309374 39978
rect 309430 39922 309498 39978
rect 309554 39922 309622 39978
rect 309678 39922 327250 39978
rect 327306 39922 327374 39978
rect 327430 39922 327498 39978
rect 327554 39922 327622 39978
rect 327678 39922 345250 39978
rect 345306 39922 345374 39978
rect 345430 39922 345498 39978
rect 345554 39922 345622 39978
rect 345678 39922 363250 39978
rect 363306 39922 363374 39978
rect 363430 39922 363498 39978
rect 363554 39922 363622 39978
rect 363678 39922 381250 39978
rect 381306 39922 381374 39978
rect 381430 39922 381498 39978
rect 381554 39922 381622 39978
rect 381678 39922 399250 39978
rect 399306 39922 399374 39978
rect 399430 39922 399498 39978
rect 399554 39922 399622 39978
rect 399678 39922 417250 39978
rect 417306 39922 417374 39978
rect 417430 39922 417498 39978
rect 417554 39922 417622 39978
rect 417678 39922 435250 39978
rect 435306 39922 435374 39978
rect 435430 39922 435498 39978
rect 435554 39922 435622 39978
rect 435678 39922 453250 39978
rect 453306 39922 453374 39978
rect 453430 39922 453498 39978
rect 453554 39922 453622 39978
rect 453678 39922 471250 39978
rect 471306 39922 471374 39978
rect 471430 39922 471498 39978
rect 471554 39922 471622 39978
rect 471678 39922 489250 39978
rect 489306 39922 489374 39978
rect 489430 39922 489498 39978
rect 489554 39922 489622 39978
rect 489678 39922 507250 39978
rect 507306 39922 507374 39978
rect 507430 39922 507498 39978
rect 507554 39922 507622 39978
rect 507678 39922 525250 39978
rect 525306 39922 525374 39978
rect 525430 39922 525498 39978
rect 525554 39922 525622 39978
rect 525678 39922 543250 39978
rect 543306 39922 543374 39978
rect 543430 39922 543498 39978
rect 543554 39922 543622 39978
rect 543678 39922 561250 39978
rect 561306 39922 561374 39978
rect 561430 39922 561498 39978
rect 561554 39922 561622 39978
rect 561678 39922 579250 39978
rect 579306 39922 579374 39978
rect 579430 39922 579498 39978
rect 579554 39922 579622 39978
rect 579678 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 6970 28350
rect 7026 28294 7094 28350
rect 7150 28294 7218 28350
rect 7274 28294 7342 28350
rect 7398 28294 24970 28350
rect 25026 28294 25094 28350
rect 25150 28294 25218 28350
rect 25274 28294 25342 28350
rect 25398 28294 42970 28350
rect 43026 28294 43094 28350
rect 43150 28294 43218 28350
rect 43274 28294 43342 28350
rect 43398 28294 60970 28350
rect 61026 28294 61094 28350
rect 61150 28294 61218 28350
rect 61274 28294 61342 28350
rect 61398 28294 78970 28350
rect 79026 28294 79094 28350
rect 79150 28294 79218 28350
rect 79274 28294 79342 28350
rect 79398 28294 96970 28350
rect 97026 28294 97094 28350
rect 97150 28294 97218 28350
rect 97274 28294 97342 28350
rect 97398 28294 114970 28350
rect 115026 28294 115094 28350
rect 115150 28294 115218 28350
rect 115274 28294 115342 28350
rect 115398 28294 132970 28350
rect 133026 28294 133094 28350
rect 133150 28294 133218 28350
rect 133274 28294 133342 28350
rect 133398 28294 150970 28350
rect 151026 28294 151094 28350
rect 151150 28294 151218 28350
rect 151274 28294 151342 28350
rect 151398 28294 168970 28350
rect 169026 28294 169094 28350
rect 169150 28294 169218 28350
rect 169274 28294 169342 28350
rect 169398 28294 186970 28350
rect 187026 28294 187094 28350
rect 187150 28294 187218 28350
rect 187274 28294 187342 28350
rect 187398 28294 204970 28350
rect 205026 28294 205094 28350
rect 205150 28294 205218 28350
rect 205274 28294 205342 28350
rect 205398 28294 222970 28350
rect 223026 28294 223094 28350
rect 223150 28294 223218 28350
rect 223274 28294 223342 28350
rect 223398 28294 240970 28350
rect 241026 28294 241094 28350
rect 241150 28294 241218 28350
rect 241274 28294 241342 28350
rect 241398 28294 258970 28350
rect 259026 28294 259094 28350
rect 259150 28294 259218 28350
rect 259274 28294 259342 28350
rect 259398 28294 276970 28350
rect 277026 28294 277094 28350
rect 277150 28294 277218 28350
rect 277274 28294 277342 28350
rect 277398 28294 294970 28350
rect 295026 28294 295094 28350
rect 295150 28294 295218 28350
rect 295274 28294 295342 28350
rect 295398 28294 312970 28350
rect 313026 28294 313094 28350
rect 313150 28294 313218 28350
rect 313274 28294 313342 28350
rect 313398 28294 330970 28350
rect 331026 28294 331094 28350
rect 331150 28294 331218 28350
rect 331274 28294 331342 28350
rect 331398 28294 348970 28350
rect 349026 28294 349094 28350
rect 349150 28294 349218 28350
rect 349274 28294 349342 28350
rect 349398 28294 366970 28350
rect 367026 28294 367094 28350
rect 367150 28294 367218 28350
rect 367274 28294 367342 28350
rect 367398 28294 384970 28350
rect 385026 28294 385094 28350
rect 385150 28294 385218 28350
rect 385274 28294 385342 28350
rect 385398 28294 402970 28350
rect 403026 28294 403094 28350
rect 403150 28294 403218 28350
rect 403274 28294 403342 28350
rect 403398 28294 420970 28350
rect 421026 28294 421094 28350
rect 421150 28294 421218 28350
rect 421274 28294 421342 28350
rect 421398 28294 438970 28350
rect 439026 28294 439094 28350
rect 439150 28294 439218 28350
rect 439274 28294 439342 28350
rect 439398 28294 456970 28350
rect 457026 28294 457094 28350
rect 457150 28294 457218 28350
rect 457274 28294 457342 28350
rect 457398 28294 474970 28350
rect 475026 28294 475094 28350
rect 475150 28294 475218 28350
rect 475274 28294 475342 28350
rect 475398 28294 492970 28350
rect 493026 28294 493094 28350
rect 493150 28294 493218 28350
rect 493274 28294 493342 28350
rect 493398 28294 510970 28350
rect 511026 28294 511094 28350
rect 511150 28294 511218 28350
rect 511274 28294 511342 28350
rect 511398 28294 528970 28350
rect 529026 28294 529094 28350
rect 529150 28294 529218 28350
rect 529274 28294 529342 28350
rect 529398 28294 546970 28350
rect 547026 28294 547094 28350
rect 547150 28294 547218 28350
rect 547274 28294 547342 28350
rect 547398 28294 564970 28350
rect 565026 28294 565094 28350
rect 565150 28294 565218 28350
rect 565274 28294 565342 28350
rect 565398 28294 582970 28350
rect 583026 28294 583094 28350
rect 583150 28294 583218 28350
rect 583274 28294 583342 28350
rect 583398 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 6970 28226
rect 7026 28170 7094 28226
rect 7150 28170 7218 28226
rect 7274 28170 7342 28226
rect 7398 28170 24970 28226
rect 25026 28170 25094 28226
rect 25150 28170 25218 28226
rect 25274 28170 25342 28226
rect 25398 28170 42970 28226
rect 43026 28170 43094 28226
rect 43150 28170 43218 28226
rect 43274 28170 43342 28226
rect 43398 28170 60970 28226
rect 61026 28170 61094 28226
rect 61150 28170 61218 28226
rect 61274 28170 61342 28226
rect 61398 28170 78970 28226
rect 79026 28170 79094 28226
rect 79150 28170 79218 28226
rect 79274 28170 79342 28226
rect 79398 28170 96970 28226
rect 97026 28170 97094 28226
rect 97150 28170 97218 28226
rect 97274 28170 97342 28226
rect 97398 28170 114970 28226
rect 115026 28170 115094 28226
rect 115150 28170 115218 28226
rect 115274 28170 115342 28226
rect 115398 28170 132970 28226
rect 133026 28170 133094 28226
rect 133150 28170 133218 28226
rect 133274 28170 133342 28226
rect 133398 28170 150970 28226
rect 151026 28170 151094 28226
rect 151150 28170 151218 28226
rect 151274 28170 151342 28226
rect 151398 28170 168970 28226
rect 169026 28170 169094 28226
rect 169150 28170 169218 28226
rect 169274 28170 169342 28226
rect 169398 28170 186970 28226
rect 187026 28170 187094 28226
rect 187150 28170 187218 28226
rect 187274 28170 187342 28226
rect 187398 28170 204970 28226
rect 205026 28170 205094 28226
rect 205150 28170 205218 28226
rect 205274 28170 205342 28226
rect 205398 28170 222970 28226
rect 223026 28170 223094 28226
rect 223150 28170 223218 28226
rect 223274 28170 223342 28226
rect 223398 28170 240970 28226
rect 241026 28170 241094 28226
rect 241150 28170 241218 28226
rect 241274 28170 241342 28226
rect 241398 28170 258970 28226
rect 259026 28170 259094 28226
rect 259150 28170 259218 28226
rect 259274 28170 259342 28226
rect 259398 28170 276970 28226
rect 277026 28170 277094 28226
rect 277150 28170 277218 28226
rect 277274 28170 277342 28226
rect 277398 28170 294970 28226
rect 295026 28170 295094 28226
rect 295150 28170 295218 28226
rect 295274 28170 295342 28226
rect 295398 28170 312970 28226
rect 313026 28170 313094 28226
rect 313150 28170 313218 28226
rect 313274 28170 313342 28226
rect 313398 28170 330970 28226
rect 331026 28170 331094 28226
rect 331150 28170 331218 28226
rect 331274 28170 331342 28226
rect 331398 28170 348970 28226
rect 349026 28170 349094 28226
rect 349150 28170 349218 28226
rect 349274 28170 349342 28226
rect 349398 28170 366970 28226
rect 367026 28170 367094 28226
rect 367150 28170 367218 28226
rect 367274 28170 367342 28226
rect 367398 28170 384970 28226
rect 385026 28170 385094 28226
rect 385150 28170 385218 28226
rect 385274 28170 385342 28226
rect 385398 28170 402970 28226
rect 403026 28170 403094 28226
rect 403150 28170 403218 28226
rect 403274 28170 403342 28226
rect 403398 28170 420970 28226
rect 421026 28170 421094 28226
rect 421150 28170 421218 28226
rect 421274 28170 421342 28226
rect 421398 28170 438970 28226
rect 439026 28170 439094 28226
rect 439150 28170 439218 28226
rect 439274 28170 439342 28226
rect 439398 28170 456970 28226
rect 457026 28170 457094 28226
rect 457150 28170 457218 28226
rect 457274 28170 457342 28226
rect 457398 28170 474970 28226
rect 475026 28170 475094 28226
rect 475150 28170 475218 28226
rect 475274 28170 475342 28226
rect 475398 28170 492970 28226
rect 493026 28170 493094 28226
rect 493150 28170 493218 28226
rect 493274 28170 493342 28226
rect 493398 28170 510970 28226
rect 511026 28170 511094 28226
rect 511150 28170 511218 28226
rect 511274 28170 511342 28226
rect 511398 28170 528970 28226
rect 529026 28170 529094 28226
rect 529150 28170 529218 28226
rect 529274 28170 529342 28226
rect 529398 28170 546970 28226
rect 547026 28170 547094 28226
rect 547150 28170 547218 28226
rect 547274 28170 547342 28226
rect 547398 28170 564970 28226
rect 565026 28170 565094 28226
rect 565150 28170 565218 28226
rect 565274 28170 565342 28226
rect 565398 28170 582970 28226
rect 583026 28170 583094 28226
rect 583150 28170 583218 28226
rect 583274 28170 583342 28226
rect 583398 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 6970 28102
rect 7026 28046 7094 28102
rect 7150 28046 7218 28102
rect 7274 28046 7342 28102
rect 7398 28046 24970 28102
rect 25026 28046 25094 28102
rect 25150 28046 25218 28102
rect 25274 28046 25342 28102
rect 25398 28046 42970 28102
rect 43026 28046 43094 28102
rect 43150 28046 43218 28102
rect 43274 28046 43342 28102
rect 43398 28046 60970 28102
rect 61026 28046 61094 28102
rect 61150 28046 61218 28102
rect 61274 28046 61342 28102
rect 61398 28046 78970 28102
rect 79026 28046 79094 28102
rect 79150 28046 79218 28102
rect 79274 28046 79342 28102
rect 79398 28046 96970 28102
rect 97026 28046 97094 28102
rect 97150 28046 97218 28102
rect 97274 28046 97342 28102
rect 97398 28046 114970 28102
rect 115026 28046 115094 28102
rect 115150 28046 115218 28102
rect 115274 28046 115342 28102
rect 115398 28046 132970 28102
rect 133026 28046 133094 28102
rect 133150 28046 133218 28102
rect 133274 28046 133342 28102
rect 133398 28046 150970 28102
rect 151026 28046 151094 28102
rect 151150 28046 151218 28102
rect 151274 28046 151342 28102
rect 151398 28046 168970 28102
rect 169026 28046 169094 28102
rect 169150 28046 169218 28102
rect 169274 28046 169342 28102
rect 169398 28046 186970 28102
rect 187026 28046 187094 28102
rect 187150 28046 187218 28102
rect 187274 28046 187342 28102
rect 187398 28046 204970 28102
rect 205026 28046 205094 28102
rect 205150 28046 205218 28102
rect 205274 28046 205342 28102
rect 205398 28046 222970 28102
rect 223026 28046 223094 28102
rect 223150 28046 223218 28102
rect 223274 28046 223342 28102
rect 223398 28046 240970 28102
rect 241026 28046 241094 28102
rect 241150 28046 241218 28102
rect 241274 28046 241342 28102
rect 241398 28046 258970 28102
rect 259026 28046 259094 28102
rect 259150 28046 259218 28102
rect 259274 28046 259342 28102
rect 259398 28046 276970 28102
rect 277026 28046 277094 28102
rect 277150 28046 277218 28102
rect 277274 28046 277342 28102
rect 277398 28046 294970 28102
rect 295026 28046 295094 28102
rect 295150 28046 295218 28102
rect 295274 28046 295342 28102
rect 295398 28046 312970 28102
rect 313026 28046 313094 28102
rect 313150 28046 313218 28102
rect 313274 28046 313342 28102
rect 313398 28046 330970 28102
rect 331026 28046 331094 28102
rect 331150 28046 331218 28102
rect 331274 28046 331342 28102
rect 331398 28046 348970 28102
rect 349026 28046 349094 28102
rect 349150 28046 349218 28102
rect 349274 28046 349342 28102
rect 349398 28046 366970 28102
rect 367026 28046 367094 28102
rect 367150 28046 367218 28102
rect 367274 28046 367342 28102
rect 367398 28046 384970 28102
rect 385026 28046 385094 28102
rect 385150 28046 385218 28102
rect 385274 28046 385342 28102
rect 385398 28046 402970 28102
rect 403026 28046 403094 28102
rect 403150 28046 403218 28102
rect 403274 28046 403342 28102
rect 403398 28046 420970 28102
rect 421026 28046 421094 28102
rect 421150 28046 421218 28102
rect 421274 28046 421342 28102
rect 421398 28046 438970 28102
rect 439026 28046 439094 28102
rect 439150 28046 439218 28102
rect 439274 28046 439342 28102
rect 439398 28046 456970 28102
rect 457026 28046 457094 28102
rect 457150 28046 457218 28102
rect 457274 28046 457342 28102
rect 457398 28046 474970 28102
rect 475026 28046 475094 28102
rect 475150 28046 475218 28102
rect 475274 28046 475342 28102
rect 475398 28046 492970 28102
rect 493026 28046 493094 28102
rect 493150 28046 493218 28102
rect 493274 28046 493342 28102
rect 493398 28046 510970 28102
rect 511026 28046 511094 28102
rect 511150 28046 511218 28102
rect 511274 28046 511342 28102
rect 511398 28046 528970 28102
rect 529026 28046 529094 28102
rect 529150 28046 529218 28102
rect 529274 28046 529342 28102
rect 529398 28046 546970 28102
rect 547026 28046 547094 28102
rect 547150 28046 547218 28102
rect 547274 28046 547342 28102
rect 547398 28046 564970 28102
rect 565026 28046 565094 28102
rect 565150 28046 565218 28102
rect 565274 28046 565342 28102
rect 565398 28046 582970 28102
rect 583026 28046 583094 28102
rect 583150 28046 583218 28102
rect 583274 28046 583342 28102
rect 583398 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 6970 27978
rect 7026 27922 7094 27978
rect 7150 27922 7218 27978
rect 7274 27922 7342 27978
rect 7398 27922 24970 27978
rect 25026 27922 25094 27978
rect 25150 27922 25218 27978
rect 25274 27922 25342 27978
rect 25398 27922 42970 27978
rect 43026 27922 43094 27978
rect 43150 27922 43218 27978
rect 43274 27922 43342 27978
rect 43398 27922 60970 27978
rect 61026 27922 61094 27978
rect 61150 27922 61218 27978
rect 61274 27922 61342 27978
rect 61398 27922 78970 27978
rect 79026 27922 79094 27978
rect 79150 27922 79218 27978
rect 79274 27922 79342 27978
rect 79398 27922 96970 27978
rect 97026 27922 97094 27978
rect 97150 27922 97218 27978
rect 97274 27922 97342 27978
rect 97398 27922 114970 27978
rect 115026 27922 115094 27978
rect 115150 27922 115218 27978
rect 115274 27922 115342 27978
rect 115398 27922 132970 27978
rect 133026 27922 133094 27978
rect 133150 27922 133218 27978
rect 133274 27922 133342 27978
rect 133398 27922 150970 27978
rect 151026 27922 151094 27978
rect 151150 27922 151218 27978
rect 151274 27922 151342 27978
rect 151398 27922 168970 27978
rect 169026 27922 169094 27978
rect 169150 27922 169218 27978
rect 169274 27922 169342 27978
rect 169398 27922 186970 27978
rect 187026 27922 187094 27978
rect 187150 27922 187218 27978
rect 187274 27922 187342 27978
rect 187398 27922 204970 27978
rect 205026 27922 205094 27978
rect 205150 27922 205218 27978
rect 205274 27922 205342 27978
rect 205398 27922 222970 27978
rect 223026 27922 223094 27978
rect 223150 27922 223218 27978
rect 223274 27922 223342 27978
rect 223398 27922 240970 27978
rect 241026 27922 241094 27978
rect 241150 27922 241218 27978
rect 241274 27922 241342 27978
rect 241398 27922 258970 27978
rect 259026 27922 259094 27978
rect 259150 27922 259218 27978
rect 259274 27922 259342 27978
rect 259398 27922 276970 27978
rect 277026 27922 277094 27978
rect 277150 27922 277218 27978
rect 277274 27922 277342 27978
rect 277398 27922 294970 27978
rect 295026 27922 295094 27978
rect 295150 27922 295218 27978
rect 295274 27922 295342 27978
rect 295398 27922 312970 27978
rect 313026 27922 313094 27978
rect 313150 27922 313218 27978
rect 313274 27922 313342 27978
rect 313398 27922 330970 27978
rect 331026 27922 331094 27978
rect 331150 27922 331218 27978
rect 331274 27922 331342 27978
rect 331398 27922 348970 27978
rect 349026 27922 349094 27978
rect 349150 27922 349218 27978
rect 349274 27922 349342 27978
rect 349398 27922 366970 27978
rect 367026 27922 367094 27978
rect 367150 27922 367218 27978
rect 367274 27922 367342 27978
rect 367398 27922 384970 27978
rect 385026 27922 385094 27978
rect 385150 27922 385218 27978
rect 385274 27922 385342 27978
rect 385398 27922 402970 27978
rect 403026 27922 403094 27978
rect 403150 27922 403218 27978
rect 403274 27922 403342 27978
rect 403398 27922 420970 27978
rect 421026 27922 421094 27978
rect 421150 27922 421218 27978
rect 421274 27922 421342 27978
rect 421398 27922 438970 27978
rect 439026 27922 439094 27978
rect 439150 27922 439218 27978
rect 439274 27922 439342 27978
rect 439398 27922 456970 27978
rect 457026 27922 457094 27978
rect 457150 27922 457218 27978
rect 457274 27922 457342 27978
rect 457398 27922 474970 27978
rect 475026 27922 475094 27978
rect 475150 27922 475218 27978
rect 475274 27922 475342 27978
rect 475398 27922 492970 27978
rect 493026 27922 493094 27978
rect 493150 27922 493218 27978
rect 493274 27922 493342 27978
rect 493398 27922 510970 27978
rect 511026 27922 511094 27978
rect 511150 27922 511218 27978
rect 511274 27922 511342 27978
rect 511398 27922 528970 27978
rect 529026 27922 529094 27978
rect 529150 27922 529218 27978
rect 529274 27922 529342 27978
rect 529398 27922 546970 27978
rect 547026 27922 547094 27978
rect 547150 27922 547218 27978
rect 547274 27922 547342 27978
rect 547398 27922 564970 27978
rect 565026 27922 565094 27978
rect 565150 27922 565218 27978
rect 565274 27922 565342 27978
rect 565398 27922 582970 27978
rect 583026 27922 583094 27978
rect 583150 27922 583218 27978
rect 583274 27922 583342 27978
rect 583398 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 3250 22350
rect 3306 22294 3374 22350
rect 3430 22294 3498 22350
rect 3554 22294 3622 22350
rect 3678 22294 21250 22350
rect 21306 22294 21374 22350
rect 21430 22294 21498 22350
rect 21554 22294 21622 22350
rect 21678 22294 39250 22350
rect 39306 22294 39374 22350
rect 39430 22294 39498 22350
rect 39554 22294 39622 22350
rect 39678 22294 57250 22350
rect 57306 22294 57374 22350
rect 57430 22294 57498 22350
rect 57554 22294 57622 22350
rect 57678 22294 75250 22350
rect 75306 22294 75374 22350
rect 75430 22294 75498 22350
rect 75554 22294 75622 22350
rect 75678 22294 93250 22350
rect 93306 22294 93374 22350
rect 93430 22294 93498 22350
rect 93554 22294 93622 22350
rect 93678 22294 111250 22350
rect 111306 22294 111374 22350
rect 111430 22294 111498 22350
rect 111554 22294 111622 22350
rect 111678 22294 129250 22350
rect 129306 22294 129374 22350
rect 129430 22294 129498 22350
rect 129554 22294 129622 22350
rect 129678 22294 147250 22350
rect 147306 22294 147374 22350
rect 147430 22294 147498 22350
rect 147554 22294 147622 22350
rect 147678 22294 165250 22350
rect 165306 22294 165374 22350
rect 165430 22294 165498 22350
rect 165554 22294 165622 22350
rect 165678 22294 183250 22350
rect 183306 22294 183374 22350
rect 183430 22294 183498 22350
rect 183554 22294 183622 22350
rect 183678 22294 201250 22350
rect 201306 22294 201374 22350
rect 201430 22294 201498 22350
rect 201554 22294 201622 22350
rect 201678 22294 219250 22350
rect 219306 22294 219374 22350
rect 219430 22294 219498 22350
rect 219554 22294 219622 22350
rect 219678 22294 237250 22350
rect 237306 22294 237374 22350
rect 237430 22294 237498 22350
rect 237554 22294 237622 22350
rect 237678 22294 255250 22350
rect 255306 22294 255374 22350
rect 255430 22294 255498 22350
rect 255554 22294 255622 22350
rect 255678 22294 273250 22350
rect 273306 22294 273374 22350
rect 273430 22294 273498 22350
rect 273554 22294 273622 22350
rect 273678 22294 291250 22350
rect 291306 22294 291374 22350
rect 291430 22294 291498 22350
rect 291554 22294 291622 22350
rect 291678 22294 309250 22350
rect 309306 22294 309374 22350
rect 309430 22294 309498 22350
rect 309554 22294 309622 22350
rect 309678 22294 327250 22350
rect 327306 22294 327374 22350
rect 327430 22294 327498 22350
rect 327554 22294 327622 22350
rect 327678 22294 345250 22350
rect 345306 22294 345374 22350
rect 345430 22294 345498 22350
rect 345554 22294 345622 22350
rect 345678 22294 363250 22350
rect 363306 22294 363374 22350
rect 363430 22294 363498 22350
rect 363554 22294 363622 22350
rect 363678 22294 381250 22350
rect 381306 22294 381374 22350
rect 381430 22294 381498 22350
rect 381554 22294 381622 22350
rect 381678 22294 399250 22350
rect 399306 22294 399374 22350
rect 399430 22294 399498 22350
rect 399554 22294 399622 22350
rect 399678 22294 417250 22350
rect 417306 22294 417374 22350
rect 417430 22294 417498 22350
rect 417554 22294 417622 22350
rect 417678 22294 435250 22350
rect 435306 22294 435374 22350
rect 435430 22294 435498 22350
rect 435554 22294 435622 22350
rect 435678 22294 453250 22350
rect 453306 22294 453374 22350
rect 453430 22294 453498 22350
rect 453554 22294 453622 22350
rect 453678 22294 471250 22350
rect 471306 22294 471374 22350
rect 471430 22294 471498 22350
rect 471554 22294 471622 22350
rect 471678 22294 489250 22350
rect 489306 22294 489374 22350
rect 489430 22294 489498 22350
rect 489554 22294 489622 22350
rect 489678 22294 507250 22350
rect 507306 22294 507374 22350
rect 507430 22294 507498 22350
rect 507554 22294 507622 22350
rect 507678 22294 525250 22350
rect 525306 22294 525374 22350
rect 525430 22294 525498 22350
rect 525554 22294 525622 22350
rect 525678 22294 543250 22350
rect 543306 22294 543374 22350
rect 543430 22294 543498 22350
rect 543554 22294 543622 22350
rect 543678 22294 561250 22350
rect 561306 22294 561374 22350
rect 561430 22294 561498 22350
rect 561554 22294 561622 22350
rect 561678 22294 579250 22350
rect 579306 22294 579374 22350
rect 579430 22294 579498 22350
rect 579554 22294 579622 22350
rect 579678 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 3250 22226
rect 3306 22170 3374 22226
rect 3430 22170 3498 22226
rect 3554 22170 3622 22226
rect 3678 22170 21250 22226
rect 21306 22170 21374 22226
rect 21430 22170 21498 22226
rect 21554 22170 21622 22226
rect 21678 22170 39250 22226
rect 39306 22170 39374 22226
rect 39430 22170 39498 22226
rect 39554 22170 39622 22226
rect 39678 22170 57250 22226
rect 57306 22170 57374 22226
rect 57430 22170 57498 22226
rect 57554 22170 57622 22226
rect 57678 22170 75250 22226
rect 75306 22170 75374 22226
rect 75430 22170 75498 22226
rect 75554 22170 75622 22226
rect 75678 22170 93250 22226
rect 93306 22170 93374 22226
rect 93430 22170 93498 22226
rect 93554 22170 93622 22226
rect 93678 22170 111250 22226
rect 111306 22170 111374 22226
rect 111430 22170 111498 22226
rect 111554 22170 111622 22226
rect 111678 22170 129250 22226
rect 129306 22170 129374 22226
rect 129430 22170 129498 22226
rect 129554 22170 129622 22226
rect 129678 22170 147250 22226
rect 147306 22170 147374 22226
rect 147430 22170 147498 22226
rect 147554 22170 147622 22226
rect 147678 22170 165250 22226
rect 165306 22170 165374 22226
rect 165430 22170 165498 22226
rect 165554 22170 165622 22226
rect 165678 22170 183250 22226
rect 183306 22170 183374 22226
rect 183430 22170 183498 22226
rect 183554 22170 183622 22226
rect 183678 22170 201250 22226
rect 201306 22170 201374 22226
rect 201430 22170 201498 22226
rect 201554 22170 201622 22226
rect 201678 22170 219250 22226
rect 219306 22170 219374 22226
rect 219430 22170 219498 22226
rect 219554 22170 219622 22226
rect 219678 22170 237250 22226
rect 237306 22170 237374 22226
rect 237430 22170 237498 22226
rect 237554 22170 237622 22226
rect 237678 22170 255250 22226
rect 255306 22170 255374 22226
rect 255430 22170 255498 22226
rect 255554 22170 255622 22226
rect 255678 22170 273250 22226
rect 273306 22170 273374 22226
rect 273430 22170 273498 22226
rect 273554 22170 273622 22226
rect 273678 22170 291250 22226
rect 291306 22170 291374 22226
rect 291430 22170 291498 22226
rect 291554 22170 291622 22226
rect 291678 22170 309250 22226
rect 309306 22170 309374 22226
rect 309430 22170 309498 22226
rect 309554 22170 309622 22226
rect 309678 22170 327250 22226
rect 327306 22170 327374 22226
rect 327430 22170 327498 22226
rect 327554 22170 327622 22226
rect 327678 22170 345250 22226
rect 345306 22170 345374 22226
rect 345430 22170 345498 22226
rect 345554 22170 345622 22226
rect 345678 22170 363250 22226
rect 363306 22170 363374 22226
rect 363430 22170 363498 22226
rect 363554 22170 363622 22226
rect 363678 22170 381250 22226
rect 381306 22170 381374 22226
rect 381430 22170 381498 22226
rect 381554 22170 381622 22226
rect 381678 22170 399250 22226
rect 399306 22170 399374 22226
rect 399430 22170 399498 22226
rect 399554 22170 399622 22226
rect 399678 22170 417250 22226
rect 417306 22170 417374 22226
rect 417430 22170 417498 22226
rect 417554 22170 417622 22226
rect 417678 22170 435250 22226
rect 435306 22170 435374 22226
rect 435430 22170 435498 22226
rect 435554 22170 435622 22226
rect 435678 22170 453250 22226
rect 453306 22170 453374 22226
rect 453430 22170 453498 22226
rect 453554 22170 453622 22226
rect 453678 22170 471250 22226
rect 471306 22170 471374 22226
rect 471430 22170 471498 22226
rect 471554 22170 471622 22226
rect 471678 22170 489250 22226
rect 489306 22170 489374 22226
rect 489430 22170 489498 22226
rect 489554 22170 489622 22226
rect 489678 22170 507250 22226
rect 507306 22170 507374 22226
rect 507430 22170 507498 22226
rect 507554 22170 507622 22226
rect 507678 22170 525250 22226
rect 525306 22170 525374 22226
rect 525430 22170 525498 22226
rect 525554 22170 525622 22226
rect 525678 22170 543250 22226
rect 543306 22170 543374 22226
rect 543430 22170 543498 22226
rect 543554 22170 543622 22226
rect 543678 22170 561250 22226
rect 561306 22170 561374 22226
rect 561430 22170 561498 22226
rect 561554 22170 561622 22226
rect 561678 22170 579250 22226
rect 579306 22170 579374 22226
rect 579430 22170 579498 22226
rect 579554 22170 579622 22226
rect 579678 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 3250 22102
rect 3306 22046 3374 22102
rect 3430 22046 3498 22102
rect 3554 22046 3622 22102
rect 3678 22046 21250 22102
rect 21306 22046 21374 22102
rect 21430 22046 21498 22102
rect 21554 22046 21622 22102
rect 21678 22046 39250 22102
rect 39306 22046 39374 22102
rect 39430 22046 39498 22102
rect 39554 22046 39622 22102
rect 39678 22046 57250 22102
rect 57306 22046 57374 22102
rect 57430 22046 57498 22102
rect 57554 22046 57622 22102
rect 57678 22046 75250 22102
rect 75306 22046 75374 22102
rect 75430 22046 75498 22102
rect 75554 22046 75622 22102
rect 75678 22046 93250 22102
rect 93306 22046 93374 22102
rect 93430 22046 93498 22102
rect 93554 22046 93622 22102
rect 93678 22046 111250 22102
rect 111306 22046 111374 22102
rect 111430 22046 111498 22102
rect 111554 22046 111622 22102
rect 111678 22046 129250 22102
rect 129306 22046 129374 22102
rect 129430 22046 129498 22102
rect 129554 22046 129622 22102
rect 129678 22046 147250 22102
rect 147306 22046 147374 22102
rect 147430 22046 147498 22102
rect 147554 22046 147622 22102
rect 147678 22046 165250 22102
rect 165306 22046 165374 22102
rect 165430 22046 165498 22102
rect 165554 22046 165622 22102
rect 165678 22046 183250 22102
rect 183306 22046 183374 22102
rect 183430 22046 183498 22102
rect 183554 22046 183622 22102
rect 183678 22046 201250 22102
rect 201306 22046 201374 22102
rect 201430 22046 201498 22102
rect 201554 22046 201622 22102
rect 201678 22046 219250 22102
rect 219306 22046 219374 22102
rect 219430 22046 219498 22102
rect 219554 22046 219622 22102
rect 219678 22046 237250 22102
rect 237306 22046 237374 22102
rect 237430 22046 237498 22102
rect 237554 22046 237622 22102
rect 237678 22046 255250 22102
rect 255306 22046 255374 22102
rect 255430 22046 255498 22102
rect 255554 22046 255622 22102
rect 255678 22046 273250 22102
rect 273306 22046 273374 22102
rect 273430 22046 273498 22102
rect 273554 22046 273622 22102
rect 273678 22046 291250 22102
rect 291306 22046 291374 22102
rect 291430 22046 291498 22102
rect 291554 22046 291622 22102
rect 291678 22046 309250 22102
rect 309306 22046 309374 22102
rect 309430 22046 309498 22102
rect 309554 22046 309622 22102
rect 309678 22046 327250 22102
rect 327306 22046 327374 22102
rect 327430 22046 327498 22102
rect 327554 22046 327622 22102
rect 327678 22046 345250 22102
rect 345306 22046 345374 22102
rect 345430 22046 345498 22102
rect 345554 22046 345622 22102
rect 345678 22046 363250 22102
rect 363306 22046 363374 22102
rect 363430 22046 363498 22102
rect 363554 22046 363622 22102
rect 363678 22046 381250 22102
rect 381306 22046 381374 22102
rect 381430 22046 381498 22102
rect 381554 22046 381622 22102
rect 381678 22046 399250 22102
rect 399306 22046 399374 22102
rect 399430 22046 399498 22102
rect 399554 22046 399622 22102
rect 399678 22046 417250 22102
rect 417306 22046 417374 22102
rect 417430 22046 417498 22102
rect 417554 22046 417622 22102
rect 417678 22046 435250 22102
rect 435306 22046 435374 22102
rect 435430 22046 435498 22102
rect 435554 22046 435622 22102
rect 435678 22046 453250 22102
rect 453306 22046 453374 22102
rect 453430 22046 453498 22102
rect 453554 22046 453622 22102
rect 453678 22046 471250 22102
rect 471306 22046 471374 22102
rect 471430 22046 471498 22102
rect 471554 22046 471622 22102
rect 471678 22046 489250 22102
rect 489306 22046 489374 22102
rect 489430 22046 489498 22102
rect 489554 22046 489622 22102
rect 489678 22046 507250 22102
rect 507306 22046 507374 22102
rect 507430 22046 507498 22102
rect 507554 22046 507622 22102
rect 507678 22046 525250 22102
rect 525306 22046 525374 22102
rect 525430 22046 525498 22102
rect 525554 22046 525622 22102
rect 525678 22046 543250 22102
rect 543306 22046 543374 22102
rect 543430 22046 543498 22102
rect 543554 22046 543622 22102
rect 543678 22046 561250 22102
rect 561306 22046 561374 22102
rect 561430 22046 561498 22102
rect 561554 22046 561622 22102
rect 561678 22046 579250 22102
rect 579306 22046 579374 22102
rect 579430 22046 579498 22102
rect 579554 22046 579622 22102
rect 579678 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 3250 21978
rect 3306 21922 3374 21978
rect 3430 21922 3498 21978
rect 3554 21922 3622 21978
rect 3678 21922 21250 21978
rect 21306 21922 21374 21978
rect 21430 21922 21498 21978
rect 21554 21922 21622 21978
rect 21678 21922 39250 21978
rect 39306 21922 39374 21978
rect 39430 21922 39498 21978
rect 39554 21922 39622 21978
rect 39678 21922 57250 21978
rect 57306 21922 57374 21978
rect 57430 21922 57498 21978
rect 57554 21922 57622 21978
rect 57678 21922 75250 21978
rect 75306 21922 75374 21978
rect 75430 21922 75498 21978
rect 75554 21922 75622 21978
rect 75678 21922 93250 21978
rect 93306 21922 93374 21978
rect 93430 21922 93498 21978
rect 93554 21922 93622 21978
rect 93678 21922 111250 21978
rect 111306 21922 111374 21978
rect 111430 21922 111498 21978
rect 111554 21922 111622 21978
rect 111678 21922 129250 21978
rect 129306 21922 129374 21978
rect 129430 21922 129498 21978
rect 129554 21922 129622 21978
rect 129678 21922 147250 21978
rect 147306 21922 147374 21978
rect 147430 21922 147498 21978
rect 147554 21922 147622 21978
rect 147678 21922 165250 21978
rect 165306 21922 165374 21978
rect 165430 21922 165498 21978
rect 165554 21922 165622 21978
rect 165678 21922 183250 21978
rect 183306 21922 183374 21978
rect 183430 21922 183498 21978
rect 183554 21922 183622 21978
rect 183678 21922 201250 21978
rect 201306 21922 201374 21978
rect 201430 21922 201498 21978
rect 201554 21922 201622 21978
rect 201678 21922 219250 21978
rect 219306 21922 219374 21978
rect 219430 21922 219498 21978
rect 219554 21922 219622 21978
rect 219678 21922 237250 21978
rect 237306 21922 237374 21978
rect 237430 21922 237498 21978
rect 237554 21922 237622 21978
rect 237678 21922 255250 21978
rect 255306 21922 255374 21978
rect 255430 21922 255498 21978
rect 255554 21922 255622 21978
rect 255678 21922 273250 21978
rect 273306 21922 273374 21978
rect 273430 21922 273498 21978
rect 273554 21922 273622 21978
rect 273678 21922 291250 21978
rect 291306 21922 291374 21978
rect 291430 21922 291498 21978
rect 291554 21922 291622 21978
rect 291678 21922 309250 21978
rect 309306 21922 309374 21978
rect 309430 21922 309498 21978
rect 309554 21922 309622 21978
rect 309678 21922 327250 21978
rect 327306 21922 327374 21978
rect 327430 21922 327498 21978
rect 327554 21922 327622 21978
rect 327678 21922 345250 21978
rect 345306 21922 345374 21978
rect 345430 21922 345498 21978
rect 345554 21922 345622 21978
rect 345678 21922 363250 21978
rect 363306 21922 363374 21978
rect 363430 21922 363498 21978
rect 363554 21922 363622 21978
rect 363678 21922 381250 21978
rect 381306 21922 381374 21978
rect 381430 21922 381498 21978
rect 381554 21922 381622 21978
rect 381678 21922 399250 21978
rect 399306 21922 399374 21978
rect 399430 21922 399498 21978
rect 399554 21922 399622 21978
rect 399678 21922 417250 21978
rect 417306 21922 417374 21978
rect 417430 21922 417498 21978
rect 417554 21922 417622 21978
rect 417678 21922 435250 21978
rect 435306 21922 435374 21978
rect 435430 21922 435498 21978
rect 435554 21922 435622 21978
rect 435678 21922 453250 21978
rect 453306 21922 453374 21978
rect 453430 21922 453498 21978
rect 453554 21922 453622 21978
rect 453678 21922 471250 21978
rect 471306 21922 471374 21978
rect 471430 21922 471498 21978
rect 471554 21922 471622 21978
rect 471678 21922 489250 21978
rect 489306 21922 489374 21978
rect 489430 21922 489498 21978
rect 489554 21922 489622 21978
rect 489678 21922 507250 21978
rect 507306 21922 507374 21978
rect 507430 21922 507498 21978
rect 507554 21922 507622 21978
rect 507678 21922 525250 21978
rect 525306 21922 525374 21978
rect 525430 21922 525498 21978
rect 525554 21922 525622 21978
rect 525678 21922 543250 21978
rect 543306 21922 543374 21978
rect 543430 21922 543498 21978
rect 543554 21922 543622 21978
rect 543678 21922 561250 21978
rect 561306 21922 561374 21978
rect 561430 21922 561498 21978
rect 561554 21922 561622 21978
rect 561678 21922 579250 21978
rect 579306 21922 579374 21978
rect 579430 21922 579498 21978
rect 579554 21922 579622 21978
rect 579678 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 6970 10350
rect 7026 10294 7094 10350
rect 7150 10294 7218 10350
rect 7274 10294 7342 10350
rect 7398 10294 24970 10350
rect 25026 10294 25094 10350
rect 25150 10294 25218 10350
rect 25274 10294 25342 10350
rect 25398 10294 42970 10350
rect 43026 10294 43094 10350
rect 43150 10294 43218 10350
rect 43274 10294 43342 10350
rect 43398 10294 60970 10350
rect 61026 10294 61094 10350
rect 61150 10294 61218 10350
rect 61274 10294 61342 10350
rect 61398 10294 78970 10350
rect 79026 10294 79094 10350
rect 79150 10294 79218 10350
rect 79274 10294 79342 10350
rect 79398 10294 96970 10350
rect 97026 10294 97094 10350
rect 97150 10294 97218 10350
rect 97274 10294 97342 10350
rect 97398 10294 114970 10350
rect 115026 10294 115094 10350
rect 115150 10294 115218 10350
rect 115274 10294 115342 10350
rect 115398 10294 132970 10350
rect 133026 10294 133094 10350
rect 133150 10294 133218 10350
rect 133274 10294 133342 10350
rect 133398 10294 150970 10350
rect 151026 10294 151094 10350
rect 151150 10294 151218 10350
rect 151274 10294 151342 10350
rect 151398 10294 168970 10350
rect 169026 10294 169094 10350
rect 169150 10294 169218 10350
rect 169274 10294 169342 10350
rect 169398 10294 186970 10350
rect 187026 10294 187094 10350
rect 187150 10294 187218 10350
rect 187274 10294 187342 10350
rect 187398 10294 204970 10350
rect 205026 10294 205094 10350
rect 205150 10294 205218 10350
rect 205274 10294 205342 10350
rect 205398 10294 222970 10350
rect 223026 10294 223094 10350
rect 223150 10294 223218 10350
rect 223274 10294 223342 10350
rect 223398 10294 240970 10350
rect 241026 10294 241094 10350
rect 241150 10294 241218 10350
rect 241274 10294 241342 10350
rect 241398 10294 258970 10350
rect 259026 10294 259094 10350
rect 259150 10294 259218 10350
rect 259274 10294 259342 10350
rect 259398 10294 276970 10350
rect 277026 10294 277094 10350
rect 277150 10294 277218 10350
rect 277274 10294 277342 10350
rect 277398 10294 294970 10350
rect 295026 10294 295094 10350
rect 295150 10294 295218 10350
rect 295274 10294 295342 10350
rect 295398 10294 312970 10350
rect 313026 10294 313094 10350
rect 313150 10294 313218 10350
rect 313274 10294 313342 10350
rect 313398 10294 330970 10350
rect 331026 10294 331094 10350
rect 331150 10294 331218 10350
rect 331274 10294 331342 10350
rect 331398 10294 348970 10350
rect 349026 10294 349094 10350
rect 349150 10294 349218 10350
rect 349274 10294 349342 10350
rect 349398 10294 366970 10350
rect 367026 10294 367094 10350
rect 367150 10294 367218 10350
rect 367274 10294 367342 10350
rect 367398 10294 384970 10350
rect 385026 10294 385094 10350
rect 385150 10294 385218 10350
rect 385274 10294 385342 10350
rect 385398 10294 402970 10350
rect 403026 10294 403094 10350
rect 403150 10294 403218 10350
rect 403274 10294 403342 10350
rect 403398 10294 420970 10350
rect 421026 10294 421094 10350
rect 421150 10294 421218 10350
rect 421274 10294 421342 10350
rect 421398 10294 438970 10350
rect 439026 10294 439094 10350
rect 439150 10294 439218 10350
rect 439274 10294 439342 10350
rect 439398 10294 456970 10350
rect 457026 10294 457094 10350
rect 457150 10294 457218 10350
rect 457274 10294 457342 10350
rect 457398 10294 474970 10350
rect 475026 10294 475094 10350
rect 475150 10294 475218 10350
rect 475274 10294 475342 10350
rect 475398 10294 492970 10350
rect 493026 10294 493094 10350
rect 493150 10294 493218 10350
rect 493274 10294 493342 10350
rect 493398 10294 510970 10350
rect 511026 10294 511094 10350
rect 511150 10294 511218 10350
rect 511274 10294 511342 10350
rect 511398 10294 528970 10350
rect 529026 10294 529094 10350
rect 529150 10294 529218 10350
rect 529274 10294 529342 10350
rect 529398 10294 546970 10350
rect 547026 10294 547094 10350
rect 547150 10294 547218 10350
rect 547274 10294 547342 10350
rect 547398 10294 564970 10350
rect 565026 10294 565094 10350
rect 565150 10294 565218 10350
rect 565274 10294 565342 10350
rect 565398 10294 582970 10350
rect 583026 10294 583094 10350
rect 583150 10294 583218 10350
rect 583274 10294 583342 10350
rect 583398 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 6970 10226
rect 7026 10170 7094 10226
rect 7150 10170 7218 10226
rect 7274 10170 7342 10226
rect 7398 10170 24970 10226
rect 25026 10170 25094 10226
rect 25150 10170 25218 10226
rect 25274 10170 25342 10226
rect 25398 10170 42970 10226
rect 43026 10170 43094 10226
rect 43150 10170 43218 10226
rect 43274 10170 43342 10226
rect 43398 10170 60970 10226
rect 61026 10170 61094 10226
rect 61150 10170 61218 10226
rect 61274 10170 61342 10226
rect 61398 10170 78970 10226
rect 79026 10170 79094 10226
rect 79150 10170 79218 10226
rect 79274 10170 79342 10226
rect 79398 10170 96970 10226
rect 97026 10170 97094 10226
rect 97150 10170 97218 10226
rect 97274 10170 97342 10226
rect 97398 10170 114970 10226
rect 115026 10170 115094 10226
rect 115150 10170 115218 10226
rect 115274 10170 115342 10226
rect 115398 10170 132970 10226
rect 133026 10170 133094 10226
rect 133150 10170 133218 10226
rect 133274 10170 133342 10226
rect 133398 10170 150970 10226
rect 151026 10170 151094 10226
rect 151150 10170 151218 10226
rect 151274 10170 151342 10226
rect 151398 10170 168970 10226
rect 169026 10170 169094 10226
rect 169150 10170 169218 10226
rect 169274 10170 169342 10226
rect 169398 10170 186970 10226
rect 187026 10170 187094 10226
rect 187150 10170 187218 10226
rect 187274 10170 187342 10226
rect 187398 10170 204970 10226
rect 205026 10170 205094 10226
rect 205150 10170 205218 10226
rect 205274 10170 205342 10226
rect 205398 10170 222970 10226
rect 223026 10170 223094 10226
rect 223150 10170 223218 10226
rect 223274 10170 223342 10226
rect 223398 10170 240970 10226
rect 241026 10170 241094 10226
rect 241150 10170 241218 10226
rect 241274 10170 241342 10226
rect 241398 10170 258970 10226
rect 259026 10170 259094 10226
rect 259150 10170 259218 10226
rect 259274 10170 259342 10226
rect 259398 10170 276970 10226
rect 277026 10170 277094 10226
rect 277150 10170 277218 10226
rect 277274 10170 277342 10226
rect 277398 10170 294970 10226
rect 295026 10170 295094 10226
rect 295150 10170 295218 10226
rect 295274 10170 295342 10226
rect 295398 10170 312970 10226
rect 313026 10170 313094 10226
rect 313150 10170 313218 10226
rect 313274 10170 313342 10226
rect 313398 10170 330970 10226
rect 331026 10170 331094 10226
rect 331150 10170 331218 10226
rect 331274 10170 331342 10226
rect 331398 10170 348970 10226
rect 349026 10170 349094 10226
rect 349150 10170 349218 10226
rect 349274 10170 349342 10226
rect 349398 10170 366970 10226
rect 367026 10170 367094 10226
rect 367150 10170 367218 10226
rect 367274 10170 367342 10226
rect 367398 10170 384970 10226
rect 385026 10170 385094 10226
rect 385150 10170 385218 10226
rect 385274 10170 385342 10226
rect 385398 10170 402970 10226
rect 403026 10170 403094 10226
rect 403150 10170 403218 10226
rect 403274 10170 403342 10226
rect 403398 10170 420970 10226
rect 421026 10170 421094 10226
rect 421150 10170 421218 10226
rect 421274 10170 421342 10226
rect 421398 10170 438970 10226
rect 439026 10170 439094 10226
rect 439150 10170 439218 10226
rect 439274 10170 439342 10226
rect 439398 10170 456970 10226
rect 457026 10170 457094 10226
rect 457150 10170 457218 10226
rect 457274 10170 457342 10226
rect 457398 10170 474970 10226
rect 475026 10170 475094 10226
rect 475150 10170 475218 10226
rect 475274 10170 475342 10226
rect 475398 10170 492970 10226
rect 493026 10170 493094 10226
rect 493150 10170 493218 10226
rect 493274 10170 493342 10226
rect 493398 10170 510970 10226
rect 511026 10170 511094 10226
rect 511150 10170 511218 10226
rect 511274 10170 511342 10226
rect 511398 10170 528970 10226
rect 529026 10170 529094 10226
rect 529150 10170 529218 10226
rect 529274 10170 529342 10226
rect 529398 10170 546970 10226
rect 547026 10170 547094 10226
rect 547150 10170 547218 10226
rect 547274 10170 547342 10226
rect 547398 10170 564970 10226
rect 565026 10170 565094 10226
rect 565150 10170 565218 10226
rect 565274 10170 565342 10226
rect 565398 10170 582970 10226
rect 583026 10170 583094 10226
rect 583150 10170 583218 10226
rect 583274 10170 583342 10226
rect 583398 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 6970 10102
rect 7026 10046 7094 10102
rect 7150 10046 7218 10102
rect 7274 10046 7342 10102
rect 7398 10046 24970 10102
rect 25026 10046 25094 10102
rect 25150 10046 25218 10102
rect 25274 10046 25342 10102
rect 25398 10046 42970 10102
rect 43026 10046 43094 10102
rect 43150 10046 43218 10102
rect 43274 10046 43342 10102
rect 43398 10046 60970 10102
rect 61026 10046 61094 10102
rect 61150 10046 61218 10102
rect 61274 10046 61342 10102
rect 61398 10046 78970 10102
rect 79026 10046 79094 10102
rect 79150 10046 79218 10102
rect 79274 10046 79342 10102
rect 79398 10046 96970 10102
rect 97026 10046 97094 10102
rect 97150 10046 97218 10102
rect 97274 10046 97342 10102
rect 97398 10046 114970 10102
rect 115026 10046 115094 10102
rect 115150 10046 115218 10102
rect 115274 10046 115342 10102
rect 115398 10046 132970 10102
rect 133026 10046 133094 10102
rect 133150 10046 133218 10102
rect 133274 10046 133342 10102
rect 133398 10046 150970 10102
rect 151026 10046 151094 10102
rect 151150 10046 151218 10102
rect 151274 10046 151342 10102
rect 151398 10046 168970 10102
rect 169026 10046 169094 10102
rect 169150 10046 169218 10102
rect 169274 10046 169342 10102
rect 169398 10046 186970 10102
rect 187026 10046 187094 10102
rect 187150 10046 187218 10102
rect 187274 10046 187342 10102
rect 187398 10046 204970 10102
rect 205026 10046 205094 10102
rect 205150 10046 205218 10102
rect 205274 10046 205342 10102
rect 205398 10046 222970 10102
rect 223026 10046 223094 10102
rect 223150 10046 223218 10102
rect 223274 10046 223342 10102
rect 223398 10046 240970 10102
rect 241026 10046 241094 10102
rect 241150 10046 241218 10102
rect 241274 10046 241342 10102
rect 241398 10046 258970 10102
rect 259026 10046 259094 10102
rect 259150 10046 259218 10102
rect 259274 10046 259342 10102
rect 259398 10046 276970 10102
rect 277026 10046 277094 10102
rect 277150 10046 277218 10102
rect 277274 10046 277342 10102
rect 277398 10046 294970 10102
rect 295026 10046 295094 10102
rect 295150 10046 295218 10102
rect 295274 10046 295342 10102
rect 295398 10046 312970 10102
rect 313026 10046 313094 10102
rect 313150 10046 313218 10102
rect 313274 10046 313342 10102
rect 313398 10046 330970 10102
rect 331026 10046 331094 10102
rect 331150 10046 331218 10102
rect 331274 10046 331342 10102
rect 331398 10046 348970 10102
rect 349026 10046 349094 10102
rect 349150 10046 349218 10102
rect 349274 10046 349342 10102
rect 349398 10046 366970 10102
rect 367026 10046 367094 10102
rect 367150 10046 367218 10102
rect 367274 10046 367342 10102
rect 367398 10046 384970 10102
rect 385026 10046 385094 10102
rect 385150 10046 385218 10102
rect 385274 10046 385342 10102
rect 385398 10046 402970 10102
rect 403026 10046 403094 10102
rect 403150 10046 403218 10102
rect 403274 10046 403342 10102
rect 403398 10046 420970 10102
rect 421026 10046 421094 10102
rect 421150 10046 421218 10102
rect 421274 10046 421342 10102
rect 421398 10046 438970 10102
rect 439026 10046 439094 10102
rect 439150 10046 439218 10102
rect 439274 10046 439342 10102
rect 439398 10046 456970 10102
rect 457026 10046 457094 10102
rect 457150 10046 457218 10102
rect 457274 10046 457342 10102
rect 457398 10046 474970 10102
rect 475026 10046 475094 10102
rect 475150 10046 475218 10102
rect 475274 10046 475342 10102
rect 475398 10046 492970 10102
rect 493026 10046 493094 10102
rect 493150 10046 493218 10102
rect 493274 10046 493342 10102
rect 493398 10046 510970 10102
rect 511026 10046 511094 10102
rect 511150 10046 511218 10102
rect 511274 10046 511342 10102
rect 511398 10046 528970 10102
rect 529026 10046 529094 10102
rect 529150 10046 529218 10102
rect 529274 10046 529342 10102
rect 529398 10046 546970 10102
rect 547026 10046 547094 10102
rect 547150 10046 547218 10102
rect 547274 10046 547342 10102
rect 547398 10046 564970 10102
rect 565026 10046 565094 10102
rect 565150 10046 565218 10102
rect 565274 10046 565342 10102
rect 565398 10046 582970 10102
rect 583026 10046 583094 10102
rect 583150 10046 583218 10102
rect 583274 10046 583342 10102
rect 583398 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 6970 9978
rect 7026 9922 7094 9978
rect 7150 9922 7218 9978
rect 7274 9922 7342 9978
rect 7398 9922 24970 9978
rect 25026 9922 25094 9978
rect 25150 9922 25218 9978
rect 25274 9922 25342 9978
rect 25398 9922 42970 9978
rect 43026 9922 43094 9978
rect 43150 9922 43218 9978
rect 43274 9922 43342 9978
rect 43398 9922 60970 9978
rect 61026 9922 61094 9978
rect 61150 9922 61218 9978
rect 61274 9922 61342 9978
rect 61398 9922 78970 9978
rect 79026 9922 79094 9978
rect 79150 9922 79218 9978
rect 79274 9922 79342 9978
rect 79398 9922 96970 9978
rect 97026 9922 97094 9978
rect 97150 9922 97218 9978
rect 97274 9922 97342 9978
rect 97398 9922 114970 9978
rect 115026 9922 115094 9978
rect 115150 9922 115218 9978
rect 115274 9922 115342 9978
rect 115398 9922 132970 9978
rect 133026 9922 133094 9978
rect 133150 9922 133218 9978
rect 133274 9922 133342 9978
rect 133398 9922 150970 9978
rect 151026 9922 151094 9978
rect 151150 9922 151218 9978
rect 151274 9922 151342 9978
rect 151398 9922 168970 9978
rect 169026 9922 169094 9978
rect 169150 9922 169218 9978
rect 169274 9922 169342 9978
rect 169398 9922 186970 9978
rect 187026 9922 187094 9978
rect 187150 9922 187218 9978
rect 187274 9922 187342 9978
rect 187398 9922 204970 9978
rect 205026 9922 205094 9978
rect 205150 9922 205218 9978
rect 205274 9922 205342 9978
rect 205398 9922 222970 9978
rect 223026 9922 223094 9978
rect 223150 9922 223218 9978
rect 223274 9922 223342 9978
rect 223398 9922 240970 9978
rect 241026 9922 241094 9978
rect 241150 9922 241218 9978
rect 241274 9922 241342 9978
rect 241398 9922 258970 9978
rect 259026 9922 259094 9978
rect 259150 9922 259218 9978
rect 259274 9922 259342 9978
rect 259398 9922 276970 9978
rect 277026 9922 277094 9978
rect 277150 9922 277218 9978
rect 277274 9922 277342 9978
rect 277398 9922 294970 9978
rect 295026 9922 295094 9978
rect 295150 9922 295218 9978
rect 295274 9922 295342 9978
rect 295398 9922 312970 9978
rect 313026 9922 313094 9978
rect 313150 9922 313218 9978
rect 313274 9922 313342 9978
rect 313398 9922 330970 9978
rect 331026 9922 331094 9978
rect 331150 9922 331218 9978
rect 331274 9922 331342 9978
rect 331398 9922 348970 9978
rect 349026 9922 349094 9978
rect 349150 9922 349218 9978
rect 349274 9922 349342 9978
rect 349398 9922 366970 9978
rect 367026 9922 367094 9978
rect 367150 9922 367218 9978
rect 367274 9922 367342 9978
rect 367398 9922 384970 9978
rect 385026 9922 385094 9978
rect 385150 9922 385218 9978
rect 385274 9922 385342 9978
rect 385398 9922 402970 9978
rect 403026 9922 403094 9978
rect 403150 9922 403218 9978
rect 403274 9922 403342 9978
rect 403398 9922 420970 9978
rect 421026 9922 421094 9978
rect 421150 9922 421218 9978
rect 421274 9922 421342 9978
rect 421398 9922 438970 9978
rect 439026 9922 439094 9978
rect 439150 9922 439218 9978
rect 439274 9922 439342 9978
rect 439398 9922 456970 9978
rect 457026 9922 457094 9978
rect 457150 9922 457218 9978
rect 457274 9922 457342 9978
rect 457398 9922 474970 9978
rect 475026 9922 475094 9978
rect 475150 9922 475218 9978
rect 475274 9922 475342 9978
rect 475398 9922 492970 9978
rect 493026 9922 493094 9978
rect 493150 9922 493218 9978
rect 493274 9922 493342 9978
rect 493398 9922 510970 9978
rect 511026 9922 511094 9978
rect 511150 9922 511218 9978
rect 511274 9922 511342 9978
rect 511398 9922 528970 9978
rect 529026 9922 529094 9978
rect 529150 9922 529218 9978
rect 529274 9922 529342 9978
rect 529398 9922 546970 9978
rect 547026 9922 547094 9978
rect 547150 9922 547218 9978
rect 547274 9922 547342 9978
rect 547398 9922 564970 9978
rect 565026 9922 565094 9978
rect 565150 9922 565218 9978
rect 565274 9922 565342 9978
rect 565398 9922 582970 9978
rect 583026 9922 583094 9978
rect 583150 9922 583218 9978
rect 583274 9922 583342 9978
rect 583398 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 3250 4350
rect 3306 4294 3374 4350
rect 3430 4294 3498 4350
rect 3554 4294 3622 4350
rect 3678 4294 21250 4350
rect 21306 4294 21374 4350
rect 21430 4294 21498 4350
rect 21554 4294 21622 4350
rect 21678 4294 39250 4350
rect 39306 4294 39374 4350
rect 39430 4294 39498 4350
rect 39554 4294 39622 4350
rect 39678 4294 57250 4350
rect 57306 4294 57374 4350
rect 57430 4294 57498 4350
rect 57554 4294 57622 4350
rect 57678 4294 75250 4350
rect 75306 4294 75374 4350
rect 75430 4294 75498 4350
rect 75554 4294 75622 4350
rect 75678 4294 93250 4350
rect 93306 4294 93374 4350
rect 93430 4294 93498 4350
rect 93554 4294 93622 4350
rect 93678 4294 111250 4350
rect 111306 4294 111374 4350
rect 111430 4294 111498 4350
rect 111554 4294 111622 4350
rect 111678 4294 129250 4350
rect 129306 4294 129374 4350
rect 129430 4294 129498 4350
rect 129554 4294 129622 4350
rect 129678 4294 147250 4350
rect 147306 4294 147374 4350
rect 147430 4294 147498 4350
rect 147554 4294 147622 4350
rect 147678 4294 165250 4350
rect 165306 4294 165374 4350
rect 165430 4294 165498 4350
rect 165554 4294 165622 4350
rect 165678 4294 183250 4350
rect 183306 4294 183374 4350
rect 183430 4294 183498 4350
rect 183554 4294 183622 4350
rect 183678 4294 201250 4350
rect 201306 4294 201374 4350
rect 201430 4294 201498 4350
rect 201554 4294 201622 4350
rect 201678 4294 219250 4350
rect 219306 4294 219374 4350
rect 219430 4294 219498 4350
rect 219554 4294 219622 4350
rect 219678 4294 237250 4350
rect 237306 4294 237374 4350
rect 237430 4294 237498 4350
rect 237554 4294 237622 4350
rect 237678 4294 255250 4350
rect 255306 4294 255374 4350
rect 255430 4294 255498 4350
rect 255554 4294 255622 4350
rect 255678 4294 273250 4350
rect 273306 4294 273374 4350
rect 273430 4294 273498 4350
rect 273554 4294 273622 4350
rect 273678 4294 291250 4350
rect 291306 4294 291374 4350
rect 291430 4294 291498 4350
rect 291554 4294 291622 4350
rect 291678 4294 309250 4350
rect 309306 4294 309374 4350
rect 309430 4294 309498 4350
rect 309554 4294 309622 4350
rect 309678 4294 327250 4350
rect 327306 4294 327374 4350
rect 327430 4294 327498 4350
rect 327554 4294 327622 4350
rect 327678 4294 345250 4350
rect 345306 4294 345374 4350
rect 345430 4294 345498 4350
rect 345554 4294 345622 4350
rect 345678 4294 363250 4350
rect 363306 4294 363374 4350
rect 363430 4294 363498 4350
rect 363554 4294 363622 4350
rect 363678 4294 381250 4350
rect 381306 4294 381374 4350
rect 381430 4294 381498 4350
rect 381554 4294 381622 4350
rect 381678 4294 399250 4350
rect 399306 4294 399374 4350
rect 399430 4294 399498 4350
rect 399554 4294 399622 4350
rect 399678 4294 417250 4350
rect 417306 4294 417374 4350
rect 417430 4294 417498 4350
rect 417554 4294 417622 4350
rect 417678 4294 435250 4350
rect 435306 4294 435374 4350
rect 435430 4294 435498 4350
rect 435554 4294 435622 4350
rect 435678 4294 453250 4350
rect 453306 4294 453374 4350
rect 453430 4294 453498 4350
rect 453554 4294 453622 4350
rect 453678 4294 471250 4350
rect 471306 4294 471374 4350
rect 471430 4294 471498 4350
rect 471554 4294 471622 4350
rect 471678 4294 489250 4350
rect 489306 4294 489374 4350
rect 489430 4294 489498 4350
rect 489554 4294 489622 4350
rect 489678 4294 507250 4350
rect 507306 4294 507374 4350
rect 507430 4294 507498 4350
rect 507554 4294 507622 4350
rect 507678 4294 525250 4350
rect 525306 4294 525374 4350
rect 525430 4294 525498 4350
rect 525554 4294 525622 4350
rect 525678 4294 543250 4350
rect 543306 4294 543374 4350
rect 543430 4294 543498 4350
rect 543554 4294 543622 4350
rect 543678 4294 561250 4350
rect 561306 4294 561374 4350
rect 561430 4294 561498 4350
rect 561554 4294 561622 4350
rect 561678 4294 579250 4350
rect 579306 4294 579374 4350
rect 579430 4294 579498 4350
rect 579554 4294 579622 4350
rect 579678 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 3250 4226
rect 3306 4170 3374 4226
rect 3430 4170 3498 4226
rect 3554 4170 3622 4226
rect 3678 4170 21250 4226
rect 21306 4170 21374 4226
rect 21430 4170 21498 4226
rect 21554 4170 21622 4226
rect 21678 4170 39250 4226
rect 39306 4170 39374 4226
rect 39430 4170 39498 4226
rect 39554 4170 39622 4226
rect 39678 4170 57250 4226
rect 57306 4170 57374 4226
rect 57430 4170 57498 4226
rect 57554 4170 57622 4226
rect 57678 4170 75250 4226
rect 75306 4170 75374 4226
rect 75430 4170 75498 4226
rect 75554 4170 75622 4226
rect 75678 4170 93250 4226
rect 93306 4170 93374 4226
rect 93430 4170 93498 4226
rect 93554 4170 93622 4226
rect 93678 4170 111250 4226
rect 111306 4170 111374 4226
rect 111430 4170 111498 4226
rect 111554 4170 111622 4226
rect 111678 4170 129250 4226
rect 129306 4170 129374 4226
rect 129430 4170 129498 4226
rect 129554 4170 129622 4226
rect 129678 4170 147250 4226
rect 147306 4170 147374 4226
rect 147430 4170 147498 4226
rect 147554 4170 147622 4226
rect 147678 4170 165250 4226
rect 165306 4170 165374 4226
rect 165430 4170 165498 4226
rect 165554 4170 165622 4226
rect 165678 4170 183250 4226
rect 183306 4170 183374 4226
rect 183430 4170 183498 4226
rect 183554 4170 183622 4226
rect 183678 4170 201250 4226
rect 201306 4170 201374 4226
rect 201430 4170 201498 4226
rect 201554 4170 201622 4226
rect 201678 4170 219250 4226
rect 219306 4170 219374 4226
rect 219430 4170 219498 4226
rect 219554 4170 219622 4226
rect 219678 4170 237250 4226
rect 237306 4170 237374 4226
rect 237430 4170 237498 4226
rect 237554 4170 237622 4226
rect 237678 4170 255250 4226
rect 255306 4170 255374 4226
rect 255430 4170 255498 4226
rect 255554 4170 255622 4226
rect 255678 4170 273250 4226
rect 273306 4170 273374 4226
rect 273430 4170 273498 4226
rect 273554 4170 273622 4226
rect 273678 4170 291250 4226
rect 291306 4170 291374 4226
rect 291430 4170 291498 4226
rect 291554 4170 291622 4226
rect 291678 4170 309250 4226
rect 309306 4170 309374 4226
rect 309430 4170 309498 4226
rect 309554 4170 309622 4226
rect 309678 4170 327250 4226
rect 327306 4170 327374 4226
rect 327430 4170 327498 4226
rect 327554 4170 327622 4226
rect 327678 4170 345250 4226
rect 345306 4170 345374 4226
rect 345430 4170 345498 4226
rect 345554 4170 345622 4226
rect 345678 4170 363250 4226
rect 363306 4170 363374 4226
rect 363430 4170 363498 4226
rect 363554 4170 363622 4226
rect 363678 4170 381250 4226
rect 381306 4170 381374 4226
rect 381430 4170 381498 4226
rect 381554 4170 381622 4226
rect 381678 4170 399250 4226
rect 399306 4170 399374 4226
rect 399430 4170 399498 4226
rect 399554 4170 399622 4226
rect 399678 4170 417250 4226
rect 417306 4170 417374 4226
rect 417430 4170 417498 4226
rect 417554 4170 417622 4226
rect 417678 4170 435250 4226
rect 435306 4170 435374 4226
rect 435430 4170 435498 4226
rect 435554 4170 435622 4226
rect 435678 4170 453250 4226
rect 453306 4170 453374 4226
rect 453430 4170 453498 4226
rect 453554 4170 453622 4226
rect 453678 4170 471250 4226
rect 471306 4170 471374 4226
rect 471430 4170 471498 4226
rect 471554 4170 471622 4226
rect 471678 4170 489250 4226
rect 489306 4170 489374 4226
rect 489430 4170 489498 4226
rect 489554 4170 489622 4226
rect 489678 4170 507250 4226
rect 507306 4170 507374 4226
rect 507430 4170 507498 4226
rect 507554 4170 507622 4226
rect 507678 4170 525250 4226
rect 525306 4170 525374 4226
rect 525430 4170 525498 4226
rect 525554 4170 525622 4226
rect 525678 4170 543250 4226
rect 543306 4170 543374 4226
rect 543430 4170 543498 4226
rect 543554 4170 543622 4226
rect 543678 4170 561250 4226
rect 561306 4170 561374 4226
rect 561430 4170 561498 4226
rect 561554 4170 561622 4226
rect 561678 4170 579250 4226
rect 579306 4170 579374 4226
rect 579430 4170 579498 4226
rect 579554 4170 579622 4226
rect 579678 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 3250 4102
rect 3306 4046 3374 4102
rect 3430 4046 3498 4102
rect 3554 4046 3622 4102
rect 3678 4046 21250 4102
rect 21306 4046 21374 4102
rect 21430 4046 21498 4102
rect 21554 4046 21622 4102
rect 21678 4046 39250 4102
rect 39306 4046 39374 4102
rect 39430 4046 39498 4102
rect 39554 4046 39622 4102
rect 39678 4046 57250 4102
rect 57306 4046 57374 4102
rect 57430 4046 57498 4102
rect 57554 4046 57622 4102
rect 57678 4046 75250 4102
rect 75306 4046 75374 4102
rect 75430 4046 75498 4102
rect 75554 4046 75622 4102
rect 75678 4046 93250 4102
rect 93306 4046 93374 4102
rect 93430 4046 93498 4102
rect 93554 4046 93622 4102
rect 93678 4046 111250 4102
rect 111306 4046 111374 4102
rect 111430 4046 111498 4102
rect 111554 4046 111622 4102
rect 111678 4046 129250 4102
rect 129306 4046 129374 4102
rect 129430 4046 129498 4102
rect 129554 4046 129622 4102
rect 129678 4046 147250 4102
rect 147306 4046 147374 4102
rect 147430 4046 147498 4102
rect 147554 4046 147622 4102
rect 147678 4046 165250 4102
rect 165306 4046 165374 4102
rect 165430 4046 165498 4102
rect 165554 4046 165622 4102
rect 165678 4046 183250 4102
rect 183306 4046 183374 4102
rect 183430 4046 183498 4102
rect 183554 4046 183622 4102
rect 183678 4046 201250 4102
rect 201306 4046 201374 4102
rect 201430 4046 201498 4102
rect 201554 4046 201622 4102
rect 201678 4046 219250 4102
rect 219306 4046 219374 4102
rect 219430 4046 219498 4102
rect 219554 4046 219622 4102
rect 219678 4046 237250 4102
rect 237306 4046 237374 4102
rect 237430 4046 237498 4102
rect 237554 4046 237622 4102
rect 237678 4046 255250 4102
rect 255306 4046 255374 4102
rect 255430 4046 255498 4102
rect 255554 4046 255622 4102
rect 255678 4046 273250 4102
rect 273306 4046 273374 4102
rect 273430 4046 273498 4102
rect 273554 4046 273622 4102
rect 273678 4046 291250 4102
rect 291306 4046 291374 4102
rect 291430 4046 291498 4102
rect 291554 4046 291622 4102
rect 291678 4046 309250 4102
rect 309306 4046 309374 4102
rect 309430 4046 309498 4102
rect 309554 4046 309622 4102
rect 309678 4046 327250 4102
rect 327306 4046 327374 4102
rect 327430 4046 327498 4102
rect 327554 4046 327622 4102
rect 327678 4046 345250 4102
rect 345306 4046 345374 4102
rect 345430 4046 345498 4102
rect 345554 4046 345622 4102
rect 345678 4046 363250 4102
rect 363306 4046 363374 4102
rect 363430 4046 363498 4102
rect 363554 4046 363622 4102
rect 363678 4046 381250 4102
rect 381306 4046 381374 4102
rect 381430 4046 381498 4102
rect 381554 4046 381622 4102
rect 381678 4046 399250 4102
rect 399306 4046 399374 4102
rect 399430 4046 399498 4102
rect 399554 4046 399622 4102
rect 399678 4046 417250 4102
rect 417306 4046 417374 4102
rect 417430 4046 417498 4102
rect 417554 4046 417622 4102
rect 417678 4046 435250 4102
rect 435306 4046 435374 4102
rect 435430 4046 435498 4102
rect 435554 4046 435622 4102
rect 435678 4046 453250 4102
rect 453306 4046 453374 4102
rect 453430 4046 453498 4102
rect 453554 4046 453622 4102
rect 453678 4046 471250 4102
rect 471306 4046 471374 4102
rect 471430 4046 471498 4102
rect 471554 4046 471622 4102
rect 471678 4046 489250 4102
rect 489306 4046 489374 4102
rect 489430 4046 489498 4102
rect 489554 4046 489622 4102
rect 489678 4046 507250 4102
rect 507306 4046 507374 4102
rect 507430 4046 507498 4102
rect 507554 4046 507622 4102
rect 507678 4046 525250 4102
rect 525306 4046 525374 4102
rect 525430 4046 525498 4102
rect 525554 4046 525622 4102
rect 525678 4046 543250 4102
rect 543306 4046 543374 4102
rect 543430 4046 543498 4102
rect 543554 4046 543622 4102
rect 543678 4046 561250 4102
rect 561306 4046 561374 4102
rect 561430 4046 561498 4102
rect 561554 4046 561622 4102
rect 561678 4046 579250 4102
rect 579306 4046 579374 4102
rect 579430 4046 579498 4102
rect 579554 4046 579622 4102
rect 579678 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 3250 3978
rect 3306 3922 3374 3978
rect 3430 3922 3498 3978
rect 3554 3922 3622 3978
rect 3678 3922 21250 3978
rect 21306 3922 21374 3978
rect 21430 3922 21498 3978
rect 21554 3922 21622 3978
rect 21678 3922 39250 3978
rect 39306 3922 39374 3978
rect 39430 3922 39498 3978
rect 39554 3922 39622 3978
rect 39678 3922 57250 3978
rect 57306 3922 57374 3978
rect 57430 3922 57498 3978
rect 57554 3922 57622 3978
rect 57678 3922 75250 3978
rect 75306 3922 75374 3978
rect 75430 3922 75498 3978
rect 75554 3922 75622 3978
rect 75678 3922 93250 3978
rect 93306 3922 93374 3978
rect 93430 3922 93498 3978
rect 93554 3922 93622 3978
rect 93678 3922 111250 3978
rect 111306 3922 111374 3978
rect 111430 3922 111498 3978
rect 111554 3922 111622 3978
rect 111678 3922 129250 3978
rect 129306 3922 129374 3978
rect 129430 3922 129498 3978
rect 129554 3922 129622 3978
rect 129678 3922 147250 3978
rect 147306 3922 147374 3978
rect 147430 3922 147498 3978
rect 147554 3922 147622 3978
rect 147678 3922 165250 3978
rect 165306 3922 165374 3978
rect 165430 3922 165498 3978
rect 165554 3922 165622 3978
rect 165678 3922 183250 3978
rect 183306 3922 183374 3978
rect 183430 3922 183498 3978
rect 183554 3922 183622 3978
rect 183678 3922 201250 3978
rect 201306 3922 201374 3978
rect 201430 3922 201498 3978
rect 201554 3922 201622 3978
rect 201678 3922 219250 3978
rect 219306 3922 219374 3978
rect 219430 3922 219498 3978
rect 219554 3922 219622 3978
rect 219678 3922 237250 3978
rect 237306 3922 237374 3978
rect 237430 3922 237498 3978
rect 237554 3922 237622 3978
rect 237678 3922 255250 3978
rect 255306 3922 255374 3978
rect 255430 3922 255498 3978
rect 255554 3922 255622 3978
rect 255678 3922 273250 3978
rect 273306 3922 273374 3978
rect 273430 3922 273498 3978
rect 273554 3922 273622 3978
rect 273678 3922 291250 3978
rect 291306 3922 291374 3978
rect 291430 3922 291498 3978
rect 291554 3922 291622 3978
rect 291678 3922 309250 3978
rect 309306 3922 309374 3978
rect 309430 3922 309498 3978
rect 309554 3922 309622 3978
rect 309678 3922 327250 3978
rect 327306 3922 327374 3978
rect 327430 3922 327498 3978
rect 327554 3922 327622 3978
rect 327678 3922 345250 3978
rect 345306 3922 345374 3978
rect 345430 3922 345498 3978
rect 345554 3922 345622 3978
rect 345678 3922 363250 3978
rect 363306 3922 363374 3978
rect 363430 3922 363498 3978
rect 363554 3922 363622 3978
rect 363678 3922 381250 3978
rect 381306 3922 381374 3978
rect 381430 3922 381498 3978
rect 381554 3922 381622 3978
rect 381678 3922 399250 3978
rect 399306 3922 399374 3978
rect 399430 3922 399498 3978
rect 399554 3922 399622 3978
rect 399678 3922 417250 3978
rect 417306 3922 417374 3978
rect 417430 3922 417498 3978
rect 417554 3922 417622 3978
rect 417678 3922 435250 3978
rect 435306 3922 435374 3978
rect 435430 3922 435498 3978
rect 435554 3922 435622 3978
rect 435678 3922 453250 3978
rect 453306 3922 453374 3978
rect 453430 3922 453498 3978
rect 453554 3922 453622 3978
rect 453678 3922 471250 3978
rect 471306 3922 471374 3978
rect 471430 3922 471498 3978
rect 471554 3922 471622 3978
rect 471678 3922 489250 3978
rect 489306 3922 489374 3978
rect 489430 3922 489498 3978
rect 489554 3922 489622 3978
rect 489678 3922 507250 3978
rect 507306 3922 507374 3978
rect 507430 3922 507498 3978
rect 507554 3922 507622 3978
rect 507678 3922 525250 3978
rect 525306 3922 525374 3978
rect 525430 3922 525498 3978
rect 525554 3922 525622 3978
rect 525678 3922 543250 3978
rect 543306 3922 543374 3978
rect 543430 3922 543498 3978
rect 543554 3922 543622 3978
rect 543678 3922 561250 3978
rect 561306 3922 561374 3978
rect 561430 3922 561498 3978
rect 561554 3922 561622 3978
rect 561678 3922 579250 3978
rect 579306 3922 579374 3978
rect 579430 3922 579498 3978
rect 579554 3922 579622 3978
rect 579678 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 3250 -160
rect 3306 -216 3374 -160
rect 3430 -216 3498 -160
rect 3554 -216 3622 -160
rect 3678 -216 21250 -160
rect 21306 -216 21374 -160
rect 21430 -216 21498 -160
rect 21554 -216 21622 -160
rect 21678 -216 39250 -160
rect 39306 -216 39374 -160
rect 39430 -216 39498 -160
rect 39554 -216 39622 -160
rect 39678 -216 57250 -160
rect 57306 -216 57374 -160
rect 57430 -216 57498 -160
rect 57554 -216 57622 -160
rect 57678 -216 75250 -160
rect 75306 -216 75374 -160
rect 75430 -216 75498 -160
rect 75554 -216 75622 -160
rect 75678 -216 93250 -160
rect 93306 -216 93374 -160
rect 93430 -216 93498 -160
rect 93554 -216 93622 -160
rect 93678 -216 111250 -160
rect 111306 -216 111374 -160
rect 111430 -216 111498 -160
rect 111554 -216 111622 -160
rect 111678 -216 129250 -160
rect 129306 -216 129374 -160
rect 129430 -216 129498 -160
rect 129554 -216 129622 -160
rect 129678 -216 147250 -160
rect 147306 -216 147374 -160
rect 147430 -216 147498 -160
rect 147554 -216 147622 -160
rect 147678 -216 165250 -160
rect 165306 -216 165374 -160
rect 165430 -216 165498 -160
rect 165554 -216 165622 -160
rect 165678 -216 183250 -160
rect 183306 -216 183374 -160
rect 183430 -216 183498 -160
rect 183554 -216 183622 -160
rect 183678 -216 201250 -160
rect 201306 -216 201374 -160
rect 201430 -216 201498 -160
rect 201554 -216 201622 -160
rect 201678 -216 219250 -160
rect 219306 -216 219374 -160
rect 219430 -216 219498 -160
rect 219554 -216 219622 -160
rect 219678 -216 237250 -160
rect 237306 -216 237374 -160
rect 237430 -216 237498 -160
rect 237554 -216 237622 -160
rect 237678 -216 255250 -160
rect 255306 -216 255374 -160
rect 255430 -216 255498 -160
rect 255554 -216 255622 -160
rect 255678 -216 273250 -160
rect 273306 -216 273374 -160
rect 273430 -216 273498 -160
rect 273554 -216 273622 -160
rect 273678 -216 291250 -160
rect 291306 -216 291374 -160
rect 291430 -216 291498 -160
rect 291554 -216 291622 -160
rect 291678 -216 309250 -160
rect 309306 -216 309374 -160
rect 309430 -216 309498 -160
rect 309554 -216 309622 -160
rect 309678 -216 327250 -160
rect 327306 -216 327374 -160
rect 327430 -216 327498 -160
rect 327554 -216 327622 -160
rect 327678 -216 345250 -160
rect 345306 -216 345374 -160
rect 345430 -216 345498 -160
rect 345554 -216 345622 -160
rect 345678 -216 363250 -160
rect 363306 -216 363374 -160
rect 363430 -216 363498 -160
rect 363554 -216 363622 -160
rect 363678 -216 381250 -160
rect 381306 -216 381374 -160
rect 381430 -216 381498 -160
rect 381554 -216 381622 -160
rect 381678 -216 399250 -160
rect 399306 -216 399374 -160
rect 399430 -216 399498 -160
rect 399554 -216 399622 -160
rect 399678 -216 417250 -160
rect 417306 -216 417374 -160
rect 417430 -216 417498 -160
rect 417554 -216 417622 -160
rect 417678 -216 435250 -160
rect 435306 -216 435374 -160
rect 435430 -216 435498 -160
rect 435554 -216 435622 -160
rect 435678 -216 453250 -160
rect 453306 -216 453374 -160
rect 453430 -216 453498 -160
rect 453554 -216 453622 -160
rect 453678 -216 471250 -160
rect 471306 -216 471374 -160
rect 471430 -216 471498 -160
rect 471554 -216 471622 -160
rect 471678 -216 489250 -160
rect 489306 -216 489374 -160
rect 489430 -216 489498 -160
rect 489554 -216 489622 -160
rect 489678 -216 507250 -160
rect 507306 -216 507374 -160
rect 507430 -216 507498 -160
rect 507554 -216 507622 -160
rect 507678 -216 525250 -160
rect 525306 -216 525374 -160
rect 525430 -216 525498 -160
rect 525554 -216 525622 -160
rect 525678 -216 543250 -160
rect 543306 -216 543374 -160
rect 543430 -216 543498 -160
rect 543554 -216 543622 -160
rect 543678 -216 561250 -160
rect 561306 -216 561374 -160
rect 561430 -216 561498 -160
rect 561554 -216 561622 -160
rect 561678 -216 579250 -160
rect 579306 -216 579374 -160
rect 579430 -216 579498 -160
rect 579554 -216 579622 -160
rect 579678 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 3250 -284
rect 3306 -340 3374 -284
rect 3430 -340 3498 -284
rect 3554 -340 3622 -284
rect 3678 -340 21250 -284
rect 21306 -340 21374 -284
rect 21430 -340 21498 -284
rect 21554 -340 21622 -284
rect 21678 -340 39250 -284
rect 39306 -340 39374 -284
rect 39430 -340 39498 -284
rect 39554 -340 39622 -284
rect 39678 -340 57250 -284
rect 57306 -340 57374 -284
rect 57430 -340 57498 -284
rect 57554 -340 57622 -284
rect 57678 -340 75250 -284
rect 75306 -340 75374 -284
rect 75430 -340 75498 -284
rect 75554 -340 75622 -284
rect 75678 -340 93250 -284
rect 93306 -340 93374 -284
rect 93430 -340 93498 -284
rect 93554 -340 93622 -284
rect 93678 -340 111250 -284
rect 111306 -340 111374 -284
rect 111430 -340 111498 -284
rect 111554 -340 111622 -284
rect 111678 -340 129250 -284
rect 129306 -340 129374 -284
rect 129430 -340 129498 -284
rect 129554 -340 129622 -284
rect 129678 -340 147250 -284
rect 147306 -340 147374 -284
rect 147430 -340 147498 -284
rect 147554 -340 147622 -284
rect 147678 -340 165250 -284
rect 165306 -340 165374 -284
rect 165430 -340 165498 -284
rect 165554 -340 165622 -284
rect 165678 -340 183250 -284
rect 183306 -340 183374 -284
rect 183430 -340 183498 -284
rect 183554 -340 183622 -284
rect 183678 -340 201250 -284
rect 201306 -340 201374 -284
rect 201430 -340 201498 -284
rect 201554 -340 201622 -284
rect 201678 -340 219250 -284
rect 219306 -340 219374 -284
rect 219430 -340 219498 -284
rect 219554 -340 219622 -284
rect 219678 -340 237250 -284
rect 237306 -340 237374 -284
rect 237430 -340 237498 -284
rect 237554 -340 237622 -284
rect 237678 -340 255250 -284
rect 255306 -340 255374 -284
rect 255430 -340 255498 -284
rect 255554 -340 255622 -284
rect 255678 -340 273250 -284
rect 273306 -340 273374 -284
rect 273430 -340 273498 -284
rect 273554 -340 273622 -284
rect 273678 -340 291250 -284
rect 291306 -340 291374 -284
rect 291430 -340 291498 -284
rect 291554 -340 291622 -284
rect 291678 -340 309250 -284
rect 309306 -340 309374 -284
rect 309430 -340 309498 -284
rect 309554 -340 309622 -284
rect 309678 -340 327250 -284
rect 327306 -340 327374 -284
rect 327430 -340 327498 -284
rect 327554 -340 327622 -284
rect 327678 -340 345250 -284
rect 345306 -340 345374 -284
rect 345430 -340 345498 -284
rect 345554 -340 345622 -284
rect 345678 -340 363250 -284
rect 363306 -340 363374 -284
rect 363430 -340 363498 -284
rect 363554 -340 363622 -284
rect 363678 -340 381250 -284
rect 381306 -340 381374 -284
rect 381430 -340 381498 -284
rect 381554 -340 381622 -284
rect 381678 -340 399250 -284
rect 399306 -340 399374 -284
rect 399430 -340 399498 -284
rect 399554 -340 399622 -284
rect 399678 -340 417250 -284
rect 417306 -340 417374 -284
rect 417430 -340 417498 -284
rect 417554 -340 417622 -284
rect 417678 -340 435250 -284
rect 435306 -340 435374 -284
rect 435430 -340 435498 -284
rect 435554 -340 435622 -284
rect 435678 -340 453250 -284
rect 453306 -340 453374 -284
rect 453430 -340 453498 -284
rect 453554 -340 453622 -284
rect 453678 -340 471250 -284
rect 471306 -340 471374 -284
rect 471430 -340 471498 -284
rect 471554 -340 471622 -284
rect 471678 -340 489250 -284
rect 489306 -340 489374 -284
rect 489430 -340 489498 -284
rect 489554 -340 489622 -284
rect 489678 -340 507250 -284
rect 507306 -340 507374 -284
rect 507430 -340 507498 -284
rect 507554 -340 507622 -284
rect 507678 -340 525250 -284
rect 525306 -340 525374 -284
rect 525430 -340 525498 -284
rect 525554 -340 525622 -284
rect 525678 -340 543250 -284
rect 543306 -340 543374 -284
rect 543430 -340 543498 -284
rect 543554 -340 543622 -284
rect 543678 -340 561250 -284
rect 561306 -340 561374 -284
rect 561430 -340 561498 -284
rect 561554 -340 561622 -284
rect 561678 -340 579250 -284
rect 579306 -340 579374 -284
rect 579430 -340 579498 -284
rect 579554 -340 579622 -284
rect 579678 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 3250 -408
rect 3306 -464 3374 -408
rect 3430 -464 3498 -408
rect 3554 -464 3622 -408
rect 3678 -464 21250 -408
rect 21306 -464 21374 -408
rect 21430 -464 21498 -408
rect 21554 -464 21622 -408
rect 21678 -464 39250 -408
rect 39306 -464 39374 -408
rect 39430 -464 39498 -408
rect 39554 -464 39622 -408
rect 39678 -464 57250 -408
rect 57306 -464 57374 -408
rect 57430 -464 57498 -408
rect 57554 -464 57622 -408
rect 57678 -464 75250 -408
rect 75306 -464 75374 -408
rect 75430 -464 75498 -408
rect 75554 -464 75622 -408
rect 75678 -464 93250 -408
rect 93306 -464 93374 -408
rect 93430 -464 93498 -408
rect 93554 -464 93622 -408
rect 93678 -464 111250 -408
rect 111306 -464 111374 -408
rect 111430 -464 111498 -408
rect 111554 -464 111622 -408
rect 111678 -464 129250 -408
rect 129306 -464 129374 -408
rect 129430 -464 129498 -408
rect 129554 -464 129622 -408
rect 129678 -464 147250 -408
rect 147306 -464 147374 -408
rect 147430 -464 147498 -408
rect 147554 -464 147622 -408
rect 147678 -464 165250 -408
rect 165306 -464 165374 -408
rect 165430 -464 165498 -408
rect 165554 -464 165622 -408
rect 165678 -464 183250 -408
rect 183306 -464 183374 -408
rect 183430 -464 183498 -408
rect 183554 -464 183622 -408
rect 183678 -464 201250 -408
rect 201306 -464 201374 -408
rect 201430 -464 201498 -408
rect 201554 -464 201622 -408
rect 201678 -464 219250 -408
rect 219306 -464 219374 -408
rect 219430 -464 219498 -408
rect 219554 -464 219622 -408
rect 219678 -464 237250 -408
rect 237306 -464 237374 -408
rect 237430 -464 237498 -408
rect 237554 -464 237622 -408
rect 237678 -464 255250 -408
rect 255306 -464 255374 -408
rect 255430 -464 255498 -408
rect 255554 -464 255622 -408
rect 255678 -464 273250 -408
rect 273306 -464 273374 -408
rect 273430 -464 273498 -408
rect 273554 -464 273622 -408
rect 273678 -464 291250 -408
rect 291306 -464 291374 -408
rect 291430 -464 291498 -408
rect 291554 -464 291622 -408
rect 291678 -464 309250 -408
rect 309306 -464 309374 -408
rect 309430 -464 309498 -408
rect 309554 -464 309622 -408
rect 309678 -464 327250 -408
rect 327306 -464 327374 -408
rect 327430 -464 327498 -408
rect 327554 -464 327622 -408
rect 327678 -464 345250 -408
rect 345306 -464 345374 -408
rect 345430 -464 345498 -408
rect 345554 -464 345622 -408
rect 345678 -464 363250 -408
rect 363306 -464 363374 -408
rect 363430 -464 363498 -408
rect 363554 -464 363622 -408
rect 363678 -464 381250 -408
rect 381306 -464 381374 -408
rect 381430 -464 381498 -408
rect 381554 -464 381622 -408
rect 381678 -464 399250 -408
rect 399306 -464 399374 -408
rect 399430 -464 399498 -408
rect 399554 -464 399622 -408
rect 399678 -464 417250 -408
rect 417306 -464 417374 -408
rect 417430 -464 417498 -408
rect 417554 -464 417622 -408
rect 417678 -464 435250 -408
rect 435306 -464 435374 -408
rect 435430 -464 435498 -408
rect 435554 -464 435622 -408
rect 435678 -464 453250 -408
rect 453306 -464 453374 -408
rect 453430 -464 453498 -408
rect 453554 -464 453622 -408
rect 453678 -464 471250 -408
rect 471306 -464 471374 -408
rect 471430 -464 471498 -408
rect 471554 -464 471622 -408
rect 471678 -464 489250 -408
rect 489306 -464 489374 -408
rect 489430 -464 489498 -408
rect 489554 -464 489622 -408
rect 489678 -464 507250 -408
rect 507306 -464 507374 -408
rect 507430 -464 507498 -408
rect 507554 -464 507622 -408
rect 507678 -464 525250 -408
rect 525306 -464 525374 -408
rect 525430 -464 525498 -408
rect 525554 -464 525622 -408
rect 525678 -464 543250 -408
rect 543306 -464 543374 -408
rect 543430 -464 543498 -408
rect 543554 -464 543622 -408
rect 543678 -464 561250 -408
rect 561306 -464 561374 -408
rect 561430 -464 561498 -408
rect 561554 -464 561622 -408
rect 561678 -464 579250 -408
rect 579306 -464 579374 -408
rect 579430 -464 579498 -408
rect 579554 -464 579622 -408
rect 579678 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 3250 -532
rect 3306 -588 3374 -532
rect 3430 -588 3498 -532
rect 3554 -588 3622 -532
rect 3678 -588 21250 -532
rect 21306 -588 21374 -532
rect 21430 -588 21498 -532
rect 21554 -588 21622 -532
rect 21678 -588 39250 -532
rect 39306 -588 39374 -532
rect 39430 -588 39498 -532
rect 39554 -588 39622 -532
rect 39678 -588 57250 -532
rect 57306 -588 57374 -532
rect 57430 -588 57498 -532
rect 57554 -588 57622 -532
rect 57678 -588 75250 -532
rect 75306 -588 75374 -532
rect 75430 -588 75498 -532
rect 75554 -588 75622 -532
rect 75678 -588 93250 -532
rect 93306 -588 93374 -532
rect 93430 -588 93498 -532
rect 93554 -588 93622 -532
rect 93678 -588 111250 -532
rect 111306 -588 111374 -532
rect 111430 -588 111498 -532
rect 111554 -588 111622 -532
rect 111678 -588 129250 -532
rect 129306 -588 129374 -532
rect 129430 -588 129498 -532
rect 129554 -588 129622 -532
rect 129678 -588 147250 -532
rect 147306 -588 147374 -532
rect 147430 -588 147498 -532
rect 147554 -588 147622 -532
rect 147678 -588 165250 -532
rect 165306 -588 165374 -532
rect 165430 -588 165498 -532
rect 165554 -588 165622 -532
rect 165678 -588 183250 -532
rect 183306 -588 183374 -532
rect 183430 -588 183498 -532
rect 183554 -588 183622 -532
rect 183678 -588 201250 -532
rect 201306 -588 201374 -532
rect 201430 -588 201498 -532
rect 201554 -588 201622 -532
rect 201678 -588 219250 -532
rect 219306 -588 219374 -532
rect 219430 -588 219498 -532
rect 219554 -588 219622 -532
rect 219678 -588 237250 -532
rect 237306 -588 237374 -532
rect 237430 -588 237498 -532
rect 237554 -588 237622 -532
rect 237678 -588 255250 -532
rect 255306 -588 255374 -532
rect 255430 -588 255498 -532
rect 255554 -588 255622 -532
rect 255678 -588 273250 -532
rect 273306 -588 273374 -532
rect 273430 -588 273498 -532
rect 273554 -588 273622 -532
rect 273678 -588 291250 -532
rect 291306 -588 291374 -532
rect 291430 -588 291498 -532
rect 291554 -588 291622 -532
rect 291678 -588 309250 -532
rect 309306 -588 309374 -532
rect 309430 -588 309498 -532
rect 309554 -588 309622 -532
rect 309678 -588 327250 -532
rect 327306 -588 327374 -532
rect 327430 -588 327498 -532
rect 327554 -588 327622 -532
rect 327678 -588 345250 -532
rect 345306 -588 345374 -532
rect 345430 -588 345498 -532
rect 345554 -588 345622 -532
rect 345678 -588 363250 -532
rect 363306 -588 363374 -532
rect 363430 -588 363498 -532
rect 363554 -588 363622 -532
rect 363678 -588 381250 -532
rect 381306 -588 381374 -532
rect 381430 -588 381498 -532
rect 381554 -588 381622 -532
rect 381678 -588 399250 -532
rect 399306 -588 399374 -532
rect 399430 -588 399498 -532
rect 399554 -588 399622 -532
rect 399678 -588 417250 -532
rect 417306 -588 417374 -532
rect 417430 -588 417498 -532
rect 417554 -588 417622 -532
rect 417678 -588 435250 -532
rect 435306 -588 435374 -532
rect 435430 -588 435498 -532
rect 435554 -588 435622 -532
rect 435678 -588 453250 -532
rect 453306 -588 453374 -532
rect 453430 -588 453498 -532
rect 453554 -588 453622 -532
rect 453678 -588 471250 -532
rect 471306 -588 471374 -532
rect 471430 -588 471498 -532
rect 471554 -588 471622 -532
rect 471678 -588 489250 -532
rect 489306 -588 489374 -532
rect 489430 -588 489498 -532
rect 489554 -588 489622 -532
rect 489678 -588 507250 -532
rect 507306 -588 507374 -532
rect 507430 -588 507498 -532
rect 507554 -588 507622 -532
rect 507678 -588 525250 -532
rect 525306 -588 525374 -532
rect 525430 -588 525498 -532
rect 525554 -588 525622 -532
rect 525678 -588 543250 -532
rect 543306 -588 543374 -532
rect 543430 -588 543498 -532
rect 543554 -588 543622 -532
rect 543678 -588 561250 -532
rect 561306 -588 561374 -532
rect 561430 -588 561498 -532
rect 561554 -588 561622 -532
rect 561678 -588 579250 -532
rect 579306 -588 579374 -532
rect 579430 -588 579498 -532
rect 579554 -588 579622 -532
rect 579678 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 6970 -1120
rect 7026 -1176 7094 -1120
rect 7150 -1176 7218 -1120
rect 7274 -1176 7342 -1120
rect 7398 -1176 24970 -1120
rect 25026 -1176 25094 -1120
rect 25150 -1176 25218 -1120
rect 25274 -1176 25342 -1120
rect 25398 -1176 42970 -1120
rect 43026 -1176 43094 -1120
rect 43150 -1176 43218 -1120
rect 43274 -1176 43342 -1120
rect 43398 -1176 60970 -1120
rect 61026 -1176 61094 -1120
rect 61150 -1176 61218 -1120
rect 61274 -1176 61342 -1120
rect 61398 -1176 78970 -1120
rect 79026 -1176 79094 -1120
rect 79150 -1176 79218 -1120
rect 79274 -1176 79342 -1120
rect 79398 -1176 96970 -1120
rect 97026 -1176 97094 -1120
rect 97150 -1176 97218 -1120
rect 97274 -1176 97342 -1120
rect 97398 -1176 114970 -1120
rect 115026 -1176 115094 -1120
rect 115150 -1176 115218 -1120
rect 115274 -1176 115342 -1120
rect 115398 -1176 132970 -1120
rect 133026 -1176 133094 -1120
rect 133150 -1176 133218 -1120
rect 133274 -1176 133342 -1120
rect 133398 -1176 150970 -1120
rect 151026 -1176 151094 -1120
rect 151150 -1176 151218 -1120
rect 151274 -1176 151342 -1120
rect 151398 -1176 168970 -1120
rect 169026 -1176 169094 -1120
rect 169150 -1176 169218 -1120
rect 169274 -1176 169342 -1120
rect 169398 -1176 186970 -1120
rect 187026 -1176 187094 -1120
rect 187150 -1176 187218 -1120
rect 187274 -1176 187342 -1120
rect 187398 -1176 204970 -1120
rect 205026 -1176 205094 -1120
rect 205150 -1176 205218 -1120
rect 205274 -1176 205342 -1120
rect 205398 -1176 222970 -1120
rect 223026 -1176 223094 -1120
rect 223150 -1176 223218 -1120
rect 223274 -1176 223342 -1120
rect 223398 -1176 240970 -1120
rect 241026 -1176 241094 -1120
rect 241150 -1176 241218 -1120
rect 241274 -1176 241342 -1120
rect 241398 -1176 258970 -1120
rect 259026 -1176 259094 -1120
rect 259150 -1176 259218 -1120
rect 259274 -1176 259342 -1120
rect 259398 -1176 276970 -1120
rect 277026 -1176 277094 -1120
rect 277150 -1176 277218 -1120
rect 277274 -1176 277342 -1120
rect 277398 -1176 294970 -1120
rect 295026 -1176 295094 -1120
rect 295150 -1176 295218 -1120
rect 295274 -1176 295342 -1120
rect 295398 -1176 312970 -1120
rect 313026 -1176 313094 -1120
rect 313150 -1176 313218 -1120
rect 313274 -1176 313342 -1120
rect 313398 -1176 330970 -1120
rect 331026 -1176 331094 -1120
rect 331150 -1176 331218 -1120
rect 331274 -1176 331342 -1120
rect 331398 -1176 348970 -1120
rect 349026 -1176 349094 -1120
rect 349150 -1176 349218 -1120
rect 349274 -1176 349342 -1120
rect 349398 -1176 366970 -1120
rect 367026 -1176 367094 -1120
rect 367150 -1176 367218 -1120
rect 367274 -1176 367342 -1120
rect 367398 -1176 384970 -1120
rect 385026 -1176 385094 -1120
rect 385150 -1176 385218 -1120
rect 385274 -1176 385342 -1120
rect 385398 -1176 402970 -1120
rect 403026 -1176 403094 -1120
rect 403150 -1176 403218 -1120
rect 403274 -1176 403342 -1120
rect 403398 -1176 420970 -1120
rect 421026 -1176 421094 -1120
rect 421150 -1176 421218 -1120
rect 421274 -1176 421342 -1120
rect 421398 -1176 438970 -1120
rect 439026 -1176 439094 -1120
rect 439150 -1176 439218 -1120
rect 439274 -1176 439342 -1120
rect 439398 -1176 456970 -1120
rect 457026 -1176 457094 -1120
rect 457150 -1176 457218 -1120
rect 457274 -1176 457342 -1120
rect 457398 -1176 474970 -1120
rect 475026 -1176 475094 -1120
rect 475150 -1176 475218 -1120
rect 475274 -1176 475342 -1120
rect 475398 -1176 492970 -1120
rect 493026 -1176 493094 -1120
rect 493150 -1176 493218 -1120
rect 493274 -1176 493342 -1120
rect 493398 -1176 510970 -1120
rect 511026 -1176 511094 -1120
rect 511150 -1176 511218 -1120
rect 511274 -1176 511342 -1120
rect 511398 -1176 528970 -1120
rect 529026 -1176 529094 -1120
rect 529150 -1176 529218 -1120
rect 529274 -1176 529342 -1120
rect 529398 -1176 546970 -1120
rect 547026 -1176 547094 -1120
rect 547150 -1176 547218 -1120
rect 547274 -1176 547342 -1120
rect 547398 -1176 564970 -1120
rect 565026 -1176 565094 -1120
rect 565150 -1176 565218 -1120
rect 565274 -1176 565342 -1120
rect 565398 -1176 582970 -1120
rect 583026 -1176 583094 -1120
rect 583150 -1176 583218 -1120
rect 583274 -1176 583342 -1120
rect 583398 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 6970 -1244
rect 7026 -1300 7094 -1244
rect 7150 -1300 7218 -1244
rect 7274 -1300 7342 -1244
rect 7398 -1300 24970 -1244
rect 25026 -1300 25094 -1244
rect 25150 -1300 25218 -1244
rect 25274 -1300 25342 -1244
rect 25398 -1300 42970 -1244
rect 43026 -1300 43094 -1244
rect 43150 -1300 43218 -1244
rect 43274 -1300 43342 -1244
rect 43398 -1300 60970 -1244
rect 61026 -1300 61094 -1244
rect 61150 -1300 61218 -1244
rect 61274 -1300 61342 -1244
rect 61398 -1300 78970 -1244
rect 79026 -1300 79094 -1244
rect 79150 -1300 79218 -1244
rect 79274 -1300 79342 -1244
rect 79398 -1300 96970 -1244
rect 97026 -1300 97094 -1244
rect 97150 -1300 97218 -1244
rect 97274 -1300 97342 -1244
rect 97398 -1300 114970 -1244
rect 115026 -1300 115094 -1244
rect 115150 -1300 115218 -1244
rect 115274 -1300 115342 -1244
rect 115398 -1300 132970 -1244
rect 133026 -1300 133094 -1244
rect 133150 -1300 133218 -1244
rect 133274 -1300 133342 -1244
rect 133398 -1300 150970 -1244
rect 151026 -1300 151094 -1244
rect 151150 -1300 151218 -1244
rect 151274 -1300 151342 -1244
rect 151398 -1300 168970 -1244
rect 169026 -1300 169094 -1244
rect 169150 -1300 169218 -1244
rect 169274 -1300 169342 -1244
rect 169398 -1300 186970 -1244
rect 187026 -1300 187094 -1244
rect 187150 -1300 187218 -1244
rect 187274 -1300 187342 -1244
rect 187398 -1300 204970 -1244
rect 205026 -1300 205094 -1244
rect 205150 -1300 205218 -1244
rect 205274 -1300 205342 -1244
rect 205398 -1300 222970 -1244
rect 223026 -1300 223094 -1244
rect 223150 -1300 223218 -1244
rect 223274 -1300 223342 -1244
rect 223398 -1300 240970 -1244
rect 241026 -1300 241094 -1244
rect 241150 -1300 241218 -1244
rect 241274 -1300 241342 -1244
rect 241398 -1300 258970 -1244
rect 259026 -1300 259094 -1244
rect 259150 -1300 259218 -1244
rect 259274 -1300 259342 -1244
rect 259398 -1300 276970 -1244
rect 277026 -1300 277094 -1244
rect 277150 -1300 277218 -1244
rect 277274 -1300 277342 -1244
rect 277398 -1300 294970 -1244
rect 295026 -1300 295094 -1244
rect 295150 -1300 295218 -1244
rect 295274 -1300 295342 -1244
rect 295398 -1300 312970 -1244
rect 313026 -1300 313094 -1244
rect 313150 -1300 313218 -1244
rect 313274 -1300 313342 -1244
rect 313398 -1300 330970 -1244
rect 331026 -1300 331094 -1244
rect 331150 -1300 331218 -1244
rect 331274 -1300 331342 -1244
rect 331398 -1300 348970 -1244
rect 349026 -1300 349094 -1244
rect 349150 -1300 349218 -1244
rect 349274 -1300 349342 -1244
rect 349398 -1300 366970 -1244
rect 367026 -1300 367094 -1244
rect 367150 -1300 367218 -1244
rect 367274 -1300 367342 -1244
rect 367398 -1300 384970 -1244
rect 385026 -1300 385094 -1244
rect 385150 -1300 385218 -1244
rect 385274 -1300 385342 -1244
rect 385398 -1300 402970 -1244
rect 403026 -1300 403094 -1244
rect 403150 -1300 403218 -1244
rect 403274 -1300 403342 -1244
rect 403398 -1300 420970 -1244
rect 421026 -1300 421094 -1244
rect 421150 -1300 421218 -1244
rect 421274 -1300 421342 -1244
rect 421398 -1300 438970 -1244
rect 439026 -1300 439094 -1244
rect 439150 -1300 439218 -1244
rect 439274 -1300 439342 -1244
rect 439398 -1300 456970 -1244
rect 457026 -1300 457094 -1244
rect 457150 -1300 457218 -1244
rect 457274 -1300 457342 -1244
rect 457398 -1300 474970 -1244
rect 475026 -1300 475094 -1244
rect 475150 -1300 475218 -1244
rect 475274 -1300 475342 -1244
rect 475398 -1300 492970 -1244
rect 493026 -1300 493094 -1244
rect 493150 -1300 493218 -1244
rect 493274 -1300 493342 -1244
rect 493398 -1300 510970 -1244
rect 511026 -1300 511094 -1244
rect 511150 -1300 511218 -1244
rect 511274 -1300 511342 -1244
rect 511398 -1300 528970 -1244
rect 529026 -1300 529094 -1244
rect 529150 -1300 529218 -1244
rect 529274 -1300 529342 -1244
rect 529398 -1300 546970 -1244
rect 547026 -1300 547094 -1244
rect 547150 -1300 547218 -1244
rect 547274 -1300 547342 -1244
rect 547398 -1300 564970 -1244
rect 565026 -1300 565094 -1244
rect 565150 -1300 565218 -1244
rect 565274 -1300 565342 -1244
rect 565398 -1300 582970 -1244
rect 583026 -1300 583094 -1244
rect 583150 -1300 583218 -1244
rect 583274 -1300 583342 -1244
rect 583398 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 6970 -1368
rect 7026 -1424 7094 -1368
rect 7150 -1424 7218 -1368
rect 7274 -1424 7342 -1368
rect 7398 -1424 24970 -1368
rect 25026 -1424 25094 -1368
rect 25150 -1424 25218 -1368
rect 25274 -1424 25342 -1368
rect 25398 -1424 42970 -1368
rect 43026 -1424 43094 -1368
rect 43150 -1424 43218 -1368
rect 43274 -1424 43342 -1368
rect 43398 -1424 60970 -1368
rect 61026 -1424 61094 -1368
rect 61150 -1424 61218 -1368
rect 61274 -1424 61342 -1368
rect 61398 -1424 78970 -1368
rect 79026 -1424 79094 -1368
rect 79150 -1424 79218 -1368
rect 79274 -1424 79342 -1368
rect 79398 -1424 96970 -1368
rect 97026 -1424 97094 -1368
rect 97150 -1424 97218 -1368
rect 97274 -1424 97342 -1368
rect 97398 -1424 114970 -1368
rect 115026 -1424 115094 -1368
rect 115150 -1424 115218 -1368
rect 115274 -1424 115342 -1368
rect 115398 -1424 132970 -1368
rect 133026 -1424 133094 -1368
rect 133150 -1424 133218 -1368
rect 133274 -1424 133342 -1368
rect 133398 -1424 150970 -1368
rect 151026 -1424 151094 -1368
rect 151150 -1424 151218 -1368
rect 151274 -1424 151342 -1368
rect 151398 -1424 168970 -1368
rect 169026 -1424 169094 -1368
rect 169150 -1424 169218 -1368
rect 169274 -1424 169342 -1368
rect 169398 -1424 186970 -1368
rect 187026 -1424 187094 -1368
rect 187150 -1424 187218 -1368
rect 187274 -1424 187342 -1368
rect 187398 -1424 204970 -1368
rect 205026 -1424 205094 -1368
rect 205150 -1424 205218 -1368
rect 205274 -1424 205342 -1368
rect 205398 -1424 222970 -1368
rect 223026 -1424 223094 -1368
rect 223150 -1424 223218 -1368
rect 223274 -1424 223342 -1368
rect 223398 -1424 240970 -1368
rect 241026 -1424 241094 -1368
rect 241150 -1424 241218 -1368
rect 241274 -1424 241342 -1368
rect 241398 -1424 258970 -1368
rect 259026 -1424 259094 -1368
rect 259150 -1424 259218 -1368
rect 259274 -1424 259342 -1368
rect 259398 -1424 276970 -1368
rect 277026 -1424 277094 -1368
rect 277150 -1424 277218 -1368
rect 277274 -1424 277342 -1368
rect 277398 -1424 294970 -1368
rect 295026 -1424 295094 -1368
rect 295150 -1424 295218 -1368
rect 295274 -1424 295342 -1368
rect 295398 -1424 312970 -1368
rect 313026 -1424 313094 -1368
rect 313150 -1424 313218 -1368
rect 313274 -1424 313342 -1368
rect 313398 -1424 330970 -1368
rect 331026 -1424 331094 -1368
rect 331150 -1424 331218 -1368
rect 331274 -1424 331342 -1368
rect 331398 -1424 348970 -1368
rect 349026 -1424 349094 -1368
rect 349150 -1424 349218 -1368
rect 349274 -1424 349342 -1368
rect 349398 -1424 366970 -1368
rect 367026 -1424 367094 -1368
rect 367150 -1424 367218 -1368
rect 367274 -1424 367342 -1368
rect 367398 -1424 384970 -1368
rect 385026 -1424 385094 -1368
rect 385150 -1424 385218 -1368
rect 385274 -1424 385342 -1368
rect 385398 -1424 402970 -1368
rect 403026 -1424 403094 -1368
rect 403150 -1424 403218 -1368
rect 403274 -1424 403342 -1368
rect 403398 -1424 420970 -1368
rect 421026 -1424 421094 -1368
rect 421150 -1424 421218 -1368
rect 421274 -1424 421342 -1368
rect 421398 -1424 438970 -1368
rect 439026 -1424 439094 -1368
rect 439150 -1424 439218 -1368
rect 439274 -1424 439342 -1368
rect 439398 -1424 456970 -1368
rect 457026 -1424 457094 -1368
rect 457150 -1424 457218 -1368
rect 457274 -1424 457342 -1368
rect 457398 -1424 474970 -1368
rect 475026 -1424 475094 -1368
rect 475150 -1424 475218 -1368
rect 475274 -1424 475342 -1368
rect 475398 -1424 492970 -1368
rect 493026 -1424 493094 -1368
rect 493150 -1424 493218 -1368
rect 493274 -1424 493342 -1368
rect 493398 -1424 510970 -1368
rect 511026 -1424 511094 -1368
rect 511150 -1424 511218 -1368
rect 511274 -1424 511342 -1368
rect 511398 -1424 528970 -1368
rect 529026 -1424 529094 -1368
rect 529150 -1424 529218 -1368
rect 529274 -1424 529342 -1368
rect 529398 -1424 546970 -1368
rect 547026 -1424 547094 -1368
rect 547150 -1424 547218 -1368
rect 547274 -1424 547342 -1368
rect 547398 -1424 564970 -1368
rect 565026 -1424 565094 -1368
rect 565150 -1424 565218 -1368
rect 565274 -1424 565342 -1368
rect 565398 -1424 582970 -1368
rect 583026 -1424 583094 -1368
rect 583150 -1424 583218 -1368
rect 583274 -1424 583342 -1368
rect 583398 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 6970 -1492
rect 7026 -1548 7094 -1492
rect 7150 -1548 7218 -1492
rect 7274 -1548 7342 -1492
rect 7398 -1548 24970 -1492
rect 25026 -1548 25094 -1492
rect 25150 -1548 25218 -1492
rect 25274 -1548 25342 -1492
rect 25398 -1548 42970 -1492
rect 43026 -1548 43094 -1492
rect 43150 -1548 43218 -1492
rect 43274 -1548 43342 -1492
rect 43398 -1548 60970 -1492
rect 61026 -1548 61094 -1492
rect 61150 -1548 61218 -1492
rect 61274 -1548 61342 -1492
rect 61398 -1548 78970 -1492
rect 79026 -1548 79094 -1492
rect 79150 -1548 79218 -1492
rect 79274 -1548 79342 -1492
rect 79398 -1548 96970 -1492
rect 97026 -1548 97094 -1492
rect 97150 -1548 97218 -1492
rect 97274 -1548 97342 -1492
rect 97398 -1548 114970 -1492
rect 115026 -1548 115094 -1492
rect 115150 -1548 115218 -1492
rect 115274 -1548 115342 -1492
rect 115398 -1548 132970 -1492
rect 133026 -1548 133094 -1492
rect 133150 -1548 133218 -1492
rect 133274 -1548 133342 -1492
rect 133398 -1548 150970 -1492
rect 151026 -1548 151094 -1492
rect 151150 -1548 151218 -1492
rect 151274 -1548 151342 -1492
rect 151398 -1548 168970 -1492
rect 169026 -1548 169094 -1492
rect 169150 -1548 169218 -1492
rect 169274 -1548 169342 -1492
rect 169398 -1548 186970 -1492
rect 187026 -1548 187094 -1492
rect 187150 -1548 187218 -1492
rect 187274 -1548 187342 -1492
rect 187398 -1548 204970 -1492
rect 205026 -1548 205094 -1492
rect 205150 -1548 205218 -1492
rect 205274 -1548 205342 -1492
rect 205398 -1548 222970 -1492
rect 223026 -1548 223094 -1492
rect 223150 -1548 223218 -1492
rect 223274 -1548 223342 -1492
rect 223398 -1548 240970 -1492
rect 241026 -1548 241094 -1492
rect 241150 -1548 241218 -1492
rect 241274 -1548 241342 -1492
rect 241398 -1548 258970 -1492
rect 259026 -1548 259094 -1492
rect 259150 -1548 259218 -1492
rect 259274 -1548 259342 -1492
rect 259398 -1548 276970 -1492
rect 277026 -1548 277094 -1492
rect 277150 -1548 277218 -1492
rect 277274 -1548 277342 -1492
rect 277398 -1548 294970 -1492
rect 295026 -1548 295094 -1492
rect 295150 -1548 295218 -1492
rect 295274 -1548 295342 -1492
rect 295398 -1548 312970 -1492
rect 313026 -1548 313094 -1492
rect 313150 -1548 313218 -1492
rect 313274 -1548 313342 -1492
rect 313398 -1548 330970 -1492
rect 331026 -1548 331094 -1492
rect 331150 -1548 331218 -1492
rect 331274 -1548 331342 -1492
rect 331398 -1548 348970 -1492
rect 349026 -1548 349094 -1492
rect 349150 -1548 349218 -1492
rect 349274 -1548 349342 -1492
rect 349398 -1548 366970 -1492
rect 367026 -1548 367094 -1492
rect 367150 -1548 367218 -1492
rect 367274 -1548 367342 -1492
rect 367398 -1548 384970 -1492
rect 385026 -1548 385094 -1492
rect 385150 -1548 385218 -1492
rect 385274 -1548 385342 -1492
rect 385398 -1548 402970 -1492
rect 403026 -1548 403094 -1492
rect 403150 -1548 403218 -1492
rect 403274 -1548 403342 -1492
rect 403398 -1548 420970 -1492
rect 421026 -1548 421094 -1492
rect 421150 -1548 421218 -1492
rect 421274 -1548 421342 -1492
rect 421398 -1548 438970 -1492
rect 439026 -1548 439094 -1492
rect 439150 -1548 439218 -1492
rect 439274 -1548 439342 -1492
rect 439398 -1548 456970 -1492
rect 457026 -1548 457094 -1492
rect 457150 -1548 457218 -1492
rect 457274 -1548 457342 -1492
rect 457398 -1548 474970 -1492
rect 475026 -1548 475094 -1492
rect 475150 -1548 475218 -1492
rect 475274 -1548 475342 -1492
rect 475398 -1548 492970 -1492
rect 493026 -1548 493094 -1492
rect 493150 -1548 493218 -1492
rect 493274 -1548 493342 -1492
rect 493398 -1548 510970 -1492
rect 511026 -1548 511094 -1492
rect 511150 -1548 511218 -1492
rect 511274 -1548 511342 -1492
rect 511398 -1548 528970 -1492
rect 529026 -1548 529094 -1492
rect 529150 -1548 529218 -1492
rect 529274 -1548 529342 -1492
rect 529398 -1548 546970 -1492
rect 547026 -1548 547094 -1492
rect 547150 -1548 547218 -1492
rect 547274 -1548 547342 -1492
rect 547398 -1548 564970 -1492
rect 565026 -1548 565094 -1492
rect 565150 -1548 565218 -1492
rect 565274 -1548 565342 -1492
rect 565398 -1548 582970 -1492
rect 583026 -1548 583094 -1492
rect 583150 -1548 583218 -1492
rect 583274 -1548 583342 -1492
rect 583398 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use vb_wrapper  mprj
timestamp 0
transform 1 0 200000 0 1 200000
box 1344 0 298686 300000
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 3154 -1644 3774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 21154 -1644 21774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 39154 -1644 39774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 57154 -1644 57774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 75154 -1644 75774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 93154 -1644 93774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 111154 -1644 111774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 129154 -1644 129774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 147154 -1644 147774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 165154 -1644 165774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 183154 -1644 183774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 201154 -1644 201774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 -1644 219774 201020 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 219154 499846 219774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 -1644 237774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 237154 499846 237774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 -1644 255774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 255154 499846 255774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 -1644 273774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 273154 499846 273774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 -1644 291774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 291154 499846 291774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 -1644 309774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 309154 499846 309774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 -1644 327774 201020 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 327154 499846 327774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 -1644 345774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 345154 499846 345774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 -1644 363774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 363154 499846 363774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 -1644 381774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 381154 499846 381774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 -1644 399774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 399154 499846 399774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 -1644 417774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 417154 499846 417774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 -1644 435774 201020 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435154 499846 435774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 -1644 453774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 453154 499846 453774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 -1644 471774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 471154 499846 471774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 -1644 489774 210842 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 489154 499846 489774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 507154 -1644 507774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 525154 -1644 525774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 543154 -1644 543774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 561154 -1644 561774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 579154 -1644 579774 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 6874 -1644 7494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 24874 -1644 25494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 42874 -1644 43494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 60874 -1644 61494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 78874 -1644 79494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 96874 -1644 97494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 114874 -1644 115494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132874 -1644 133494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 150874 -1644 151494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 168874 -1644 169494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 186874 -1644 187494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 -1644 205494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 204874 499846 205494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 -1644 223494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 222874 499846 223494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 -1644 241494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 240874 499846 241494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 -1644 259494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 258874 499846 259494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 -1644 277494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 276874 499846 277494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 -1644 295494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 294874 499846 295494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 -1644 313494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 312874 499846 313494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 -1644 331494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 330874 499846 331494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 -1644 349494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 348874 499846 349494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 -1644 367494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 366874 499846 367494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 -1644 385494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 384874 499846 385494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 -1644 403494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 402874 499846 403494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 -1644 421494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 420874 499846 421494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 -1644 439494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 438874 499846 439494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 -1644 457494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 456874 499846 457494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 -1644 475494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 474874 499846 475494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 -1644 493494 210842 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 492874 499846 493494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 510874 -1644 511494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 528874 -1644 529494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 546874 -1644 547494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 564874 -1644 565494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 582874 -1644 583494 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 489650 202322 489650 202322 0 vdd
rlabel via4 496510 496305 496510 496305 0 vss
rlabel metal3 594426 7336 594426 7336 0 io_in[0]
rlabel metal2 281330 499912 281330 499912 0 io_in[10]
rlabel metal2 289226 499912 289226 499912 0 io_in[11]
rlabel metal3 595098 483112 595098 483112 0 io_in[12]
rlabel metal2 304514 499912 304514 499912 0 io_in[13]
rlabel metal3 595672 561624 595672 561624 0 io_in[14]
rlabel metal3 589064 590184 589064 590184 0 io_in[15]
rlabel metal2 327866 499912 327866 499912 0 io_in[16]
rlabel metal2 335426 499912 335426 499912 0 io_in[17]
rlabel metal2 343154 499912 343154 499912 0 io_in[18]
rlabel metal2 351218 499912 351218 499912 0 io_in[19]
rlabel metal3 594538 46984 594538 46984 0 io_in[1]
rlabel metal2 358610 499912 358610 499912 0 io_in[20]
rlabel metal2 187768 594426 187768 594426 0 io_in[21]
rlabel metal2 374066 499912 374066 499912 0 io_in[22]
rlabel metal2 55384 594370 55384 594370 0 io_in[23]
rlabel metal3 392 586712 392 586712 0 io_in[24]
rlabel metal3 392 544544 392 544544 0 io_in[25]
rlabel metal2 405384 500710 405384 500710 0 io_in[26]
rlabel metal3 392 459368 392 459368 0 io_in[27]
rlabel metal2 420840 500486 420840 500486 0 io_in[28]
rlabel metal3 392 375032 392 375032 0 io_in[29]
rlabel metal2 219506 499912 219506 499912 0 io_in[2]
rlabel metal3 392 332864 392 332864 0 io_in[30]
rlabel metal2 443786 499912 443786 499912 0 io_in[31]
rlabel metal2 451346 499912 451346 499912 0 io_in[32]
rlabel metal2 459074 499912 459074 499912 0 io_in[33]
rlabel metal3 392 163352 392 163352 0 io_in[34]
rlabel metal3 392 121184 392 121184 0 io_in[35]
rlabel metal2 482664 500486 482664 500486 0 io_in[36]
rlabel metal3 2310 36904 2310 36904 0 io_in[37]
rlabel metal3 594706 126280 594706 126280 0 io_in[3]
rlabel metal2 235298 499912 235298 499912 0 io_in[4]
rlabel metal2 242690 499912 242690 499912 0 io_in[5]
rlabel metal3 594818 245224 594818 245224 0 io_in[6]
rlabel metal3 594874 284872 594874 284872 0 io_in[7]
rlabel metal3 594930 324520 594930 324520 0 io_in[8]
rlabel metal3 595672 363384 595672 363384 0 io_in[9]
rlabel metal3 594482 33768 594482 33768 0 io_oeb[0]
rlabel metal3 346276 499240 346276 499240 0 io_oeb[10]
rlabel metal3 595672 469168 595672 469168 0 io_oeb[11]
rlabel metal2 299418 499912 299418 499912 0 io_oeb[12]
rlabel metal3 595672 548296 595672 548296 0 io_oeb[13]
rlabel metal3 594370 588616 594370 588616 0 io_oeb[14]
rlabel metal2 539896 595672 539896 595672 0 io_oeb[15]
rlabel metal2 474040 595672 474040 595672 0 io_oeb[16]
rlabel metal2 338408 501774 338408 501774 0 io_oeb[17]
rlabel metal3 343616 521304 343616 521304 0 io_oeb[18]
rlabel metal2 353458 499912 353458 499912 0 io_oeb[19]
rlabel metal2 214354 499912 214354 499912 0 io_oeb[1]
rlabel metal2 208936 595672 208936 595672 0 io_oeb[20]
rlabel metal2 143640 590562 143640 590562 0 io_oeb[21]
rlabel metal2 376698 499912 376698 499912 0 io_oeb[22]
rlabel metal2 10528 595672 10528 595672 0 io_oeb[23]
rlabel metal3 392 558320 392 558320 0 io_oeb[24]
rlabel metal3 2310 516600 2310 516600 0 io_oeb[25]
rlabel metal3 392 473984 392 473984 0 io_oeb[26]
rlabel metal2 190680 472304 190680 472304 0 io_oeb[27]
rlabel metal3 392 388808 392 388808 0 io_oeb[28]
rlabel metal2 430738 499912 430738 499912 0 io_oeb[29]
rlabel metal2 516600 310912 516600 310912 0 io_oeb[2]
rlabel metal3 392 304472 392 304472 0 io_oeb[30]
rlabel metal3 392 262304 392 262304 0 io_oeb[31]
rlabel metal2 453978 499912 453978 499912 0 io_oeb[32]
rlabel metal3 392 177128 392 177128 0 io_oeb[33]
rlabel metal2 469378 499912 469378 499912 0 io_oeb[34]
rlabel metal3 2310 93464 2310 93464 0 io_oeb[35]
rlabel metal3 392 50624 392 50624 0 io_oeb[36]
rlabel metal3 2310 8792 2310 8792 0 io_oeb[37]
rlabel metal2 518280 331912 518280 331912 0 io_oeb[3]
rlabel metal3 593082 192360 593082 192360 0 io_oeb[4]
rlabel metal2 519960 376488 519960 376488 0 io_oeb[5]
rlabel metal2 521640 389928 521640 389928 0 io_oeb[6]
rlabel metal2 260778 499912 260778 499912 0 io_oeb[7]
rlabel metal3 595672 350056 595672 350056 0 io_oeb[8]
rlabel metal3 595672 390040 595672 390040 0 io_oeb[9]
rlabel metal3 593082 20552 593082 20552 0 io_out[0]
rlabel metal2 286482 499912 286482 499912 0 io_out[10]
rlabel metal3 595672 455840 595672 455840 0 io_out[11]
rlabel metal2 499128 498400 499128 498400 0 io_out[12]
rlabel metal3 310856 503944 310856 503944 0 io_out[13]
rlabel metal3 595672 574952 595672 574952 0 io_out[14]
rlabel metal2 562632 593418 562632 593418 0 io_out[15]
rlabel metal2 332962 499912 332962 499912 0 io_out[16]
rlabel metal2 430136 557340 430136 557340 0 io_out[17]
rlabel metal2 363440 595672 363440 595672 0 io_out[18]
rlabel metal2 356314 499912 356314 499912 0 io_out[19]
rlabel metal2 217336 500318 217336 500318 0 io_out[1]
rlabel metal2 230888 595672 230888 595672 0 io_out[20]
rlabel metal3 166432 590184 166432 590184 0 io_out[21]
rlabel metal2 379218 499912 379218 499912 0 io_out[22]
rlabel metal2 32480 595672 32480 595672 0 io_out[23]
rlabel metal2 394954 499912 394954 499912 0 io_out[24]
rlabel metal2 402402 499912 402402 499912 0 io_out[25]
rlabel metal3 392 487760 392 487760 0 io_out[26]
rlabel metal3 392 445592 392 445592 0 io_out[27]
rlabel metal3 392 403424 392 403424 0 io_out[28]
rlabel metal2 22680 440216 22680 440216 0 io_out[29]
rlabel metal3 595672 99344 595672 99344 0 io_out[2]
rlabel metal3 392 318248 392 318248 0 io_out[30]
rlabel metal2 448882 499912 448882 499912 0 io_out[31]
rlabel metal3 392 233912 392 233912 0 io_out[32]
rlabel metal3 392 191744 392 191744 0 io_out[33]
rlabel metal2 472234 499912 472234 499912 0 io_out[34]
rlabel metal3 392 106568 392 106568 0 io_out[35]
rlabel metal3 392 64400 392 64400 0 io_out[36]
rlabel metal3 2366 22904 2366 22904 0 io_out[37]
rlabel metal2 232386 499912 232386 499912 0 io_out[3]
rlabel metal2 240394 499912 240394 499912 0 io_out[4]
rlabel metal2 247842 499912 247842 499912 0 io_out[5]
rlabel metal2 255682 499912 255682 499912 0 io_out[6]
rlabel metal2 263704 500374 263704 500374 0 io_out[7]
rlabel metal3 595672 336728 595672 336728 0 io_out[8]
rlabel metal2 279034 499912 279034 499912 0 io_out[9]
rlabel metal2 212408 392 212408 392 0 la_data_in[0]
rlabel metal2 337400 198730 337400 198730 0 la_data_in[10]
rlabel metal2 354536 102480 354536 102480 0 la_data_in[11]
rlabel metal2 281960 5670 281960 5670 0 la_data_in[12]
rlabel metal2 287448 8302 287448 8302 0 la_data_in[13]
rlabel metal2 292712 392 292712 392 0 la_data_in[14]
rlabel metal2 350840 112210 350840 112210 0 la_data_in[15]
rlabel metal2 304304 392 304304 392 0 la_data_in[16]
rlabel metal2 310520 3318 310520 3318 0 la_data_in[17]
rlabel metal3 357952 197064 357952 197064 0 la_data_in[18]
rlabel metal2 321944 3150 321944 3150 0 la_data_in[19]
rlabel metal3 216944 5096 216944 5096 0 la_data_in[1]
rlabel metal2 327544 2758 327544 2758 0 la_data_in[20]
rlabel metal2 333144 7350 333144 7350 0 la_data_in[21]
rlabel metal2 339080 5726 339080 5726 0 la_data_in[22]
rlabel metal2 344792 3206 344792 3206 0 la_data_in[23]
rlabel metal2 349888 392 349888 392 0 la_data_in[24]
rlabel metal2 356104 3990 356104 3990 0 la_data_in[25]
rlabel metal3 379288 198184 379288 198184 0 la_data_in[26]
rlabel metal2 383096 102130 383096 102130 0 la_data_in[27]
rlabel metal2 373352 3598 373352 3598 0 la_data_in[28]
rlabel metal2 378392 392 378392 392 0 la_data_in[29]
rlabel metal2 224840 2310 224840 2310 0 la_data_in[2]
rlabel metal2 383880 392 383880 392 0 la_data_in[30]
rlabel metal3 391272 12936 391272 12936 0 la_data_in[31]
rlabel metal2 396536 198338 396536 198338 0 la_data_in[32]
rlabel metal3 401184 4200 401184 4200 0 la_data_in[33]
rlabel metal3 404656 4088 404656 4088 0 la_data_in[34]
rlabel metal3 405160 197064 405160 197064 0 la_data_in[35]
rlabel metal2 407288 102186 407288 102186 0 la_data_in[36]
rlabel metal2 424536 4214 424536 4214 0 la_data_in[37]
rlabel metal3 426384 6104 426384 6104 0 la_data_in[38]
rlabel metal2 435960 3150 435960 3150 0 la_data_in[39]
rlabel metal3 274456 44520 274456 44520 0 la_data_in[3]
rlabel metal2 422744 102984 422744 102984 0 la_data_in[40]
rlabel metal3 446712 6776 446712 6776 0 la_data_in[41]
rlabel metal2 453096 4102 453096 4102 0 la_data_in[42]
rlabel metal2 426104 104650 426104 104650 0 la_data_in[43]
rlabel metal2 428792 105490 428792 105490 0 la_data_in[44]
rlabel metal3 469168 7000 469168 7000 0 la_data_in[45]
rlabel metal2 475664 392 475664 392 0 la_data_in[46]
rlabel metal2 437528 198912 437528 198912 0 la_data_in[47]
rlabel metal3 463736 195720 463736 195720 0 la_data_in[48]
rlabel metal3 492240 4760 492240 4760 0 la_data_in[49]
rlabel metal2 236264 4102 236264 4102 0 la_data_in[4]
rlabel metal2 498008 392 498008 392 0 la_data_in[50]
rlabel metal2 447608 199010 447608 199010 0 la_data_in[51]
rlabel metal2 450296 198954 450296 198954 0 la_data_in[52]
rlabel metal2 452984 198786 452984 198786 0 la_data_in[53]
rlabel metal2 521192 392 521192 392 0 la_data_in[54]
rlabel metal2 526568 392 526568 392 0 la_data_in[55]
rlabel metal2 532784 392 532784 392 0 la_data_in[56]
rlabel metal2 538776 2702 538776 2702 0 la_data_in[57]
rlabel metal2 544432 20160 544432 20160 0 la_data_in[58]
rlabel metal2 469112 197946 469112 197946 0 la_data_in[59]
rlabel metal2 241864 1582 241864 1582 0 la_data_in[5]
rlabel metal3 472360 198184 472360 198184 0 la_data_in[60]
rlabel metal2 561624 2702 561624 2702 0 la_data_in[61]
rlabel metal2 567560 2310 567560 2310 0 la_data_in[62]
rlabel metal3 526400 190680 526400 190680 0 la_data_in[63]
rlabel metal2 326648 198338 326648 198338 0 la_data_in[6]
rlabel metal2 329336 194530 329336 194530 0 la_data_in[7]
rlabel metal2 259112 2310 259112 2310 0 la_data_in[8]
rlabel metal2 264824 2310 264824 2310 0 la_data_in[9]
rlabel metal3 212520 25144 212520 25144 0 la_data_out[0]
rlabel metal2 272440 2310 272440 2310 0 la_data_out[10]
rlabel metal2 277536 392 277536 392 0 la_data_out[11]
rlabel metal2 283864 3206 283864 3206 0 la_data_out[12]
rlabel metal2 289576 5838 289576 5838 0 la_data_out[13]
rlabel metal2 295288 1470 295288 1470 0 la_data_out[14]
rlabel metal2 351736 118930 351736 118930 0 la_data_out[15]
rlabel metal2 306096 392 306096 392 0 la_data_out[16]
rlabel metal2 312424 5782 312424 5782 0 la_data_out[17]
rlabel metal2 359800 109746 359800 109746 0 la_data_out[18]
rlabel metal2 323120 392 323120 392 0 la_data_out[19]
rlabel metal2 314104 197890 314104 197890 0 la_data_out[1]
rlabel metal2 329560 98070 329560 98070 0 la_data_out[20]
rlabel metal2 334712 392 334712 392 0 la_data_out[21]
rlabel metal2 340088 392 340088 392 0 la_data_out[22]
rlabel metal2 373240 197946 373240 197946 0 la_data_out[23]
rlabel metal2 351624 392 351624 392 0 la_data_out[24]
rlabel metal2 357896 98182 357896 98182 0 la_data_out[25]
rlabel metal2 380184 198296 380184 198296 0 la_data_out[26]
rlabel metal2 383992 102242 383992 102242 0 la_data_out[27]
rlabel metal3 377888 8792 377888 8792 0 la_data_out[28]
rlabel metal2 380968 2590 380968 2590 0 la_data_out[29]
rlabel metal2 226744 5726 226744 5726 0 la_data_out[2]
rlabel metal3 388584 52136 388584 52136 0 la_data_out[30]
rlabel metal2 392392 2366 392392 2366 0 la_data_out[31]
rlabel metal2 397600 392 397600 392 0 la_data_out[32]
rlabel metal3 402976 4200 402976 4200 0 la_data_out[33]
rlabel metal2 402808 102410 402808 102410 0 la_data_out[34]
rlabel metal2 405496 198730 405496 198730 0 la_data_out[35]
rlabel metal2 420728 2534 420728 2534 0 la_data_out[36]
rlabel metal2 426440 2478 426440 2478 0 la_data_out[37]
rlabel metal2 432152 3990 432152 3990 0 la_data_out[38]
rlabel metal2 437304 392 437304 392 0 la_data_out[39]
rlabel metal2 232008 392 232008 392 0 la_data_out[3]
rlabel metal2 443576 8190 443576 8190 0 la_data_out[40]
rlabel metal2 448896 392 448896 392 0 la_data_out[41]
rlabel metal2 454272 392 454272 392 0 la_data_out[42]
rlabel metal2 427000 110530 427000 110530 0 la_data_out[43]
rlabel metal2 429688 118930 429688 118930 0 la_data_out[44]
rlabel metal2 472136 25830 472136 25830 0 la_data_out[45]
rlabel metal2 477456 392 477456 392 0 la_data_out[46]
rlabel metal2 482832 392 482832 392 0 la_data_out[47]
rlabel metal2 489272 4046 489272 4046 0 la_data_out[48]
rlabel metal2 494424 392 494424 392 0 la_data_out[49]
rlabel metal2 238168 3262 238168 3262 0 la_data_out[4]
rlabel metal3 500248 4088 500248 4088 0 la_data_out[50]
rlabel metal2 448504 103810 448504 103810 0 la_data_out[51]
rlabel metal2 451304 20160 451304 20160 0 la_data_out[52]
rlabel metal2 517608 392 517608 392 0 la_data_out[53]
rlabel metal2 522984 392 522984 392 0 la_data_out[54]
rlabel metal2 459256 104650 459256 104650 0 la_data_out[55]
rlabel metal2 534632 392 534632 392 0 la_data_out[56]
rlabel metal2 539952 392 539952 392 0 la_data_out[57]
rlabel metal3 544152 4424 544152 4424 0 la_data_out[58]
rlabel metal2 470008 127330 470008 127330 0 la_data_out[59]
rlabel metal3 284256 31080 284256 31080 0 la_data_out[5]
rlabel metal2 472696 197050 472696 197050 0 la_data_out[60]
rlabel metal2 563752 2366 563752 2366 0 la_data_out[61]
rlabel metal2 568512 392 568512 392 0 la_data_out[62]
rlabel metal2 574728 392 574728 392 0 la_data_out[63]
rlabel metal2 327544 192122 327544 192122 0 la_data_out[6]
rlabel metal2 330232 108850 330232 108850 0 la_data_out[7]
rlabel metal2 261016 4830 261016 4830 0 la_data_out[8]
rlabel metal2 265944 392 265944 392 0 la_data_out[9]
rlabel metal2 217224 3094 217224 3094 0 la_oenb[0]
rlabel metal2 274344 4942 274344 4942 0 la_oenb[10]
rlabel metal2 279384 392 279384 392 0 la_oenb[11]
rlabel metal2 285656 90678 285656 90678 0 la_oenb[12]
rlabel metal2 291480 4046 291480 4046 0 la_oenb[13]
rlabel metal2 349944 106330 349944 106330 0 la_oenb[14]
rlabel metal2 302456 24892 302456 24892 0 la_oenb[15]
rlabel metal2 307888 392 307888 392 0 la_oenb[16]
rlabel metal2 358008 110530 358008 110530 0 la_oenb[17]
rlabel metal2 360696 102130 360696 102130 0 la_oenb[18]
rlabel metal2 325752 2702 325752 2702 0 la_oenb[19]
rlabel metal2 222936 1526 222936 1526 0 la_oenb[1]
rlabel metal2 331464 2422 331464 2422 0 la_oenb[20]
rlabel metal2 337176 2478 337176 2478 0 la_oenb[21]
rlabel metal2 342888 2534 342888 2534 0 la_oenb[22]
rlabel metal2 374136 102410 374136 102410 0 la_oenb[23]
rlabel metal2 354312 2646 354312 2646 0 la_oenb[24]
rlabel metal2 359800 4410 359800 4410 0 la_oenb[25]
rlabel metal3 378840 198072 378840 198072 0 la_oenb[26]
rlabel metal2 371448 2478 371448 2478 0 la_oenb[27]
rlabel metal2 377160 2702 377160 2702 0 la_oenb[28]
rlabel metal2 382872 2366 382872 2366 0 la_oenb[29]
rlabel metal2 228536 9926 228536 9926 0 la_oenb[2]
rlabel metal2 388584 2310 388584 2310 0 la_oenb[30]
rlabel metal2 394296 2310 394296 2310 0 la_oenb[31]
rlabel metal3 399112 197400 399112 197400 0 la_oenb[32]
rlabel metal3 404768 4424 404768 4424 0 la_oenb[33]
rlabel metal2 403704 102018 403704 102018 0 la_oenb[34]
rlabel metal2 406392 102242 406392 102242 0 la_oenb[35]
rlabel metal2 422632 2310 422632 2310 0 la_oenb[36]
rlabel metal2 428456 3206 428456 3206 0 la_oenb[37]
rlabel metal2 433720 392 433720 392 0 la_oenb[38]
rlabel metal2 439768 2422 439768 2422 0 la_oenb[39]
rlabel metal2 233856 392 233856 392 0 la_oenb[3]
rlabel metal2 445480 2366 445480 2366 0 la_oenb[40]
rlabel metal2 451192 3206 451192 3206 0 la_oenb[41]
rlabel metal2 425208 102130 425208 102130 0 la_oenb[42]
rlabel metal2 427896 105546 427896 105546 0 la_oenb[43]
rlabel metal2 468552 2086 468552 2086 0 la_oenb[44]
rlabel metal2 474040 3262 474040 3262 0 la_oenb[45]
rlabel metal2 479248 392 479248 392 0 la_oenb[46]
rlabel metal2 454440 107856 454440 107856 0 la_oenb[47]
rlabel metal2 490840 392 490840 392 0 la_oenb[48]
rlabel metal2 496216 392 496216 392 0 la_oenb[49]
rlabel metal2 239176 392 239176 392 0 la_oenb[4]
rlabel metal2 446712 198842 446712 198842 0 la_oenb[50]
rlabel metal2 449400 161770 449400 161770 0 la_oenb[51]
rlabel metal2 514248 2030 514248 2030 0 la_oenb[52]
rlabel metal2 519736 3150 519736 3150 0 la_oenb[53]
rlabel metal3 521920 4088 521920 4088 0 la_oenb[54]
rlabel metal2 531384 2254 531384 2254 0 la_oenb[55]
rlabel metal2 536872 2534 536872 2534 0 la_oenb[56]
rlabel metal2 542696 2478 542696 2478 0 la_oenb[57]
rlabel metal2 540232 4256 540232 4256 0 la_oenb[58]
rlabel metal2 470904 198562 470904 198562 0 la_oenb[59]
rlabel metal2 245896 280 245896 280 0 la_oenb[5]
rlabel metal2 473592 102186 473592 102186 0 la_oenb[60]
rlabel metal2 565432 2310 565432 2310 0 la_oenb[61]
rlabel metal2 571256 98070 571256 98070 0 la_oenb[62]
rlabel metal2 576520 392 576520 392 0 la_oenb[63]
rlabel metal2 328034 200088 328034 200088 0 la_oenb[6]
rlabel metal2 257208 7462 257208 7462 0 la_oenb[7]
rlabel metal2 262360 392 262360 392 0 la_oenb[8]
rlabel metal2 336504 107226 336504 107226 0 la_oenb[9]
rlabel metal2 580104 392 580104 392 0 user_irq[0]
rlabel metal2 581896 392 581896 392 0 user_irq[1]
rlabel metal2 570360 100912 570360 100912 0 user_irq[2]
rlabel metal3 214200 198184 214200 198184 0 wb_clk_i
rlabel metal2 216440 115570 216440 115570 0 wb_rst_i
rlabel metal2 22680 98672 22680 98672 0 wbs_ack_o
rlabel metal2 23016 2366 23016 2366 0 wbs_adr_i[0]
rlabel metal2 87472 20160 87472 20160 0 wbs_adr_i[10]
rlabel metal2 93464 2758 93464 2758 0 wbs_adr_i[11]
rlabel metal2 98168 392 98168 392 0 wbs_adr_i[12]
rlabel metal3 258272 197176 258272 197176 0 wbs_adr_i[13]
rlabel metal2 262136 186970 262136 186970 0 wbs_adr_i[14]
rlabel metal2 116032 20160 116032 20160 0 wbs_adr_i[15]
rlabel metal2 121352 392 121352 392 0 wbs_adr_i[16]
rlabel metal2 126728 392 126728 392 0 wbs_adr_i[17]
rlabel metal2 132720 4200 132720 4200 0 wbs_adr_i[18]
rlabel metal2 138320 392 138320 392 0 wbs_adr_i[19]
rlabel metal2 30352 20160 30352 20160 0 wbs_adr_i[1]
rlabel metal2 144592 20160 144592 20160 0 wbs_adr_i[20]
rlabel metal2 149464 86128 149464 86128 0 wbs_adr_i[21]
rlabel metal2 283640 195426 283640 195426 0 wbs_adr_i[22]
rlabel metal2 161504 392 161504 392 0 wbs_adr_i[23]
rlabel metal2 166880 392 166880 392 0 wbs_adr_i[24]
rlabel metal2 288120 165928 288120 165928 0 wbs_adr_i[25]
rlabel metal2 178472 392 178472 392 0 wbs_adr_i[26]
rlabel metal2 185640 90328 185640 90328 0 wbs_adr_i[27]
rlabel metal2 190568 2254 190568 2254 0 wbs_adr_i[28]
rlabel metal2 195440 392 195440 392 0 wbs_adr_i[29]
rlabel metal2 37464 392 37464 392 0 wbs_adr_i[2]
rlabel metal2 305144 193802 305144 193802 0 wbs_adr_i[30]
rlabel metal2 307832 195482 307832 195482 0 wbs_adr_i[31]
rlabel metal2 45528 20160 45528 20160 0 wbs_adr_i[3]
rlabel metal2 52640 392 52640 392 0 wbs_adr_i[4]
rlabel metal3 236152 198184 236152 198184 0 wbs_adr_i[5]
rlabel metal2 240632 198786 240632 198786 0 wbs_adr_i[6]
rlabel metal2 69608 392 69608 392 0 wbs_adr_i[7]
rlabel metal2 75824 392 75824 392 0 wbs_adr_i[8]
rlabel metal2 81200 392 81200 392 0 wbs_adr_i[9]
rlabel metal2 218232 103138 218232 103138 0 wbs_cyc_i
rlabel metal2 24920 4830 24920 4830 0 wbs_dat_i[0]
rlabel metal2 89208 392 89208 392 0 wbs_dat_i[10]
rlabel metal2 95368 3206 95368 3206 0 wbs_dat_i[11]
rlabel metal2 100856 77070 100856 77070 0 wbs_dat_i[12]
rlabel metal2 260344 198730 260344 198730 0 wbs_dat_i[13]
rlabel metal2 263032 112210 263032 112210 0 wbs_dat_i[14]
rlabel metal2 117768 392 117768 392 0 wbs_dat_i[15]
rlabel metal2 123144 392 123144 392 0 wbs_dat_i[16]
rlabel metal2 129360 4200 129360 4200 0 wbs_dat_i[17]
rlabel metal2 264600 192416 264600 192416 0 wbs_dat_i[18]
rlabel metal2 140112 392 140112 392 0 wbs_dat_i[19]
rlabel metal2 32088 392 32088 392 0 wbs_dat_i[1]
rlabel metal3 144648 4088 144648 4088 0 wbs_dat_i[20]
rlabel metal2 281848 114730 281848 114730 0 wbs_dat_i[21]
rlabel metal2 284536 175210 284536 175210 0 wbs_dat_i[22]
rlabel metal2 163296 392 163296 392 0 wbs_dat_i[23]
rlabel metal2 169624 2254 169624 2254 0 wbs_dat_i[24]
rlabel metal2 174888 392 174888 392 0 wbs_dat_i[25]
rlabel metal2 180264 392 180264 392 0 wbs_dat_i[26]
rlabel metal2 186760 2254 186760 2254 0 wbs_dat_i[27]
rlabel metal2 191856 392 191856 392 0 wbs_dat_i[28]
rlabel metal2 303352 118090 303352 118090 0 wbs_dat_i[29]
rlabel metal2 40152 2254 40152 2254 0 wbs_dat_i[2]
rlabel metal2 306040 192962 306040 192962 0 wbs_dat_i[30]
rlabel metal2 208824 392 208824 392 0 wbs_dat_i[31]
rlabel metal2 47264 392 47264 392 0 wbs_dat_i[3]
rlabel metal2 54432 392 54432 392 0 wbs_dat_i[4]
rlabel metal2 238840 182770 238840 182770 0 wbs_dat_i[5]
rlabel metal2 241528 199570 241528 199570 0 wbs_dat_i[6]
rlabel metal2 72296 91350 72296 91350 0 wbs_dat_i[7]
rlabel metal2 78232 3990 78232 3990 0 wbs_dat_i[8]
rlabel metal2 82992 392 82992 392 0 wbs_dat_i[9]
rlabel metal2 26824 2310 26824 2310 0 wbs_dat_o[0]
rlabel metal2 91000 392 91000 392 0 wbs_dat_o[10]
rlabel metal2 97272 2254 97272 2254 0 wbs_dat_o[11]
rlabel metal2 258552 105490 258552 105490 0 wbs_dat_o[12]
rlabel metal2 260834 200088 260834 200088 0 wbs_dat_o[13]
rlabel metal2 114408 1470 114408 1470 0 wbs_dat_o[14]
rlabel metal2 119560 392 119560 392 0 wbs_dat_o[15]
rlabel metal2 124936 392 124936 392 0 wbs_dat_o[16]
rlabel metal3 201544 21000 201544 21000 0 wbs_dat_o[17]
rlabel metal2 136528 392 136528 392 0 wbs_dat_o[18]
rlabel metal2 142856 89726 142856 89726 0 wbs_dat_o[19]
rlabel metal2 33880 392 33880 392 0 wbs_dat_o[1]
rlabel metal2 148120 392 148120 392 0 wbs_dat_o[20]
rlabel metal2 282744 104706 282744 104706 0 wbs_dat_o[21]
rlabel metal2 285432 106330 285432 106330 0 wbs_dat_o[22]
rlabel metal2 165816 4046 165816 4046 0 wbs_dat_o[23]
rlabel metal2 171416 46830 171416 46830 0 wbs_dat_o[24]
rlabel metal2 176680 392 176680 392 0 wbs_dat_o[25]
rlabel metal2 182056 392 182056 392 0 wbs_dat_o[26]
rlabel metal2 188440 8246 188440 8246 0 wbs_dat_o[27]
rlabel metal2 193648 392 193648 392 0 wbs_dat_o[28]
rlabel metal2 304248 115626 304248 115626 0 wbs_dat_o[29]
rlabel metal2 44520 30632 44520 30632 0 wbs_dat_o[2]
rlabel metal2 306936 125650 306936 125650 0 wbs_dat_o[30]
rlabel metal2 210616 392 210616 392 0 wbs_dat_o[31]
rlabel metal2 49056 392 49056 392 0 wbs_dat_o[3]
rlabel metal2 237048 197946 237048 197946 0 wbs_dat_o[4]
rlabel metal2 68040 33040 68040 33040 0 wbs_dat_o[5]
rlabel metal2 68712 2254 68712 2254 0 wbs_dat_o[6]
rlabel metal2 74424 2254 74424 2254 0 wbs_dat_o[7]
rlabel metal2 80136 2254 80136 2254 0 wbs_dat_o[8]
rlabel metal2 85848 2590 85848 2590 0 wbs_dat_o[9]
rlabel metal2 28728 2366 28728 2366 0 wbs_sel_i[0]
rlabel metal2 36344 2422 36344 2422 0 wbs_sel_i[1]
rlabel metal2 43960 2478 43960 2478 0 wbs_sel_i[2]
rlabel metal2 51576 2534 51576 2534 0 wbs_sel_i[3]
rlabel metal2 219128 198786 219128 198786 0 wbs_stb_i
rlabel metal2 21112 2254 21112 2254 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
